

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
IjW7TWFm3KgKMVpjP6ygVFbznd+FPstRLfWNqknIMyJ8+Petd/t/6GqRoQyK0IrljIinM2bdWJa0
fDJ3MPtw9Q==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
UvNKMyHYO7foasAmwmJQ3tldmK5UlvU00Hek+aRbgGk6YIL2wKvqcEPGh5ETO74ijwGAvqxMIzHY
TFltBE6SamLP/WdNmQrPYW7w3MUsI0kqOCrTm8t/idnF9PrPu7oGcqQOKgEL9TdLr8AiGPxMaTqm
RolVqrL5+MLQUExAiEI=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
PNtXSVfX23+g2jfFVAmY1gVTdgATPD6Pj0CvTFTcyjPgCqWueeWwGxBdUCyveVP0AR4AXhg5BMqS
swJmZHRRVxLK7chH1J36nBeqWcV4Cq9cum1SQO3mjOEFHjjww1gv3Syi5yvtavbjLEw67RPpAjWb
wGU7QnwyMZx9hDqpFP3fyW90vL4XtJgukKYllA0qQBTiSmrBn21pyJ9cYMDxpvvQP5BV4NShpZhg
zzkA1x8gP9y4KQI9v14pxrT0WuSxZryUyPmQ5W9a6Y8hhu2e/avBbJfLfFK3LQs0GjiyU5OCYucA
xgLgol580NBlFGs4egghWLU2W2ZIG3bP365kcQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
4NMgVcG/CD5nY3o8ZGR40DBBMRryZWMdVNLVI7r/3Eqjonb7qXBHUdyBMZ2ZrEGS2SvsDUjJgBhV
7Ye2FRVYMA6C8fO9Gvvb/NTvkgPEUt3/CpLmvd6uHfzJhZpCPgOZizH7l8eVTs5/5Dzk3s8Lb1+v
McDyUPxs7gWYFY6Kt/s=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CYzL6f5k8iw0M4OnZdKWiKrhYgoEN5rM49URJ4pWhYABCXwsXbzkKBP1HKzismQoFmpnCYp7gP2y
8XHYPCjw5cgF0kN+RIbqzAue/ip6jOWpvxh52l+Dr1FKbEKKlc+eGqdiUyHqyWhyXk7kS1rnL2M0
dPIhHdtAg45aF3CV9I0Yfm785rvdlRxCuJxvYysuQmn7I9400WGnoDreoZy8TyJwVpKslU++ac0z
NMGJiqWSaJ5BtPnq22hKmi0+OI1P20R1Tb3MR/4AkIXR599Mw72F3kOIfreQDWeUyFpuumt3Ih8v
i9EtFKN0BDgWwg4dPIqAasEI9Dq2Y2YFyfIArg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
n39IbVRxNKZUsCubowTOOzNhNKrmcNv6OW9lv+Cdwtajc3xH44RGP8csfxiS2Vot0/o1hPNTds6Q
i9DjURZuo/DvgqI78TPWwH05tplCjF7YcWQT1m7pL2ByzPcgtdMJzS3ntk6kIvluRN1g+EqNtNQn
+ZbS+aNTF9yaB3l4/MmTSW1lzPrFdFNmEP8V+78jFSDjYYSdZB4nBJ0hkjbBWNGp1ANOLzYbAv3J
n4nd6wlsQpTbPQRKUcvjIwL2GA1XrlDW9MpyoUdJR0TSc4csSnUfQpcya+VvpkcbgA5MF1EuObkG
FqQJHPtbbC/CLIorgSIgCDIQsvlH7wvr8D7S7Q==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 425872)
`protect data_block
eCzUWnw+8Rpc3KguUrIuRlk6B3XlfzD/zgfk4gzs86FdocAztCAc9Dk4aVgU2jFfbUYN+u8XCn5c
fI9De7ZP9NXG/OlAHxsNfzkLaDDEXbVYHAWAOZk+1Z94WwjChJr1Zr/2y1ZNo9q4HZbrimkxnPFT
Rk/VqWFiA0MBpRnlLPOlRv7eU4vY6f5VUdw8QlGdHK436bSHajsrP0tcXy/8ljbmehgZUq2PT0B0
vGX4hUV02DVngIzkwUBnvHEKPkilwD39RMmvRkBzkg3pI81FvsXw3SwEkxPrgx8s7Yp24jLof2As
v60WNQCnsIITyg7IldniZry4OWxEov8dhD4ywwRthrN9syudcx+qskbDTJMMRZVld0Q0j/s8M/1Y
pcznAsajVaF9b1OeM987VUn9JKHOtWsupITzX7oX1REWNhY7dbktYLR86TbdJkZoKhtRd8/3Y+FN
QhPE77f15jNw4JW2dH4AJH78Rs1Sb3zXRN5S401zjMJtYgoxV6DI4UPdNsVC/XuXPvaUFgjgj9X6
V92jmQducEGJFsmJazJTfGKmRP2EZHwvikioMm5a6VomOj058LFvq3xR3WxzBXa3lWKf3wA3Tc6x
w6QnP8Aj2IgFXiYv9eC74ePSQFA732llKNRdbEHKkm1VyeCIwP4Crx4PbbNpvUgrysNXtBS+wEfz
5hcdzSoDVuyfPGQlPoY57sziWUArCQq0Orerz24p6v+zH3EDATr8tDmvTndf59/OuPrxNEdKCUX0
Ko+nGhrDP2GEIog4xqFf6rW/WYI4rMqmvMlfb3nKNWQZocl9IM+bb7qJFQ9AmjwcNTSmpU5BvoyX
yAmh2nVXUmIxYQbv4B5dCn+ey3E2pWZLaHMzd8xOJGDcpTQdxa5UVjmQJhMqJBSDJGQIEa5h6FW5
vSR5y7DP8wnKl3DGbIDoGVb67k0x2ss/DcBEMlTYVDfIDdZsCOhrksr4jrnfsu2ZRdznLuH6arFp
cyuAQj6uvrotaAGisW7uaC2YU3nmc+l5Jz/hEzsJoXlyN0diN7FzxIxnf0WFacUp3ATCl15wwtE5
M08tXLMKZu4UvMY6Zo7PQ8JwBpnqXdCmYj1oqP1JaNsIRDQpKyfTXGgvW63dKi4O4zeTd0f0W7Zo
MCR7O6aYYCVt0dxLSVvw62euyT/oDb/5RZ4TXKlyM2Tt84eJEumoHlKRkvLZtHha3pnGbxPBpSkH
7v1n3qiZW5dL38ONCHrNdJg5GMZuvh7HydmebGtUvj8wKi717eLBeXqbYDl1XfY1XVt4SBXKCkpT
49/gpNHshiz4JMFLXQHRheZzaAOBDoS85+mwBN41Gsxoc+9rukqO7Yrbd6xIk3IPD5mDp5UmCoOw
ZeI2VVjBfg9mqS/a7B1/x9Z9U7dHHMynz4+2hZyxZXSNyJj0z8U8zfOAsn4hp0LlvNXqox/HIP9T
C+YUNRyDCFg8kR7GdlFh6WcmExb8dOaCeNTCoMhscQU6zSXaV6y1WB4f2k2PW51W6cr2JNMv1IKS
qiXCsbkxr/gYvTNZ5dRgtfDh7lhIX5cGCT463gnFqb3YdzUeaTlp18xIdO+ZT6TsgKWKMgbJ6lvB
Bs2A6sW7nN60FVZn7M5XgZD3hl7AChgw85i+KZBrrbpnK9BC/821PZ+Prif1laoAN5O1C2kGwauY
A3UYWZEJyDR/IPoEbwPwY/t5yXpX7n6rtTSIz0MMzDSD24F/8gv8jDYS+FuaVI8UZ1DX7VuIDDzJ
Pq2OpXHQsChsanOeZfhasVzK/As/ZbW8VhNjTv5ilZN7DIFFQNY/lVIPzbaBvNYUQEJ6EupfS/mt
zK+EZfRGHDYYzSSSgibJaSWZGqPHqcCy0AGyqWg130coRW5nL8W4J9CDnc/4rkdGJG7s/3BatWIX
VFASiUcM6ay16/leDchf+45/y45Ajs/ZL6n+TBmNTsMlAMm6X9tyOKg6BHeOvu+ybWtw7eeyHvb4
cDetMs3acyJsL4EgJF4tSMxwF+USkySSNJnzRjrtQjL67j0QReUlbFTa1HQNSLmxuobK2fAz8qCU
lUI9hNmb3BCU9tVLShSGs4VjtcxVa4gybwSKr9rVa4fHo1xPA09ZSHzYvYn/rlS2M/9icsYztNLe
5gJLsgu6Sl8PsjZqXW0ZemMxPIX8W2YxbOalS3CHVM/GNjy/XeeElxNCIzXqpg1nh6XDZ5tutUG2
wfROMijuaBqoXvKB1ZEb7FXzrWhaGrMf3GhHqjPavJlfkFdH9h+RP2wvRgzNH1imnDPLpiBTi7W8
qwSktfkKS8UxJcGqdGxqCgCE5zvKPxNPf3Fyng+/ZTcDANfdC3Ssljl1wC6FyT/Wp4Y7nrVTQoYc
AA5o0dFtLMLPfoa7bgzGd6DwambNWar1g0rcEJHht9SNGPH+6bFaCXzgkV7ltjNiwdOr2atrCpIW
f+3ugvI8fY4maPTG4keTURY61qvIRCVOXuuSLlm9DuPGi1GLt5aMv6mp+ly1Q88Ti6oHBHHuuj0Y
sBvN3ECxr8KtGcvUp0mBYh3ycOFHtOlgs915Z/dsNqnwno63BBCtHZkMQUi2AF4VpcMo2KMFTCmm
tvzaFGE5RksjjGwbz51D5JiQVot9TOWVDhcffUwzw13pehzQpmN7C4I7Y5eBvX+XP5eBIYd0ck1q
wXs+hdcjMtJZMFOn9DDzVcZsHomEpeX9IK6pIGB3wkVTvmwiSMSxzL0geCROPY4wY50brCWofMqt
tQTcdtJocBD3SSmi5gqWPyTqSP/2bO0758EimMxnFWN42nPTqhVHVu+cSiQhmCraNNvPsr5+dptM
8PLt6Z/OpX4+LJn5uwmzpFwxeFa/T2N2RF5LjprBQIFXuZZJfLtIfSnAWbnPmsODWsLXCbXV1wxu
0GCykxb4+53cESMaYQ9v5HeYJUHabmWDgXFjsIzFL6dHlh1TPzlECci8tTw3CUxWDsobKLBuct4J
ec4AIoBAqANYNe3zj6wyKztc+EaU8UQZNPZIRSpE8OuKdwKrzymdOzBuz5M3LO3gZkKNGLcfTO0a
JaRUUk2Nqe6815o1j2ACj6fYV5sO3atVVu0vy9B8g8NrGwkFnmVu+I5jB8cApo8q0q2i5mPI+vyF
iInOuzWaRP3ROdMq3OljoHR1NdeANAGHSfzwuhPcjh9Wb4xukXE86IzASZHWmigpgchnL3Y9bdNp
GK7rmwXP0jUL630RSbzKhHkiFfnTkeTqgkq7X+zidcyPyLqd5qlnyRsXNaLZczQRIiHHUp2u1Drd
ugpqC9XIHEJpmhMhZog3mHyK7dXEDa0m4IDGgDjRCisIs34wm/p5N4aU40ArWNNlEALXlxMJXhn1
xqizO3vt6azAPjr9KGPSnoX7ddDfJSme2ZHrZC+OR3VCmiDGs3iPg6J/RtcTpyR0HWzjhbSYSMIc
1rEBFePRISMnbtUWj0Y/XZZWPAOvaRecu9TaBYogzK5YTSgGnR9geE8Zakengr86/vy7wAdQQcU+
p6rd2cSHEL1f/XfjsYp+oJd+OJvhO8yWl6wfAaWou/Igw0iW/frNTgRZkfD07E96T8c9zeBxi1+k
IX6EqO1yPEFmC2HKxgd0Fvz9mHlO/AYG74OIwGwa0l3CUlqcg3IdRR0XOhX66S1ic+00gnA3bUGa
9e2b87eyZGDfiH89h/NNQvTMvS2aaZTh05gmKXjm3X1AfjsQncl10OBgJnQVZd+2uSTtBuVlhU6a
kBpBg0KhEmP4W+lBQ0icBcK+5R+JUS8pP4pNFPNo50s260MCPohBwojW/O/jfE6E6w1oRH9I9fAx
KmSf1/WqoZZbqiTBPkp2jZDmsIz3AaHroqxYiYrUUGjJdNTkXWec9yVa7YLHsryS0HWleXNpQ5TK
FOrI9o5U5dSkuNC48dx0LFXvR3b9cmofbVxxn3kmXUXgI3HK4CfHi5HiJ3tG3mDLdtrn68qXW+Ka
NeSBGmfso3hEXZ+Lm8uUvCimwSA0cirRumwAdHZpcUfPD0dP2eSruwyHGgAkCrOIp7yyTpjfRoCz
RjRTdIqhTfJF0uSBZ/CVB6fFQudVWBSZutPDni2mqacObNiL7vzAy+MF1mn3VZTuJHWEYRMCP7VU
hpSy+bLPhzlXT9OOzYslTATRau1ARn6iRGXK0k9aaB5qEx2XCsDbtxg0k+HjLOC/fWT/3g0JZ4q4
ZnBugWLTDal2vI5lvcOCzhxB7ElWCKVa8qQfWEQpiv5YwLDwXB3umVBkIv0k4ldHOK0LEpuXG8MP
cBrMNny/aW2hFNYe40OB9KhJggmvrtN89HyVAdkV15iuaN6/PndLXwLGx6S8GrMR42hyRAzfCs3g
BusbKwjpbk/sVGYZvFoctA8clpSz1wafRugkRSt2YT7xAE6Xl7gJ50EUFqE7E5WObTE5TiD8XoEZ
+WePTy8DInhw3xvyirphNmzvJZ8rzZbjgWSN4Ccqzw1uGxk548rFOnfCg+59XE325nz10Up7ulmB
YU9YP7W8C3vbNXPdGJVoA0qG+mEVVnnlBvnL2gVC1V4l0wQG6epS4eFr7TsJlQEzOKtN0QVw+PXY
Y3LSTYvTjrH77nJKhKMuadMM9gCaqqQWfrfWMlSWKFAKKHSOXwc9yP3H03BCyqAkKerw5MYGeFIq
33pwg1p9rBuTtSQkN/LKNj+b9mVAqMtBmYJRRKI/YLYpCJGnFiHd5Pjgqs99TOO9RoSsmNCSfjn0
oqZNUQ7jA6u6Wg9Kp2Dfe7baWJRF/MtvWJ8hNn32uGEGpeiztTzjT/UHq4X8PMq9roj5cZt5az2n
rfKGybqCVwboPaOJefgN0IZUO2xy2m7wZNlBP0LTkfGatJ42Jt3UOoFx7GIweYI/K/fOtLKr9tkO
0CRJTjbbb/0FXTyepa15N/tBo/nlmLjmb3mdLgt+YkYAjzvsi2dtPQDux3hxMhL9FZVjYQU3g+0A
0D9WmyuVBUDoYnNAmTWYDZmZePH5RW/+X8SDwBrszPj7LFCp4xr1sJ1aOSAoU2nBUYwV0PG0yF3H
Ig4ftVLSPBli8uiL9ExLLlST+Ob/ygmIAlGJEvw1mzk+CzzJFlqwTatJx4bHaP/I8K3i/b59mmwd
rAfRlIiRx8ZyBnKIk6P8njiFssJUZm5H39LVSGTPwttGkTEVY8OOLXpulAsoz5ImbTjvhoMvfTpB
bySerNEvXEG8+eGTtdFPLC/eNJ/udbl/Cg1p3wH59Tt/iyPkGX0X9Q3U0uEmeJIHB+tpaQrYYWut
1WIYM0RP5Paxz4ghMzP61IwgMORYi352EqWPkd31kzQqJRIkiHV0u6PloSgOODxBjmpktJDA9YHr
tBmoI3wtJfZhhOGWKTTdcw9rbS9pTw7U5jAPtPHzISAJPG24ZRoouzxAXF121jo9NvmZJHgiHxfd
tMfHV3N3GOwXh8VsnuDnP2/QAbPrgJGOtbxghncPohUYkkIGia6w/cC8Ke1EoqQiM/UTkJG6QnaX
QV09Mw5eihC9n1VBVrv5u0d1eYsOBh4Bgj8nYJsutxbZf4dkZS/9veCXpWE8/h5goVskq8wchzWA
xk3ZXMPO+m0UaiPh1JhBvy6B2G8GkckVTfjbLXl1ltVddGUbbeQhazWBCrVaoJHZkUT/Y2CP0r7K
KFZi1rQNOZ0ggSiu7HADNwPgZPyTB2qbr32YrZ8mxSnGabDTC655814qtgEtqlKuFmn6I1+3DTTp
SgHAZgswg/fPVTJ1L5+QJps7KRb4OaQ7x5K/JjK+Uk2ul7yL+BB8wX3oU8pzgfgNpMYnZ6NcspJn
4TjKTJn8LsrEj4tNabDNpnjRZzliuUE0LqZWMLP83fd+T0yn5Xssp9/nICReu/4uLbhtumNwgsVW
FGnfX6uUwKuOOEM5yzXUxNQaEChFjcqvySJcQKWmgC5OcJ7dYuhHW7fwZWQc6wjIasuzgP3hKikk
3UotmfgIMKSoJotub8zPl3+lyTuo8VeiseNtI6F6e8/K3YZoLHbthYBqXKBgD13Nty0fy2JQeFLj
YVgZwI1XQBwW6O0eYD+uiUuOdRc7/K51d+5Vh+chbdCVRbMjReq2T3AB2kmzPTu9oy61MfDm1Hed
YsmENRZbyFsEenfYq+/dxwWpJh7EhIy4ko7XcguRndfuTlnvpk3Ezhf//UldssWGJ5D0U3Vy0FKM
Oe/hseIlPgRhotoQzGSuIr6GWI/AyqmFswDhc88nrOpPPQt5yOU0K8gxzZ862eeJ2kdKgWmwi7Fz
lAtwdySoOUarQyhA2/uG7LiBya3A+0A9nhOP6muDJSFbsISxriKH3QUmT00g/cyYA4r30lvdfTyw
5YOEcrWUP0aJYrz0/BaroAXlZcx81e65foZoKWVVn/XloAeGSujjZfnBcnD3ZWZO0umIbUquUIBK
VFOF/FpCFhwYnhzKH2yromWhSEBAMZw5uJykt6NZLk6BVNY9uF+tyaOicJ9yLivpmG8XzQlAe7ZS
lJXCuuTv4f86qm0Tukn2QpjVAgTIzxjYb3K/x3mY3ZvbzLwx1CS90w4iaTc6/cEYn+0HsQN3dxtr
vrT/i275Ub9KCHBLkGq+kMTvHO/o2dHDcPWbNN1Gb1Qv/9ziMc2jHvkEGTfVstylTCFqqXaT3LRF
oV0CHQMedCP/alAaFlGxxO+dzrZn0WLbvNagYgVSvwJukuVct370S5aGme/M7zNsxI7q+iNNUMcb
3L3G14m3x7zI8K/e/g6lxCt9uFTf/rj4vpjbKI6HxV3mzIpyERhyqC3w6QGKyYOL83kuVPr4xtPv
UGtCM1brtYS8xKiGGIyc2sO+mAZ52eNv+zWogdD1ofH6K0xrOtGxlii3K8hLyePI0Nq0stnuB5d9
s50jGz4BQMlBDfiDTZtpG2e35+SAza2bJQNgiHcmLxLAOJFve2JIED4u63FaRcOY4gTRWDHQATdY
dn/jGB1WVmqlv9eTTMfqxSTOnkFynCNBc3xkVHNL8jqZzzs9BidsXll1TW6RJHokd8Ii7eeJcd0Z
+4y7ZyN3oJ0+CooURweOEtTB2jn/1Rfpejbxq+4mQMIdAYCKpo3fwjDF4F2o/I3aIaCAfhE1GmpB
wn4jE+JQXB+N4+ty97jMl2bKSeSVwiNtAsILus/5SDRVi/F91n7gRnylVja7JzuMjLy4s3tPtL9G
RiPwy28mQ56vXQC1b5d0kG72XxVqs3raWB42jVYjNjmUn85dyZ9vJ4v7MDY/0QznoxfNIBJACRgc
zgxY0qqsY4fOz+TuvLqDKPWsDBsw0PAmyMh82krd3Udbc3/tpRFibA4IXFrLHHT+dRmam4eal2RI
UQy3qIGKGz9ID7MeFO7MdyZ0Tf2ujxVtaiRQH3scwLyBXCc5oiYpiwTpV1OEnJYHGh1IOlC5rnZz
fic9U7fOOxTr0DfHXgUvMFunr+qg8baSlhbtv7YKXGv7QCI1P8QCEB2SIGOe4Bm5I2jCG9o97OVe
+BoAN2I2PuFqTeH1g0tZWaAvcLRc10oneZDzhQomZ0Qh5IAKsrvSxxKc9vNSf6AmXBKs/8u08Tsu
tl/4makg33GyaGaY+4UO6D6sKaJSwBgGo2ajDYd/RcVQeIABtVqXHLFi+YBJ0GAKXN1tVQ5pV4vY
yUHBvq5SrnfAnbdDIPlzqy8MJOmca2iT0ApvJRcEj8pPfUMHQALgE2qjakMO2J3s1q6WdIrr8L29
9+ZvHXVrud0ZiPDC61AIIJB2greV0RY/Wbi0ps2fBtVGyc11jiI3SmBE6wPZAhW4uRa5rDlYdAEB
gZfT1oJhy1gyxzqjy0JvvvS+9xl2dBMSoPHPVhISJrd3SDxw8g2GI3TlJyTT5CIGI8xvTDFvs6j9
1dJs5YOBtgJyRADPq3Y7/OGjth+9EYOUSPkUFCKELA7bViwAfl533cvhd/wUZk4jspNqAZty28Rp
cCIlS/kXZWz1p2XCExOjMpto+TFZjT1pNTUVr5RiFpIAB3fnQ+7cxRJTjHfydsROOXrBPwvlLHfz
6+p8pVyPK5dGuCsJ8LSMLtQtsIKOy8/RjkfS3mRGueLfU3nJiwa5Z0IhjLlXsSQf2Z0eudIt3HXC
lgWcaalZMac7p1IfKp9cbgaeCP2vJ+uG5j0jlBTMVueLhLcbUrQiSbsN6BJS9gCCoJPK9VuTB8dQ
q456f9yb6T8LyIZ0MggiRdXQG4G+FurtCwVCHTwcQozFCP3MQFV+BTKzkI2PEM++IMWfb3ylQs1X
ydVoBwwL8qY5KHgXyu7DSZz2+XqWiKWoFYMbHUKfbG3bv2FQ8MXpoAtdR7nOE7QNzEvwDGce2Dht
/8rTScu3q1trCKzjxDg4r4LL8IxkMaXv7+D/gIzBj4SZNCNGjackZXVzo2rSqXbvc5/WKrw6jCZN
vv7rBTfv4fYWn3BGfO5z+4Zwr4V5Sl+Kjc2oh+xWsxgDvawfQjTlMy8d0hACRCusK20ZXa/TNLIj
cd1F9GfvBdxyp1uZbPQDyd9e4pNf3KIYYO+973eMGrSV2Iq2PmPEF+GATSULXNewf/sDcpx4hNo3
BiMk0cHDiFrN4kK7QeN+Gb0cZH+3ok8DhbopmCmoAttBA4fjhqPYUg/+Zk4YpnNmpuUF/csPnlC0
dOeOIWL+FG+MeWrZwdTW5JR9pq9A0sc4jnPA77k3MrXzjgfqnSsglbHZKYro349C4Qf8tOzjf9FK
alXLmfqMiMX6K+P6sT8uCCjim/OrOsqv2WwMxnmcXDwyYxeQtTkEy5Xc+oXs52bFXtCwNYLYYtox
553HHxf3zdSgxTogwbx4jjR0kyFZHrvTl6Serz0UKWCvfIqVt4hTGBMhDzFQ04hll+V2HBs8fd6G
Ow211HBWf4iZypr1QEqPiNvPxjGL1w3fn3BLBlpJaClBk53aL+fz5yCgepQELF4T6RUr/md/DRIe
YAi3HuNh/Zvde5CcR1HsAJaPHnoO074vbJUz7DyB/Wyj05wBh6GSAAjALOeiXRJQOh/C8FV8tDmt
qX+Pn0d7Lz1ixZYLb/7kUMXAkIOsbg9yt9pClVagWAaDh/GvDgNuBMXG/nCZTD4+yj/ArpnxXAKB
JpKMByTqQngr9Rw2IfX7e4kBS0xrC4SMvyQ/Pwolr9zGS0Kv910basSXlH8KZ+WrPFLKu1LtGC18
j33opMeqhWMa1q3R9joteqiY5CBM5TqJiB8ZXIsz4nPtzVgmp5V5Iw3rY/aub8MsyuPE//xOCf0w
lis9ASQJkAyRS4ZWkIZzILHEwqw7l376oDHywX8lUDIKH3aSLTFVKRVr0LFkjvmuXbj/R6P+t412
HzaHSFgQmPotCnuD6xS00E2kmooDo9HlmjvtgJWM7v4DrVIQcZCgLsrgqkwEwIBqHtPQmK1mnxl+
3pb1LX9uTGdf5AJ02CMwo4IYSpzbHE3iTRanEv1gxsqnweDTHUFVa+3URmLVNALTJMBDCuxWcSAU
GERO+tisvvHIP8TnL2l16ZT8VnaSBbZztak36FS1Iq1RZM4lwlMvXrMNaZF0Zo4G18T23gSqMeL9
l/6Uub1V+q+ki/5r2IjZCNHowA2wpdWQx48u4xG5Eowwbx95U6hEn1SwW9VY0SRZFMUaM1dN5eIP
vSHvNd3sXchocPzZ8H5LGvGi98XVghaDF2DXcV6TBzBSgNgH/xnkvfAp8na8EUru6knTvGy21XQW
+890XbZjbFOXXCb4orSBsNW7iaFAhf0H1KL1NGkWjAtQmly08XePGm17ZQ//Yaol/k45/gKi7NFA
jTXjefkkbKh5SxpK1JXrbxKGSySw4yB7SoHJe9AzysOoYOOgjbRss9Wbdxu8II4e43yFxfLk2jjZ
t/xbBlEv1TAgac14Owqh0zKXqPjOx+4KckXpn/HWIICeKqdy4DGafuuQMq6AF6FIABt9lDKYHJTR
lqh8KWOpDtg3CT4/qkrJZLvHf+o/RCbM5Ys1kHxjzVXPRNjm4Ud5r+Crww0tichTvkn5uA5cSXHr
7ILZK1D3p0MeaEpiYPjyaGUppG2VRIs1/UPqwHr/OJP5H3UoNTj1alfZJTxUXiLTuqcKLok9zwmm
XCzktDJ2b5M/L7rOIKPWQi0xpRPmJGrPWv0ctaYaTGwgRIbBogkjjs0nFVAo0CCi8nVi7KRqA5PX
wbKCAqwOpFnTbvfk4DtBToYlNEtaL/UXLHSHf1Rzx6ecncNPVHK/pqbywm2xg6rAbSpqvhg8WUxC
jQVtmb1odez9nTzjemY8FBEsAkydeqUNtjW060+kNuOaSoPXudBflfyOB0tVFgk7cpBJLa8aqyBS
d0DR5lLqV9LvI8ZVkyhZah5oyOpes3Yxsz/JvB8LOD+/D09kwMHBfNOe1idrTqB9czFPgSJBn20I
ylUH8GiHjj0vs2zR9819mCuPwNEBW06weLAfWNICHPdDcWGCelCtu7h6/y8M9rYb9gncsAKkvVc1
G8YETsNYbL/MVu4duupOvdaRDVIqrq5lBft8JmSSqv2RbaxRAe3s+sONixM+9Ye+3MF5UmAf9/rB
XPUrrwH8nqXxik6RGVcL6+oI36A8FuVriYcqRrwPfcHg7N9hMJ27Gg9ZHZs7HP94vDDJGXDSfvUH
sPR3xE47zdIrsb80jqQ2wBx99OVvEaKCDMHUWOj+YW7HVKO3Oq2gYUviFL2qVED14+ZHGEh90wLA
nJFwjYwdI1SUYJWCeGU4jJGnr6indWuPTtHL4cptnVH6TcKsTx7+nqTYT9HtkFu4AugSQ9nWz3GM
+zq2+ySvG0TETTlTorQQ1/3PHtggsHb7Y6LOVU+8d+3OsNCp5Fvi1lF5FoEl5qegeVX2XTeaD/Yt
RSxzZplpkXBGJAVAa6U44cUpOKB0gG1WvVF7CRk5cddZRSjAqBiCehNaN84KV+R68XwH3zTnB5O/
VcUFAJ8mfHiwa/KrrfifTCB6MvPmIVRRDXC0PuTAp1f1hlNYQe5/YCzsDCNrm/GUZBInpX4cD+xM
0vEfcR9cHEbP5XXxFiFaf2KyyYdfChtjN7b8kjSaZ81/IS7P0m6mejDLIVFwsQAEQ0pfPP2SwujL
tLRPhVuOguJCvIGSBv7uKEtTJb6Uv9IhEmgyRnFL/jpFHt78lZ32xEJOGk7+lncx1qcvSnXdyg7d
mkFrLKNNwKtwiYanpc+Ld1KtfoYKA4BUJIs230S1QzpaZlwyd3Tuv5IR1u1ywQtguyVIuuGB7n+B
E/ne3IiqnMsOVQ7ePxPF9PfWcRhDvZ9loEsuMUxDMqg5iqcD3+9Mx3pKiwJYgekVgc+rNXtB4bMp
GizolvN24kK9FzxvcseVsDW7tevTs17FTMxNVtzLZSziyWfw+S+JsffMKVr1lOXK00A53bFDlFg3
0IhW5cHOi1syu4MrvINj0ok8GkE4UrnR59vaJ+yx4WwZNTNQvxKdSTjhtNPRK3ABf60DQjOF7p6/
osfRsCVKmyb+Z2KWyZ/Or08NI9vfn3FDE3chZFaQ7nXMj/T8jz8+3UHRUqIRHUiMGXpJwyevmz6h
lYt+EqC8XxWOAq9ga6E5iCT1ghGJP0d8XF22F96dowgq/3K+0RfjgsTaOyRObNkQ7mFCb67oGfHC
0Zv97Y3FbWfViq2SXngMTf7+MTK+eClivQ527WGcLacI40pbQxo0Ackar0l+96hpOwc4KLCQ/tIA
GT0V6AhMNpiz5XGL+KbKSKJ0Mi3Bz4QS3Ny6uYVKrPjXN2ISoREZsRrY2SkkHVM9Zj/qtcGFX9r8
hld7rVQaLuYm/8gG9ihEEswo5m1A6ZDSdHDNv8Kl8rRKadES/6w1k78FF2oVkHQtCHrl93L7nfmO
DqoGaETvu6+PmsayYRhfASNT89MScPKAT9T1LBHaHgA7fyCR1P52kioVtqjdSHBFuAjl4o8Uu2qd
XEqnjUyTMeImgjZAUJBNLq962SFgFuOOX61qn1wWfS03+QI3f9GHKFPhFydAjAm3rg4TsPLwK7pZ
YU4AxHbiPCHewK8iuM4v30idJEwYTxYzFJiU4GQk+5h23zKcYKGxhu33biVPV+9NB3jkk5PFv2RL
meAMfmztQRaJX5emHVvYv9PTCl1hP0ugX0cNLy6w0AsKI5zk1PGhkyz6FHDFmnUTY9bbVDMALcmU
ZJd73R42eIEjuheBow0hiOGsi4LwO9qiFBW/IXHczZ776/w9cW0J/DWwY0OBW6P1lonHYN/3Nkvx
rxHuiYnW1Pp/3hn9ZwScRI0KrGxQqnZrh8OjiL5QSjsbeS6/Jdz4oiSXCcnrplJW6PLNKbliwhZt
j328L/GjkeqJBDcwIghR6/rwdY87GK+ITTtggqsJVxdGabj7qbUZjTpNX8vjO3NI1In3v0FBLkH7
6oe0IWTElFRoTf/5OK2w09ILd7yHmKnvyJw+tKQIk8OQo1tUImJgwMvucES+Usi+Em7N5ivN7axr
xY4iRa1YK25i0fNwFTHetZ60UabaMpZB95PYUVbiNFvF1z3420iuAOO8+lm8xkcoI91aVrMHJ1sy
LfaPaPFkm8VIhlP/VxSWTLJ+EoekWmnkvZ6pOrl5M9L8rj4XSRufKTl4rbnN+rNqQROGfVLK/t9R
TeP/XZUbnhMk2+rTJudqOUx0hGHKSuXCfRJxfP5uprH2lP7V5t+JwNnJ6e9LYsx095KhbtZeRIcw
Ggp8aX8HlaD0aa42AYXz6/5JBEzV+1f5o/geBcoT1Er8TIn0AHAhtDFdXZZhkdVuuQifA8f0+Fdt
dOq5MU6nE/jC18EJVAl26hy4PDJ+1E4UUKWumPnRYnG2LxdMlr/vRmMsk9G8HYs3vIYgeSbw4FbQ
mseB18Yvt3bFJ7WrXwls8dRGYYQK0gcNmlQ+QQbRQo9TJUcmSmRp7ATCIhfOfVR/cN5nDn0OqXt5
Se3j6BvNrb/n81xQkZJ/OeLCMss5CYHZo2IW1pV321xWvtxFUB1nxkpZECSIS1q4ITT9wi/fcnNf
lhYEA8E+VTZeboX5zj/f2HpUZO/s8vG3dK0sHzy3GUMYVb6Zq1jzwLLQvXsV5DO8W2Q5KU44HjGK
FmNbI3qf2jQ9YBHWC4BM/HLcYxYTNSSSqPAfgcX9FUrj/QRMLt6kOs8G+2+eBeCLHFja3nKdnXis
fygZdkyhCs6T9gsekI0NCNLb7dFm5J+UVX9O0T7GBiUUZU5JaztzDAOwDBvmBEhQlSCnYn7Hwrud
1rwdW2SUOhX8TFDqCz8yzJ64MjUBxa5iX/+bQ8e/Kh2XL3WnZSzrnaiqwAvBvvGXPCPAQpWfyMkE
fY0ISUO12kltPrTlXA2qL6FzW1xYXSKtvUD24P3KF/ol9G3nXoVMfdNWnlWfubBLHalERDwvXqOe
LhH3mf4KCNe2eozKa2oMxPOxE2rpH+xrBzVzzwtyVd6PpCGt54YGScBSiv6JTsxHzgPxjqBeo3+Y
PX1QD1wHcg8cwdIQjVUYhZNDK37OiaUGHGQFuZ5KOHxqTloXyKvTuTjDAXmlqAAMWRM1gLiip5nX
D59BZnD0v0J7nP7uG6U78YvynWIaRQibYtJ081OwlfT6j8d//fDo1aUw/onJivC6bgQjfuK172mn
pwbGo4H7uCBI3i0pv9Nu9DHaiowt+TLOQwg/PQlFufW+z9Y/TH8oSrCfADZefmDT+PSiDIXp4yrn
/8tDz2Ec5BnD6ombm7fEVRc6qDKBzTY7NLwkT+MT5yv66ZcUI56JssRaT/fcRoIzoRszpkOn54VA
XTmKrBszaPezZwkFMRgFAEO+JcfryOhN1cuUiknBOWdJqA1FO1WiBpiBEEBJ4KrPbx1BEwaxVV6D
coaPL3X9BNn9YzeMtUR+6FUYWX/noyZVFUv5kloPa785TRERHe8H/qaIR1/xyVzxytWNK87Qh8q6
2N3LPe2IjfGT/yADeMSJY+TCaVNIjkN1YQHkvMXq2YGqwnNZYCRAoHMB51zr6ly/mvjPcnqm1Y3C
uh+qWwsUVg+jZaFb0v2Ar91enj6maW95ympM4mu8bSdQVqwN+LXxQcHJLPs2WuRpabAFrq5IE07T
lMWOGPNvIwg7nV8vdXXawf0DrqR7H/5xmx/6CQ8IVEOgGyht+MUb9IZvI70s2FU4g86xgzQwM97e
3I0qaxboe1HMRHmpAHfDmaiOhKsOv83kvRbQbii16Rz6tdmVGvAfgd1YJf+gyXEbA79tCAfUlvZE
aoO6BcgdIi7rG1plE+BdzLwb3+IwAuGqBlObSy4/VmgEwyX0SLdeginweTqS0viv3bjdZM94n1nq
ZFqpwJSZTHWoE8t8woXqzlGV4a9PMu5apzTNVPl8O5LEaTRNCS33+1CCeCMpSs6yJPCa7IebXZ/f
SwADmaT8RqhWuduqW5flt2Nlh3AST2cTqBQrbvmD7sOAZBkaCGcRMWP2ibjKMrcNIL7nG0F+SBui
rVHsXLaBpK4S5vcNX+hPVGpYxk+ITZdd91sjaSQITsHUP9LVeKoOl/CUA4kKGY39aVFcffO+Tb3M
tZLOAzx9UMMq2y8tHMEtECqzfmFSPUwAq0Igay68xH01ng40jd63dohSEJf9bOSM6RLpcofFeBMn
ekOktqOCryKIOWLEN0SGFtxY5XMrMQ7t4E/vn08byc+dB93IAtplopdWMEfbKzxYV6zEi1raxvvR
i+jqfqSsUgX5Fvq5MCapDcg7H/vnWZBgSyxgC3FjPZzlAZeFUDmhDChHCdjAYVaF1uBgeT9xjQS1
49vWmUrzURTZii4kgyHrkvJLQc3NMoqlT9Q2u9rcM9iKPjNE2dqUxqb3duoZxZDSkuRJG8/aana1
o4yPizRTffP1d3h9lWnexnOsTzFS80oGSoh95RurVwBm8ven4yJ6Y++8/2BN6JOykB8x0mPNTEO9
cmXS4EgacKxLOZ0wYFC9Iwy/BcB+HTJQQMGlxCYU5ItqBaLCe/uubAue1tUE1XkTTfDUSlB9jARi
TotL4X3/8IXirK7G3VsNOQhG/3JWJ5JMxpHEvVyPbwhdX9M5VwBhrdBECyLKRYi0cw7rX55TOrqG
+sGv7qYlIC/E23lfONsfqnvQxzc0ZcRh3xBN2vZRJJ6sEfPxeq4hdISSCMyn8eSVdi2/TytuRrwL
N4TmKz02m3GowmJpQc6ldLPwxBFLDCbqPFEMU+//9VYtWZrFPL9h2g81YVmGAWuATtj5fbN96xvJ
yKQajnDPqjeGXqbLh/B0Yyn0t7J9Vd9RxV/zj69v9vVeg9HZEHmbPaURpmkRRC83NzGZwIMhFbAn
38eX2T6Se6GEXwyw/qrCw19y4ITT2kG/vkYu4V8BvY9+0gb7hAwafEQ6rBKqTXUCIEHBFA9BloY/
igrLg7xb97RONq9Eac6S9H6+WDMZHHOua4JMVQ7kssHlw2JNqMOZn8N6/rTIwJXUnXE0obS8FVrp
qPj44Qibb0WiSGGkqtB8uwfJHd81wqcicvW+g/2Y8DIVSRIjhirC38+YPdoeoRNM/vfyPq1WbGcK
a7URvTWbDbSAxO7vywY3F0rrSOh45AYe3te1+LlLNs2UfSDuDmO/xrADAiUBtJSHKhWuN2/RmBbF
8/EcF03gcxm05IUUtMnChldf2nA0qc5mk42jULODIuHabhpbBKWxUpvsSb4hkShGh17JGRZxNYzR
TD0bLhyJn6XylT9beAEuMy2C7r0lTjKpgjcUXT0OloTeQcPydU/FTi+X2SGywoIKb1SlT7rsjRwB
jKCh/OxCl0pYY2r96Ed9WoNTbKYaLTl0lccgRHtUMI3AK6BL277j1D225fBhR95OhXq5ATM09Bb9
K+7Gqb1LLfrtgejuNTHFYOMw1guYtryBrGxpQ7ZOxxsQTp7NpJgdG9uKPMZW5Fb6xF1SHy52WPEH
lqFyA3TlgzqMfhuYrIF17K8wnt96cCyZ1DMWttwV2sTEacIQasup2TWb9n/SH0VwkdwqpPPMvQSv
dN5EN8OvfC0YlN2NN1kDCoBKR8Mooins10BJ2DbKMtKN0NkJ06oEIxj/SvgZ38VO9z8nbzxZb/io
X8uxqxjkW/9eIszCq7EQZhL6VLrNiaNz+JP4iFhNzBGlVYrRYqRedqkXnLad6T3qFDrTl85dXc+a
dnBu3JnSBLqpsCvDvHR651UmH+3YKdFzJn3n9KUeXy6MQUqRtE8bHVN0aftpEtz6tGYs4txCieCR
xjvhrYu0CgfIGshuADaXcl07ndb44QiBUUuhrjBpgDigeYKRWcpIuh9rttCRNBdjG4wO0I9ftbY2
fwXBdkkH+p5NJxrdYOTrXm19S1hpIO40NAkyZjLQfeUMy51tZyCT6pmcOXxXwujNFfECN9Y0GRQL
QW4+eO5meZLe4uw3vbyJI+XaKFBdB93BwEyIXc3grLONTjaUbFTU7+u4IyxEGmzk1F+2QkyxodvY
Crotrl2fmBxBrOexDncKP1+wyOcxP7C+sVwRxKdHTZxBU1oj0T5UyGU4mE79PYackwhSF+olH6xl
4TaypIZVIIeKfMe3MhKPyceap7JKweHeOQM1SaRNmLtScm4Wvv+kTrInwBwb/vjZhWodZSIvVQoT
kTUHsEq+vFE2feu8XKi/bMye8YBcuwIyWZeG1d3wPDqFPuMhdzPMENcRKH5/Cbr2AR/4fJRvOyaY
yQcoVtXUXQN1lyxvYrt7chnrB8gFeQUNQ1Bvd0LMt4AZ9/6ZnF17tamSRRSoE1Gy75WfSLQg0E8+
io+dF1Txud64caK85h/IZEfERlcRK0OEs079D7rqFDr7G9OS+tJyvbZnAa9eLWE9CqJSCe96xbwd
dIL+jPKUgkIVh9CtrhwZPdpxe9jAqh42rGQqs3GiSOK3c3xA18fX0IZcZyMBr7rHxxvqh371GSPE
3zfjpp2S0fPoJ5g9liMEupjaaICtVVlJEV12uPlcfRLbZqOC2mj4v0IyBnJIIEgmeaG/zthDGRWR
H8rA1xwWjtd092MnPKANRRS6VUSOoIa4DYYZrvqrNURlzgGElSn+fMjgYUAv2QEH3aCzUO+w1S0i
Oi7jd975/cur5XY2U9ZJXy/i6L09xdSQ4tF+1dt+niSEprYEq/Q/xjvmiqT/Ap4n8+/hSH4x90GY
SdB1wBjR1RlS7UjeLMsJmjvcwoc7Mdupt7ltIvsio7lwhljDqm8StBUb8+IIFUvCLk5519xDGwDW
Btd4VeXqDJDX7J5Va0Y2Lzz6pTy5YxcGZc1hrMN2CRoIXfdAFVao6wzCZrwZYR1LYmfzOB/RXedr
9NpuwjDjO2YEjY9Wv/XllsmirCG0/IwCa12oxHvcbYI7qV4y5Vy/aDLCKB756q+FZiB/R+sz6izA
Te9FjAnH8zWW1nz6/upSNS+rfbpm2ao003xNZ84wIbH3XLHXvz43cMfCCFH2j/fFMaatJ0Lq0Gu6
mlTKopIZ9s3uVkuorT6dUAAmdhyAbOqBVU2FMp2wwrKtOmRMGGIswAWA0555WlC0GqG+aKv5Hkm2
x5P5tR/1Css3D2pXE7GpJplOK+U5axu11EWGLGHyKnRna9S8FbC1AxScDmeU+gKNXKx81MLmf3q0
ZFbDBoWlefb6pCnpOohKTvvm721WWc4w+Bn0aBn5HXwKgw3fj3KBUXZDHlhP4m+kaFBGwbFmi6Y9
NL9xM/ArP1VdP1H7uF8wGS/C0TKwA1i5EXLYT7qwmkTCKYitTPxOzUIi84Agmt18HmTEiDkPsz4n
jodrQ18EaLX3tAUPrmlC94XL1kHYs/4fGfOwOuLVdBa28zlJ8yvpaT5gq8oZtMOm6xghjFrkW9DV
0NQrHjW/A34BDNL0TGDzYHkV9xL7QK6hNB0MTtqBNmaTzI81TN1Z3YvyHP1T85abpfKn2sAi7HwM
rXhdvXRvNr6DI9yn/I4z87K2IVWAlKhAgtpW8Jsm7c9QhKBGYhcqzWC+/DTjC88GmGDJKbCPQgDV
6w2guHCP6OZXevdx7r86F7RC4p0jvgx+jrYGbiGvAjzr7Opas4nnFLX8N3ABBFlpxYGDeRmnZOOI
jUBrcAYtsNwJf+qGhz8OyBhX7JoeThUZJSiefnEvM0mgQ/TsE6lgdCitgU/pjP6Z3J84BqpSc/jR
d4SvNQvAFycbj0ycGQHMf1V38xzYhy7JDDPEt67rkx7HNlk8Noql4XzHUYFdvydI/nhlhlGNGiya
lrPuldDrb5oYjsy3xOabnpjjv3kbqz8jcl6a5b665BKPx9EaMWXOBmk+ikhabIL9MCShDIxUvnyE
Lk38DkuTpFaRh+owiFY/Otu+OQ3ZiueItF5JNqp+GOHNVbJZM55eaGih0eQ9I8hz14xJWEk+y+KM
uSmXM27SAhowtwl82Vj7xxiZ3uYQWCGPJ6YtANneVy/EWoUk/HE6y94mjrEq6FVa9YACL9c6SSOk
peU/79I9SmQXx/V2G8k+bYIFVg0iRlORLy7HBX4aKCrudIEy97sDFEo5WyNBWu9fpCZHtk88lTcD
KWviO/jAzvxuyI9kcP5UMuka/wZUx0p/o+A3TB6ZQfOaDiEU19FEE8nf7HpOWHJaTIXEmAbNoAgb
BwH1XOzBeZEtM+14pFVisqGEUceiolIm0+EXaBZROj0wZmTIRdYkZtpvnhaOA26aSNKdHVwD+v0S
9mv3OEXkm6iTm+Dte9hlq2KM0eSDim+wWWYi+yhridtVdbo9Ae4NH3avsF15FsjLlOkVry1+wpPi
XKfiYrQLzZdmOqnfa65PiTOCFeLzue/gbs4uHPX1UErDVA/jLQZ86Sy2otpyb7sBRN9HrGpvxjAH
6FOUzGqiyRctY6t8W+/z04rGwIdXpoh1f1rGbMXQ6V290AtYCCnelofPqzCaBgSgzZeijGSnOEQf
ZjwqB00sHaxjS+MV2Wu5S26ZC+GtevIbUh+nwpIkLbQmF8huxAc35jI6tBfXiukggFDWLGe66f5D
xh59z/v9JHR1hhWh0kNFHmR5P9beq+zMJNQ04OxlScUuDCsbGc1cnP5DY0fcUYDb01tKu1GlrJiU
a+ypN6wxPHdmWnkaKTiUmAQpwPxCmTzmXFzk4hlH+BeegNtu6Upmv17C+s9qt78rBSOhO/Lr8LL4
SAHmKjSL0d7Ba/nnZ2tEpQ6d12vFQjv9zrDRI0kMKsIH7ep4hj4AtEDVa/69lw/VQsFQrt+Zjtku
P04NbAyYQMceHjruLxIJ/HTTVaYsSNMe4LT6G5bI9D+z7hEuuDb1mHObTaUYreMRlk5avzOAU9x6
qzFpTbKZDgheaiSKP1sJVh1mQVwag8liQ+5Wy9nasyWnq5O/OD0mWq8XFGw5U3xdqm5yF5pay7rR
0ZqerWS6h3wHpzRee0jPba8PHkwNoodKgM9fwwODZ9f4+HxhBQBKnWk6a1bPE4NNDqf1GcepM4eK
HJSPhemLVxgzQW5u3c9DgxgUJ3t8UCAtdw443KsaYzZfvpqtCrZEl+IHrdBmATQyY72iQgv4x3KO
i1waG+cxkwh1foTjaHJP9n6ZVgpYUOkeQQnYj/RfUrw+kuuVTrmiKC1olLdOFB52XLpaqWlT/Vq9
MjyvW0jRerjNcgrDCjhl2i+KFDVZHZJ4LpabiPEo6QG/+1BkEeVYyo2SGC/ZFRHFY4m1IUovTACB
G2eNFqsgGeY1G7GQPP4NOpfvxgeJAYnQldcgBblQaAkdOBT1lZn++7qmGE72DxLB/ynwXlJmyflk
Vwi8nViHMdO2NRJb3bx2oDEdnketSgdynSO7x2P5IpEi2FLpFvmtNCp7mzLXJbQ74z2ovBiRleSK
BEcYLuvAgn/nNKgHiMezuoSuatEEZ5QrKvZsyZyrPJBTxJ/B+Ie6ENvNePd02qzsKA/ibJk6vMI8
s8bop0+WHrB5JltrGNui2wzEGATNCYIxLBThul7sw6Z4wcuwomCXTCgrUQhsQbDpmcpfKoPhOY02
UICifQ+/MyvxiukSmWAid13SPLxqKkThBYnPmUs2Kb3KFY6k6aIPaNoGP4WtCGwi5h1iqeVotVE6
D7HQ2ZPe3SS9Ij/srZkBz5nMHouFGy8M/vLa4qvst8U11XbfRLkyjAT76r6XJ55mY1lRESz/W/I8
IGGzi/lfd8TByiBHd7c3yqXfDqDiCLLgt0VGgatI/b9VR5ceEFgdOfiLw4Lzow9d3OFtZimiUZsf
Jx9qMpGu4L9/r8q1sWQ3KS1MURJyuzXCWrAf2HTCaXpx0Tq6C8wYiAA5NE7X7IJOM27lNqHUxm9I
Ul2Rb1sgHcyEE2Ob0JETQyV+9NjAUtlZ0ebtJ/p8HzJYQHd+uHwV++SeJofQiwXJ6NsVVVMk2f6D
lLQFfeelPZAmHQPmZ23NTNN0NEGZQmzTHw01Z0t2wlID0NWstC64C/oIeqCTQAaIE8jLa8oJe/5e
lWz1Zl//U4d0IK66KSxtnORJIiCDgkul79mK9fM+HojRcG/mSZqRvCvqkxANYLknlYeGWWsh4+Np
70dpDUT6k1gKV32e6Wj/h0byyRRRPhmnMX03LEuSpBCBm4M5lKuFBV2D4ckbXZ9F0/ixVTqhObPD
Ua5SnzMjboWVZOCNhay3KkhjF/1zJwE5ioNp72Fao0cM8HJ3PQ9IFoXYWiMckATVm0RXOTF2XEmR
c86RUzGHE/yNv1ggl+8dINJJTYlRvUgy1YETceVuABr38lrfViqH5sx55XLNzWHtvSgypdQxb3r9
kk0v1mUk51ZUJZ3YmBLBPgQ8rsnSl+5fwkoUWFmdX4JvLMzne3JAyi/XbQYr1ed1PXje8Ssh1N/d
BkS/tAMdv5mH6HHdo4gU4JUybHsvL3a3KA/EIyINic9G/DOjavgW9lFK2BIFnN8f/iQxkNvwvgvO
k1inTLYSyisi6K1dCRBbr4RwFcXC67EO/nGX+i0XU9UF5bi6kOU6XwOYvb1tcqNTjLUNDR1Vez4u
P5esS4KcjDf07SdVJKZJiTfq0wl7M1ZhcEAYK/zL0GLToJz5MUQF7ZcdAHulpsXzFulI+1cZZDsy
402/+O8OeCyTiuXKYj/1PrAfX6QDVkGncWd+Fu6bq08n+y88Yfc3z0v+brX20Ykm7nEUSOqH6bxz
miwFuqwF21Cq1G38ExpirxAfB9PadXOCK9fUoqEGsq75NSjuOv60VvH0ko0M+jgEOwvCc4Gm9UlQ
d4FRXXeHpoK7z9TrFy8clsJ3SLZ2kl6Fp02HUDSUYSMnYfYY8safUVBR9K/bhSzIMtScxXJZzwDn
L8MZlHV+JKpn3oydPuqah/OpHKMDlmRaqvkkKIbQ2BnlqXRNyr5pqqRyy68loFFGA+2mwveXyNtA
pWIYO0nIqpsQ+EcJZMfj7sPic2lAr6n0G+YVjYIQWdUJGCtgw49GqSpEA/ZPN3MtNwOcbJLcifL9
MtIOss5tOZkhmgg8Y391CZ/H/YKzo27k/9M07fSY0HDB3WzwFawXNPwO0GdqgoRHMnwt5/G7x5U8
uLLDJcehXZYaAC1wySmTXz+oHqSBJZIRrhQE4YTyUdvdxQFegtYzft3LVAiFK14Uy7/omYQcwFS3
27ONi9IOkmwB67uG6fKfbNvrY0W0zPhgZKTqLrn+wBi08uiA+0Mn0iolnO1EKPYeEqjZx3t+cYZI
lglwc9yQHEd/BmUDUcFi/EO5Tds4BYqhFL1JsWeEs2UNQFX0fzEWXhq8oaSuoamhwjjBekan/9A1
Jn+P23OeKmFxo4Ifm4LgEzKkrIyAnJlUuiMxoec7U4JEH/KBM2i17lK99LNdv3fGu9Gr3CilIAmP
TA/ykm2J4ObNJo5A1rIR3WanhcARFveqY5ikCqtIX5G4LIeP8jXtvvK425+M6B/nHyFdtvB8l+QO
YVKJa6+IXZf/qU6P7ZmTDMAtT2tmBXcSTHBteijpiKtuZFgU+0lEFftn25e7H6tDX7hfJ4nJDi7x
W/AQ/WPOCLdBzTzK1YHdfXcrHTy36K6PsC5bWWItkd2a+FdKOLgJFe6qhbRndJjbV7isxQy0qS0i
88rNynV+9wCN7swvAdjMWJiVTBi6MUMKr6SiPXFizeHprhYmTbSYPCxKzgLsPWZ9FwkYnZHfxKEJ
FlvSdnlt1tceiTCXb1QUcjrd+k/uWDmsaZMjTxzYKWL0bqbiU7YYgdzyxh/AtJvSOf7lhrBqrEdU
2Iu7kA/jtIGOrWFo5nfe2e5DfghbbgZTZ1/Oeq0xiRhj07hx/DSUsnzk7JbZ6l0WzqfGE7uFU78c
tUi0xF1Wvmy27uegD+0tzX/54cRFraeO7p77RWdtKnDMosxRcjbo3Yc1tTnV9TGv9WOlElLW//8A
/tavLfqwRH47H07tiAemtJXe9G2QX+hMdLw8yTLcuhbDLeUkSj+3FJX8d194G4va/fAanbREgTaP
bWuGmB/UgdsxMVaf1fGKKtS0HrTFq2gQOGj6zKKlQQiZx4MGzFE545VwBhZW+pQ1/6RcxDXAEzQB
a8JjonNvOb0ReLHtmABdz8ykbr3/TiGVx3TqgnNz16QdmQH9e83tYUlGenS6NE1nYGIECZcKqtqS
F6yHxWNV0hiyutqdZ+UvRHjzknjuSAsmwTtOhw3kvwugNuWqBGpD5k3kfRdK93B7IPU4JmmS6RuF
vE6u62YgQTvCz6F3JXc3H5/CH+36ZKjWnq499DvWMOmX6hFuXp6KRFPDWinl30ZfHG8BN7C1Ppbl
4gwfi0bmSahvOVdN8y+uQKFcCp7VbuFVKtYY9mY3EY/g03JtXrU0dfok5S2+XY0egtl0DzQnqIHv
kyyN6NmHr8POAay9UigQ4hpbqmkDJX+hMdKISogqiaBPmthChWOh177zC/egRuCLqqCnEZT6LP2z
0VWrYpi+eHRwaXtgsREwUgWG2HZqw/5UcOqVpjIfkUPdAmkTw9ygXkdfGBe9eW8dffQ0DRP5w4Iq
g7IPgTxkegK8ap1wRP0L9F0+hQNabGmSLXlhGbn7g/DQOgXIkylc1NLAuDhjuI0bfmQtovQiIaJR
1bHVoF99Y0+0UD6UPd/RYk7nBp3XBLNFKX712t+rXs3+NNgNmDUNct+PGpj8LtPVHMf8KEqHZa17
0WEAeU5T+soqkX6TcxaVGMXzv/solcm1ryZuRxz6X2gGnAgstwKxYUroRDrjLft80aA0Bsj4ft90
aSRhrfSd5HoHxufk9ifdPuc87zeBKpi7gWjfN/L7U+zbxCDkEz0FbB3TgNlqGsj944+vHd3KRZPG
k02zKO4mdEDr3XeKNE+/S9POr/8hLWR2tEJGxAtWM6SAEbo1G6PvM7mUvyllkNUDXF5MHjM8ZC11
qH2KQmJ7OOqAQlmyDU8pJ5xLDHZUH6Dlm4RhNyriuZ+l2COYlIgrBNztcBMo1+JXh1tZJEN7NR4B
zYzQRn+9mX8tmKByfa6+tjzeJk62KpRsHZzY/13EVhm7DTH1FQ91diz1ALayaS0z9LTiBSoEISDD
d8b44F6tEgNDn+QDZ1vGTLNkDnT4y3kNbYaPh/LwE9cNuazakka8K4SOHwTUFSDcQSfQ4YYkUZ6X
HbfnHvvvN7iCwAOCLr5AduWhI8y8dMc/kOvMgwQUTP21swlqGHLMHjcsrYXhkDWCBQ/cd7PedxIO
qi5R1YDmrceKRwVpc8QyTklPnoPDCUPyW7CXukNkak7Eq8BC4BathhSax6CullvFvpTHsOlNcKhx
wOSI82GCKBIrEjlTosPHp/CiAL/YTEBSa+sfVifADZgJCKFSLMehhd5OESu23VqCLdS/LQkcAjfN
xLKLAoJ0n+capDfSIXPqBpt+FVbWz+PIxl2sbptVB6oIfgZxY3CsPdyDu/lb9TUIEwQpjudxJ6Am
hH0fATkeSqpEQSvfxhM6xQZ1xA3q06KVYVnSBKDa04UGgnfJGB1bbKLja/A6vsXLBgXKnFXtSKAv
4/ewipikNNdTBOGYSnmH1QKe8urogzkGiUjNRFBDzZLx/q6ZXxZyf+PSZ5hg6BYxi/8m0O+Tub+7
DOZWBJ2Pi8x/DoYcb43scaecAFWMPZquluX0WKNnl+CkkTvcYtBS5gh1Tm5mQA8izgu/DSktbD82
6vl9Fn0NsYade1R5MQS/4uxz7L+z9Pb2Zy2x5+lISJrLPykK6ThQOtQjbbu3IOI+g9M9WIXzdEqW
c/9nEuTYq0CBItBXXpN4YBbDxJ70Q8fZv7mQo4RlUReSBOnfZUBNYZS5wuBXPiCJRztnyRaYweZu
NBmvMtex3ZeQSKNtBVwyMnvBE3Q2EF+nfdRsTxFoTeD2vCQgY+uaDMhoDz7eovfDsUknklh+/al5
5fzvo9UQjzdtbwBE7NUf8IYf63ZYf8y+H+fwPzyuHyGMfgtdfL3Tt+Kfo4PuhkmqF4JyfCDNB9d8
DzxJ2SkDNZeUjXHxCajVhSDWVPqCGQgu13/lP1S41Z9+EKUOb/SGwdY/oEQzOleEEm4TLNoaBiY4
8fz3NbPVg3PnsfenqP1jFBCXG7N4ZubQcPM5D0/4mGcndon5KxDEtJZDNOYB1EnnQWWRlEXwZfOW
83fuvozWe8/h0ACNhEvUyZ3L5n4yOwDCAdxI4tLAvoGBK1GL4b6alYvd5bBTHmFq/XlAGnQYeZHk
zFsKenWYhv3+kCVvVqxO3IO6E7u52hYAvLckGS9IyaNjM+ORDEUrK6n/zppxHSomHvteXULmHo/W
ccbwqc2seiZHNhnh82RlHIxnseyV2sBB986mA84nKibxmQrmxHQrodq3gxcY75VRn1AG1OmCCFqO
0THmHmwmHNke4AhCa7ZBHxMnZtpxPyk/PnUG3xDn/BmBkSgYgd1I67Vl5Z9R1UN3r6zEU0bcKuZP
zdeH9BVNXnNxu3qV/zxTicdy3Zcp6ijGOshHteaZqrEYWZd2xLhaNsQr4POlawxIiQ6MiBHMXa8N
xhj9mZEDkIQwct3j/VSZ6cShbTGgV7nWhOhsAl42su6wJcCB9so1KP3r25kEk1MBqZt1qoa0PnZv
LTtWhom+W/f83eAPrQF9xxLnh5tkAt2m5GC7MyeNQsrvn6NSDaTFPXiFvEGCah5iQSPaoSnr1XBq
LxZ1s79evut592FXUSaGumFNaXKNRSm8CBybXl/Sl4r4dv/XYsCYTQ3LObvb5l1iAJzIo3JobBL6
CH10gkr0p/QuavLiSNjh/mZlQYhXCTPiKcVBpxjPLs0BEKgn2EVw1VGW2k5OO/Ce/kCAUQ9AYwRa
a7TWWGycga1fSyn7G/jHUxa10a4Vw+5RwNX7MxqEPo1KYMTfNH1KI/u4bi+s7h+duJDAXC4QKRyL
Krfiu9idPMcSbBVj/rSiSn40jPFhoYlOoiKy0nEsJCMXAjTdHvx9TVpc/lFoaq7n4QZK9V66578R
ifKhD3XFstT252jKrvFdDkuGljQRTcJMDEzOf4Zt5BCy0FWuND4OC3nT+8aWvr4NP1ds6nnJDjVo
nQJn4prhYr0667q//rn/G1JqxKrBNjeZ6WXO/pwp2dVwv41cXq4fsK+BDFpm5cM236616Jqmliri
xDCzw8wiF3mzb2xoEe0Yt8IFGtg9M00afo8uPO+isUkjCni6pmw7yj8UXphs4p7TtmW+QTWaa+hU
X7sbrt706v9rjYkwRlzRrfdwswrZ0cn14Kt2RT5Yp5GWKHj7JdjUvEKgvDS3vNBYKnzb+tyN2uKL
aOtGco6rBqxFIgDaQH1oekP6bMYllKodsSJcT/mbd1gJ4J6KgIBaIEHNdpVM2znOhPkVTaiijeKN
Z+eYj3QVIoP5e3eJxs2fvZ95U47Wy5L64ZxawrRuWzx3rXDsb3j9Qz2bN3SWm8IGWcMFxVwdXOUh
m1/RuelJFLZhROoxV2XYBwEgd01CvGGiO7l9LuWN2ZDc8NZIS65C9KqcUJPgEpueJFjyavzqoo4J
HMht20gFgYr3vHny5vCRKGjoMCcdM261YjDnileyXCre5SiuIOgAUpJux8d2h2ui3NHzDKIOFo3q
C5JxD33YYQuTa0lDih0wPuVpl47EVytF5mAtFDF6JAES0kPzwHvmVbzAj7qk1hml39dHX5hmzjyQ
zYTuHL/U3hH9KEkFCoSrgOYIDmIUqaELbIhseoTNQMAn/yQnu2/KSFwXCDqtZLmCSesemsH2lXuW
QaDC3F28NM/zJwzY0jFu8G9HNKwlWPVLlEh711BVcg00MZVyWsG/B2O2vRTxZHaB2CdNW7qeG6gr
gA3vffU9tG5ayTedvuL58+3CJF2yA+Iky65faBalyRqM2aUlFZgHRqp0jeyXF7RYILasN4a4AfIA
RM3kguCvBBdKhnEKZ3zQMB9QLfppKo4G0KrhCfRA+L3rD/YOMWiBycmYUzMenJl/jSe12n3U6k5h
IxnHvH0CFlJFSm7J9oPldzOTmhGTac5HI2Qe/HyZ7lFBMqMVy0t8GthIJ4B8lmD7roCOopd2gB3W
CJntwZj/irgL5pSArpIaJGc9A4JWDu3TjGe2Vq5Zuw6xnqWLEqE58x7t5pVDIhR+3uFaRxirkx9U
L3Q7ZmMcV0hcXCG+pOFzofwEPOmG45nHXzoztz+9TAKOPe16ehxeK4Do4Hyr25PY++XCe7m3gq/u
GUzcKo268GKy7mPnd1uqP6sCMicVad7U80p90E+w8G8n/fLe9pNbAxdeIUT05P24T58hLQUIYQ+4
OGRZlOHqg+84tdWrB3ldIOY5sw57Yr9KeWQBo9GsRBwpOPt5DVRXYY4XvtMPslYX29oF4HqkKXzU
1jBb0Gq6QNxsLWu/uv3JmK285IUAfY0hpYVbpNPlLLZtFR11LpuCcWmTHHTRK1CpHqHqdLZaoAIk
uFBNsbe8NjrnTJHzNmwkM93bZTKNokTDNQT6e6ku3x2W2Fk57IwaPUJy7MyZib1uiOe3ZA74n2xt
R7Y39YKPBN3eZk+HqriIWvW6hqrvl01cCPRzGcnvYGIOeEqm+C0c4rQWCIJpuMbi+KNbdFuXwWr3
VZg7SHn6LZDE5zA1XpBpubOE7FNcWpoKzomKkYpyY4zihA/H601aWQfAWNSEN5VleXiQ9Zb9Btcb
uuhPv883L3kei/qtg+pQOeREIIBr4zb/dNt1PH3fXh0t7mElpfj8CO31sxuhINSa8kSXRZjsiyOV
QMvSv7FVyE3Jl+OD/g31NWXmr1tLgsfC3AHle43FLCS0adeXZBgqHRqj9pGY8ApOcU1xhMmOGK19
yh6+twtdiccSCdjZNcOCCt+NyhtPrxb5kK3JPsmIHIHhAvytxU+twb1o3A26rfOQpFSpkMhv1e0U
D9ZUcP06iIQnFKL1FW4fx7TwzkloFx/Ma6nqUm3Hc1EACaTV37D635XO20rFRFVIq3sc+1I912XE
dHKZumF9Xi82PGwBapTlNS3KPARai3IS63HUeMyGVM4NkJb5mULAR1adKi7rSYU3Sb4WY0lg/EQ7
SYJ7Yyvzc+YEoDPE3wtlVd8Wo4YpEgimUiHOS2/LIfxl7Ozz3knFyiZLy0niAzSK/DckcL1vQwKj
oo7BwpWS9KZNzCfj4OVJrs4vesOUzN/9Maj6HNrr8vehiNg487nHaj+aQVY9jcRqsSLt2KYAipFC
LjtQUjczfivGt1SBFyjfTNTBrzN36pOHAllK5UGu0+T1oDw8Mlq0lRx5vve1FtosGjTJEpIFdPJ9
ZQcG7ncH1ePv9wNcsyobvF5ZguZldxJThJWgpvaN0v4XjxiaNO7dJ/QtKZtVflgyKfIOG8kOjQu3
zDC5w3GQRdxw0Z/H9+z5+gf+gNZIUvx2v/tTEUgU3U0Zuy7C9z3/i13YYCytv5ncTXJAVfR6k5Zo
/h143bHh/iRwmGmo69tQcA0OZtii15MyGpoLff6fKXjRwGZGgRwZZ9jJqDDNzbzMy28OnY1yE0lo
srMtLZG222O5rwwmDEaQEsWu2PRnhvswlZ5/UZQyKbSd3Tm4iIZhAoAQ7rTK8K63REJdSSrmjKIy
s/Oq8ZdxP1auI82s2FC0m4dKWPjtXauiQgXVrS3vAwE6iiK5dxybByodp/zuhq2MTavxnoK2uVPg
FQxJM8OjyZXSypEsy/yX5Pfndoh/VVuSwT6ClXKb3Y4luYWKsI9ZqGu0mixgFPlJtqHUUY0HGNk+
VcmCUTl68eTQoJdbNWlGO0XyICcBoFVl502yxfIY1z9qreq6ZnWBcaGMjsF76Sd+gND76Pf5U7wY
JCtrokn3PEvwh5pDdK1JvK/ZgVHCeEdL6gbSBFzAwGr8NWd8pq99Zob4mLFfXv0Rk9Fl4JOd3B/x
T3guh4KnI83EziBKbsU1vfNBLbz+Cjx3dhCBzrTI+RaDsqhcCLsWuhsXH2rhAJ9seTUtqb9VWQ+I
Bcc+Y4qMiCB5y23W1e46zyMgftU9FHCx9ZkUzsb3nh5rorXhdQMMT6r2+GulzDbwBNYSLWNSoe7W
UnqIQY1W0wnq8AsdMR8QdPf5CjuvlM712PpG6L8STLo4Tbi2XpOQSRFAN/EPQuAbA16/NUNbRxth
YoyGPXFM8iDSNFIEiEt+J7xcOAagyDEsb/35znaJ8Bx0LMsC5HifpLM7yBTgZ7xM06CQC9HRntNZ
d+dzCV8EobyApzaja/AFzmtHnMxbDXb3EOr2uk0r7KiDXJoMiwpZOVJ3R6L3q9k9RGY+cT/clD7Y
o71uDe22w+Qx6P5Ve04m1m+Zo/ArVR6Suv2XaXwl1SbKF+hwlGkYRwVZh/P5PLuVFAxbyue2GjEW
R3gNIfNH/W0bBUhUsJbPr/TR8QvdNsszjtxyRNyIlVPcXOiJQSuU8zPmCvVgtmN0cIWOJXakhhSn
xZ4ZI1DzqFp/ej9Fa8gMKhlRqJe9HYbkrFKxjZFimvP0mFn+EjVcwN/2hI4H2a4/DP21O+YfXig2
B9228yid+0m/Q2dSuP6SmM/foMpaElFdA5cDTCn8xVwACC1Z8gzX81Oim57MPJu4ZcUSyNAQz1X1
Qosuqvph8W4/WgQHmtZLYGnWCmO80NBRcA+Jv4NHoPvOyBefreACO84wh/7b6+rG3UT1rIBtxlw2
H9SGge+7g0FL3DXJR/6cFpZ02wqFA8FXMwWjUvHkS2TNq/pieReFaLLp4Lj28fFjDDr3okL8aVae
L050hFjnNHs24jVbYii5V9iT62/G/C6WeRlVNo/vYIYmRqubB/lcqT3mvBYadB4C6dGTGDJ+DaKa
/bPIMvyaZc9rs6jJwHmMq0ccb+W/BT4JBcsEUtGOVs/WMcsySLmzmTEXlK6nkAMUbCHhxd6HmCfL
no+fpK7HFqZOwW1jNdMeUH9OS0aF0DjkzPLeAIkzZzumP4EA48tjvH3oJrtShRnei2+nxYmSLcrW
ERVKkoAYmNGty7lr63m/Jvd6zU9T472blh1U79KfHY26dyVYdxFPc1yjstzd8wnz1qVoKOJZtmHr
fBLy7+kiE3a/GsjCcgkioHfM4djPXTBH5za/D3GXwYc63z//4lgnnNWWfx6vZacoOMHyQxYO/mIV
H4zT+hSTQaeGQIvB7MV0xeoaLEz3xSPL/QinrkokHOGc7vXTw7Ug4IAukmOg+uD/T5o0O7pJV4Iq
/wr/ENGRojSTQzJoy+HGCTk0U4n7hC4KXuz2biMEov4B6Qkp1T8g1qrJfdOXBXiTWNav7G94K88Z
SsRlfh7On+Fk5RDyQUdVGn3a64CEfxqGxXLZO0IAjVFoJq2gJNm3WnK8Fhmds/NoArnMJ0koXxv8
aazIEMmi9ONaeu8lsCmAiAwpMD7Ol0LkJUPAIGsG8ytPj2+fKk4vB2iLSMHDrzk395Q4S1yifCq2
1FkmOjRPoxoX36/y0MOvBm4SsfaS+vQ9iq0gRQpx/8HNLTWMUeqFvw03FJsO448fl4eNaFKejIsW
SeCE06joTR3Gc6t5MCgPA2Ylp+Elq0BGTI/JW8fO99l9DKBgnTYFLtYazw1isP4ycN/fykoXwE8B
tMYVWI5R1BwIl2iwwCpN7BV8JFkIfNqt5QjQfEo18ybw2velqFBIXdDGslAmJaGf9dzh51kTG8iF
oxp6XJwT0shu5JACgXJxswwTggQGbXpOHOYcLWvYMW4lIQCtBgDyywu9M3N7Z7dQGExh65pn33L8
e0mwBvBFcIDWEVh6MpmbKqpPjPpw6B0U9farKku0n4jiDdlhe3SpSww63dY99846PkRl0GX4FQGl
gpB/j3JzL18o7lXrS+LioIay2owc7V6/zbgdaIYYwANC+Jt1VtBRbETofeF0v26G0RSE4FXaBPjQ
abRki7dDNL+Mbthf5L9US3BNdK+aJT42Hs+bkKMyBPSJCrJL1QRVcqTs7BSJTNVbOsxkRZmpFboz
WfCrBJPNhhT4YZXRJ4OzkA9+5J9gR0OQvvRuAWtSe2ZsQo2JTqyieTINnd17yHsTGeqSjLv2LHKH
ONnCiiJcA86iWS8XmsxSA/Zyou0WKgODjaanL99wB/gSW1HV+MVc2X5pZc+22L1pMJ3mQ0o+Lirg
ysIe50lGO2J1zVUdXo0B8ij/cOE4DHoYPZbAxWsp7O6y42mPSS/ylF5180YnaA5OjI9Hdmoj9HR2
l4MD1tp5GcMr/ntQsjA3nqSr8ck5b5i59oWa8zjvNDn5PnvOT/D5WyWqisvhwXV4I7V1I4Zn6eNn
6dpAL9OJlEG+nqUYDQ3W7XjvnHxDZQHxpv2tnEpRRsIU5VMd7uusBRim7V7n1cbPpwpBYhsXVltC
xJggAkJkakfiJ8ZT+WpPLa2tPHZyEQnmNhSBySseV0CAquxP33E7e+3vybr6tUQLJlJh1NDB7ZTQ
qasZOLsxk4Y3aDW3GSWGmumSQITypzXvSU886B2HqFxQENI5DXPObUYJLx8TaTVd5lfQz2KN8m9n
tRXXewkIMHjCCRezxVBg2IKKhyZtbzcYGQxFonA4mBurWGb6csfRTIRiiWL8UIJZPGL3dTdjzUyH
cXE/tu/iu/r7gdW3X6MOhqITPxPSZCOTfUDpYoVdUMs5/8crgAk7/7oekGJ0hHIKFmoLqX6c+yAA
z0W8QMNFPyP8z8Gu6vhETCHRr6doKANNoqvqxNWFskXdfkYT5Rs2jziY2RxUnI83WM1jQMx3Jw9l
iiiu2vQKZeC/5p2ji7n4CRn7nUHujgTqzoCtykos8vaAQ7sho2HIT1UxcHWfCT1tqBBE4CaKuIEP
+11Mu8pIURapn3MDVUCJJ+6p8wymsZYdouFWYfRLq4mokeIu20Wn46Ur2LSzettWX4zCnnVT+tHV
QYV2hyr8mitO6UKdOhc62gEsZaEipT7NeHp2QF7m9uL4KPhnfncdwsIZ5oEo779Txy7R0XE/jZQI
N5wN2spHwR00L0+Rr7Ip/nLRYExrYF9KRf4NVJeth8T5b63Z2sGjfO1XPFtqXJJ0o8CpOIOJdXyi
lbUib8uFJt6YACrWUy76uJprL2LaxUXW1SgQ6UbmMnkT1SHVJL0mSRB3dtXzz47NPoy7C6fkA0Uj
B+FXulAgQ1hxiGmA4KATUAP/mDcwoShsYhFe8YTKNDmKCpITrdZWaRE5qJw9P1vnqbeaU8UNhzl/
nQjq23gv5qk0gXgSXgL4DByQ5lxgroZ6GL4AS0mdIdY0D5+2Dml8GEvBKyLD8Nsar8B3SAqF4CBT
h3i3i/G8F56jTPNroLo2rMcAHgmRKvJ6v9hqPIzSAXXqgRxS7zGR01iBeIMGObe43YW2QvLZSAzS
ADiBwT+oDu6NEb0etwcT3BZneptsQRUHobEkD26xiiSdvIC8hMjaTbAwpMAYxAuC5tBc3guSg9So
hFdqAJKLD6VdxlDrwwmLs084MuUCdmZPEnB3xToY0sZi+aJjHz8sfZfLHiB7HMnOUoSYj1/P8JNH
q/KgBMSZHJV35ilS/6dKBl6sHqbExFcwhXtNL8R1rcpYk9gXeahfqjckC1PSjkuUIby49fHb8nan
Zb20qrU+rZWPAAjoiMPz9WU1k/N+TkRivzzfnuDD4JekSI3sCuD9h/DVy3Ee+uKxaBITZ+lpXHXr
RkC8sXg+C+VIQhevvW3ifJO/pTvdFgI4/PQAetFG3aGm7C/5jJ9sOvM+fIEWC0sKZI2SX4TYvxLx
pOfH013eK7uWxsrpZ5ylWpGSF+Wj6IyEW7ZjV+bR23aepuOdszs/PdUDjeuta+S54kA0d2tjuBoy
70KtnPvyLIJs9smEWpmUwHzzgfqKMQso2TOaxLACDNrSsX5skljZAx9gMqnneBUKBoD0jm473AHV
AgJdKMT2dx3CaKn9QnpcJsP5QJROaUS8cRwIUaA2Wdl93nzg4IEOLpQybXIpt8N0Am65ASo9dXYM
ZJrHyjQGF5Zobg0QnZCx7FFM+whjgAJ+roaOr30rmokEuuq9WrsxW/+pWTwl/r9hOh5PIfzOMbzg
hci8+elXMKFeOdBcQDc7ywSUzXfKRZO0W4E4/Bllox3kvbe81lNGgUtTZrLmnU/6Fh79gfYjT7ed
8ugrQpehm5j6FNjBSLQsUg1Uz0tTc1xfVnsKI1O6psbxd69g9yA2GAob/OxNdK3BS8dyA2x1HoQn
COAD7w/+BpTjCSRdwL3zB4iMhTvsCvYUe0igQHYOplxm2VFg0pciNKBNx++VZdLnvPaF6/wq4nSW
9Dyykc9F09U6JrLDAcmCAjP9USNGI1tGwi1KM8A+vQzvvoDpvAO2sSc61hi6PnG+JlBQm3QDq9G3
fzA31sZQcU7KK8h/LspEysH0ixsCn01Sux/VT4aAU6nSggo+ffPLw2RrBWC5346s1SzzLnSWnVkz
wGkR18vmr0mOQqWYOMeDhtDKxbaogLa4cfdbHHFFZ8hjjHO5LmOk9RSRQSZ7bJpxSAovquVZBvgX
og0YoTeVeBzHiIqMXeCzWxcpoNDdyGfid8JHq8DowgZOA7HlPKrHm5XrKNxLiEe8Sp/yd6iHMz8u
td/LZ8IfAwRHhAfUBmlwbT92GyzehuDm8L/A6mqYncMpd2d8gA/MBzpB1BWbJW8Jy4cs7yKQJa2B
6Y/EJg2Z4N0yuVKK8XFZGtstlbASxLu9GAgVEbRUE4TSFRtVJXO+AQY0qTtfQKn51cUAeA8HvLgn
DF9UAMjBRUbgAR2hCWkn27n7vCWVSJ2dBFFLPzBExkgzVKFt9i2U6fMnMXonidrA0HAptABZQd8X
EybuBdmKZ7w9z8pGSuk7RMKYqpUFm7Te7il+MQD7ocZZT28cJ6psIqdYgj2yoVLK20u/OxItLXLZ
6L3Tl6lsBzDWj/WWAan6fgGx/jFm75gYY7fAIt9w1wR8HJvIEZ+zlEzBjMshHz/JJNRnnDgz067N
f7vWX2ubl6ZAYB+5bbfavpw/k1J2yacx5fHTIVRL3WQ7/IQGskcVKfwBAIhfSAotAwo904DQl68z
1blWThiP4Ex36XVGxsPu7oyX7xEOpQ3SC2iaXuqqkq8porzK5WUJqMVnEDJL11RDtjmXXkbDVPey
np1V0DYlORvONVzIH/481tA4hgQw0NffzUmb1W8sIpy2M5EbIJMIcq5dK3pzTnI7J+3kOKOv5Wd0
lIixOqbj12X+hldRBRzntgUCH+suUVboFQNk5mHs5TqkY66sG9WgXhaBeZINlz2GyQEJEc4Rnt9e
TUchJ3yngjR1Q0WLE76gs8OSDs4lfnS/uqHMvnKLfDWqCn1laQbXl8LmSN5yiPIyFDIkgoJdhiDL
FF27y28MlNO0acMAw1BSRNbaG5NcvyE2Hqsq+JTJZ/Xcx6Brn36UeV4y/yECF4svVVfy2IYCLeYa
u/dJ53orj4nuHquFPuTshJHu7Ir3y8wQHwG7E7xXDfHaMDPp7MDOFuEBjdti4vcUxBHZis/EXeXv
6bLGsawi4tQ3g0PL6hYSL0fvcv+yFum1tELnuTq941W3PRbM/eTgqQSUvVmiimpZXqUZcR9a2eju
EwNw4xRXMC3aMgMr0gUq7yktfHLAzI0PXpDz5fcISqQ7j1lYp7RMK0ONIf9TgvIvpqS561PRoidB
z5K5sPdSnhPef0aHjv7jab9TUeoZyifAcGmvh5rmQAmwNY8hUHlUtx17h/BQ3SeWSYI3KXsyD1YE
zP7+NsbSpVZ+A2KwefSiaVENNaXap0i+rmFeZA2HUXsxrKdZ1O3ix+hS1UWN+f75tPRY8u0BlNWW
ruM0K8bf9FTYxX7Zs+NVt8E9ahC0eiSO5O01gioxsiKzaQUrBAgcdBBDSL7XqL42NSox8IcllhDg
4MQtdDoR8Rv7bthOF3dZLqCvKBO8U4jWAWnHS/IfwOOnFFtzA9O3BARG1HGZiwVYFppHOZ5nNTkI
IShkMLJTPtIED8K+U+kWyFmRHwc4ipGvXAToOPRppF0ZiEbNYTFz4DvfOQi7KF4YtxJrBVpiBV7l
8IBU63VdTmsbv/vY6mjW9B7kSEyemTmbFm+egZdtM6aIQjzpUV4YhRvVtCfh0yI9ITItZi8nBbH6
vMeD/YpiOwcO5LReDztboeFw/VMF7CRjMPnT9Ttibj576prsHTH/09PAPXp0nxmOYSts33jVJxNo
cBc8nslldM25BLtySA8xCV46G/rYLsnGP4Cj+hNa1r6TeLwpGbdqnOSCpCseC3p+1sjlrPFsBjGe
COTCSmzGs0EUDvjtjWkShAe/c+g6VGfmxGqJC3qJ3RAfhHWKEU6+698rvhq1yUyzWnV1gCAwoWFb
SABP3mDug9hcaDC7ELOdaLSN/88nnSrW/cYfDOqw6f9/T5Lw+/3UIG7A7wAVTZgyjL1L3oz5RJei
y9yaBaVWxuMNngbdYpImSHeV4Ndo2ZUn+LbYO0sLnnBvimfF1+BbriX+kX/ohkhyZMo5eFlbXBlr
nC23ghtCTUhK94V6Qa9JWeNW/9NiHHFwzFNer44sZirzFtgdI2Xavc6JIvcca//Wyrp8wKwoEzPx
q1YRYS56Z8QuIyT472vn87tAUWtJmROS7zSLDmJfiNuhUoJO2OhExjORJQtTNtDYcNklWn/DdyBH
bZzBMNq4x/z8mT/q7KIfRNAWHJUSwiLSD2NSrtH5Ay/n+gfnh4sy0JQ4luXvqf8H/fDO7rALltBp
PlJXVrJEvj4PjhJ2t5m5KrBGuiIkaeiDu72Ulrdjp8DsPSG7FA2CRHoI3jD1Gn5TlWW+cQfxav2h
n5YmlVCDb/YBPLugjgdz1HH6Jm0zrrZTkk2WWz6pTp31NkAJYZcFXd8nLkg9MlYd3wX5+FMG5pwh
vAqAAcL/6n3H99V5BWgRb9aZqN55uEepQ2eySFEZ54myv6Tl4Z2IUSE0P6Ofr5Ktj5W8d/KtsaiQ
QELWuUdIYQMMWRiiqZF2to5Y7P1xYCU5Ot4kvyZnKwyll8oo3YFVT3/XyPyVZWFj+l440BRcpWbc
uX+A9F+ozdWpyaVTnTcyGoT88H7IBUm6agMdnpiLLamQ1f0YbyEiJv1PHbg/RDshhZzehVms7LvZ
xkejFaNgpoVTpdIDMVVcB8ZICPNQCUy2zFwGYVaFOMPgMMNo9XtxYayqzumrPC9Nz8rnFcJcYK7Z
+qH1v/vyGGFV01icXHAaJUVUAn7oGJxj45SqTaoWyeyhYQ0AmnEMvOaBIyGvmxEkBKMSa6CzvjDO
4Fqw3lTKoW9KKE6mepKov/e6erL4gj76h3Tmioilkzvpv6tkzD0CQihtadYd5Dhqy6nRyESPPaRC
xnZOnvKclaXkjAkEpxb6vS9Y5PXjGO2rAK5BVIgGmWkenENMQ3u1MoQffPI3qRCCnA8GuNHmYVrV
YSgHtuA0sp3I7omGKoVHKZjuMavZPLfu02apN5BJujj08eW5rmjgs0xyr/lzp3qm/imKz5m5ckfg
6a6Xq7vDloQ4wAhxI1zsDHf86UDHlnNfaircpEPZYhpAIRlSkaOSvpvKLxSyHWyqGGv89d0J/giv
AstDBpqpUuVVYADQRl/OsvNLeo60SZqUgW1jFEihdlxJPSf34NYvN2WSnSbY8aAqu6ZO1P+IzEqW
H7i3cD/+LVM7kgpJJMZDgBPQz+gGPghHgWZmS4kKgjI/dKbWB/Tin7p+Djs87Z9k3kg1gVuHCfsF
kd3hc0+kGcB9eIJlhTsR19rx4POd0VTLEOhn9HTv89ct7oYQe77mfs+lGra6lh1+L0njYfPK6wce
WvjTjUtZmRsfMYb4HKfegiUqRuHx0xQSKtC2vsuPYQnN77AI85NcNoJir8aXD7+aMxaakUHC8sQh
0PNw2iwvBw/04gX+cYHORKtdO6jX0WqBVIal7UKNUojAe87OJSr7TPVEmWDbzrq5AGIU0CdLSJpN
OhgUfeP7EF0MWzt+389e/oQXTa7MITgNkSBINnMl2wiQqgzgNBpHmq8QYKKJuS2uK60AaizD+Kxe
48ZkMWfRv+Y3xV8hVDuVDJ6RLVBPhf6Q2Acl7HnBgSKztuhMLPk6IAAOY1nX5r/zPKA2tu6hsbd+
G5PiPIrmmdXHULEm4I9uOsuW2VTg2vlLGjx4SwMRWYj40UdZoKqc0RK63PWK7jNBywvLBQ2+oytj
unq1PpHz/bo/C9brkP6oZ1tpp4kA9xO5esqMxa2ycEPHLYVkLwmr6Z0utdgPiiolEz6OaWyRYa8B
/VyNtWy1m7t0uNRnfyYPnYLjcrhugmixJLYpr4MroW59lZIJXMC2N0IM/LrmvjmQmYQ+2Jftqaxl
M+D4jfcRQK6Vr59o6fOFRWG5tPNkofofm6tcTdoxabtJ/Pblo+mRhAj4JfBU7QgU8sfqtgP6VM/X
c+8B7kYWPSOOQOmV01aeNpfoQ1+hYf2Io1PBpvqp2d7OnwrZZYpyMDILh95in9ETKUH865cdrlbj
gQsPku5IeVeVAkcDpDC/fw5otnz3/cAtIjDTs89+bUvdbrhuf1XQaHxI2WGqtA8hCPw6avU3h8tt
TuezrIT1ngikCngquBhSA6YQ+b6GePsCyXWAugt2+i8LNSVs33HYm3fn0hYn590NfTnwqPl7JwPn
M34vgQwoF2UQvvktDScMdg+J0Dzt0t/dOQDLzCddpIIxR0bFzOb+W0A9+dFw1U76s+aOzNqVc0Ki
s6+1pJRA116xp64Z98Ol4AL0vTyD0kiOGXZ3iMxL96Dvw3rsl+1zEJOvXFyc5QG+hWePJ7e2hGBH
kJg6iQszI8dXFG4bjeq38v4T0ZFFkEewSQwOjHvlisd+jl1ugIf8eXsiFP+ic0V1NTxnmy081gid
g8ynpTJQXfz5sPppEfiQrfhZeeGT3b8zcIWH1CNnh3tck7WzsG7kM0LPm4E1Z8IR92luWcpYPewo
GKIs6nmC3bLsIsaqyQreQtlb2dwHUhbOzv66+/61aw2/HNDu6MidGu5RFXPeTOW43hxzl33fW9oh
phadzEJ+vrklCADOkIq6LndRFdpfLPe6VVnEHQ1pRYzcxJQiBxwXDHgnqpr6dmYTIQ1kQlDlNzps
2c0DfV9DBDjz5536fqUyddMG0IyaesEovGod8JzNBnPpB9SLtzRoE4M1smSP62eId0WhnnbeXpZp
JiFxqi4nOsE103sBcP+4e/WT8pip7RjlHTtuzKbkaQN9wCeJS6LsOVG0GXrInemcVspJNrjrPc3C
hdpsgwYXcIT2r97NCrhQx6i3ryoaG9Jq971ipLRR8/CxXZ2MOuxWxoLxw/Fv9t8mOBozq0RJLoYG
vQuLWkf+u5tVUt9eM75VwnwIslgVqrwuZAcnzYKentnNMStWEbAZObDOe/auJ/2omoK+c84QK7CA
K3kYuRSnHs9szRp+CtgqxpQDQcfG/InB5lfulAuarrC6M4B4b7l680PsUcm5r1k6sYIS0p4JjEA1
0KTddpma/xPPKiltAaorIJ+LNFMF89NpQVLDVUvL6YX6Viz+TJNNBc3pVA5sxpbKfkvcPrFmQvP7
abX6sjvvUfWxNoe2tMRBs7nc9948FnIi3Bh+Ov6zKGXCKC2ANtbDWQt1BGZf9PF3Ns0jbhmkKR0u
d1/IwBgcpEJH8Ah6Y1ZXFJ4MIF3IJUG8eoQRNPjpW+DJvmNHxIGkCqp1XwVMncAOfRcxe/R0LXCb
wHXKaTLfkMGH5wpXG8r3bv7ws9vaQWVwO8764AFfx67wcnSkvkRXvhkvh6Lkz2yRZYj1Nn64PGkN
vvo9yH5xrZ+NVA3HT1fKbda0tkmXvFBU3qskqrc/raEDDTb7JGPj1eOHKCe5IEuV2tsDS9Esa25E
5IGD5g9r32ypD03k1Dtb+99Ai+WU00teCcVVuft7KW9psW/Emh5LdKa8skG9eQd2a76vyiDJ8cre
2n/dC0w5Nwq6jjUzWQsSMA3XeyO9v7wWQOcpH3SWFIITro4OmJpFIDqIziM7ptqWuW7OfcjUdpqL
rnA1o9zzqr3DcBPVHiyqmrD69BPBStgGXcQkujAvAZFv/x/enC6WaUcLgfKTamyv2ocCdOSEZB/e
KCjsuiUVls716SDOdfGXtxm/rngSxC8p6KTUwipK0uKY3Jb9Z1oUvkxXpGCuT++iW1D1g08Oinex
btsqIZgCQXxc3jltf2EL/Zt5kyXW2KpgRwzF3U/J9EfL8D3og5UHdWlam4Pqukti5Kae1PJXIi2f
V+EJTXMocH3jrtXXscIJ4G0M2+XpFZT7nkBEqOKEfiffe/4E0D378vbq/pb6AXtoGdANV6viQw8t
G9rdyeY4SHt/hu7fIP+PHsskswG2JRwcwP598Vg6OW3KDoJ5HB6KTwk7CIj39103iYq+rYX6W664
KruopKOdNxsQrgErvObEaik9VrexIJi34g018dG1Jf+As0ax70g+EpIBrdpFsghuqRyzYDtIwuH/
qtgD37KBYZZHKlcyWQRt8/d3MvV0WywAVoahaMHxyQPFn36HV+TFGgtsaIlqoA/3L+UP80W5/jNp
g2mlYcaUZ6tsx+ZUCanL6G9SQSXm7y6AHDYszEOknLs/lxS4eNjDsKtlTfCiiCgPw3/0Z4Z5jq7e
TvpYMPuJ0wET3Tk1IsHQhLvSW2eFsQG3EhKjYvOMuV9taK5pdpW+sfktxr0ySLoHiqjcI7Dozdh4
YIr+q5Tq9GY66Gv9lsbkTb5IiMDQle8CbX5tbmAZqrV9zExGLPUPI5aVL/iOV4bemYet9RKjUsEn
uq4ZdC9FBsBCq1PnaYK1fzaF3+RiKau4tLIH7znfNv7i8sCJZ8RIp4fqpu/dXTGUfO8LYtqtx+R5
e5G9cGWkqJGAdH5J/SR8uoommActV34LA26QhUWC39pXpLFcqmvR1I2bCyCJOqKA95BmYk6eR29r
INgXTe4ccqNvEluzbYCyoZgJy6MpgfHp2XUplkvSo7idYjMG9AqHapsvIg/LfuDWIz4qMJJEX7ok
Hfg+OGswUdPdoNgHMR9QZOUmZEkSXuBOEIW7XLg1eeXuHJO9HkA6dJ01SMQB4rJaW5802Qo2j+3N
UqKv9quFNfOhSytjG4ZRyuiFJJQ4PZ3VGk593k9NZR4BF7XwXjMkkme1bwE3P3DtTL0nSzeUB9YL
ny9DN0H81DZIAs4C4fqn3zehPBWdLCR70SwTWM3zogbd/1B10HHcXD+KMYh3VxOq16EAPkOFEME6
73J2ME03yTWtAPu/Q7JB/3ESB9Dolonwx+MgcQsrHKCnqZXOZysBjvQuY1Q3vdCW4YTKMdIXUIY2
LKVEViJo2AVfymwDPkAINe5cyT8TZ/GyIKSNAZUKOJmqqP5vbAzeGyEy5v1CUobXY5m0dBrLi0jN
e4TytOZCJVO3B43w2sbAUOY+f1IpAsn6d8q2TKZE7jBZ4cHTCBys2JMOc0LqZi2HSXFM1hdgKSeh
1WbvG+wtCLTdxVbrGw+rfRZ1NyPMCKKJE082X8icppyQjGiq8UisxgIbvoWbcYNYhI1wiYoGkkcC
bRmHny8r+/zMo8WMohGcdeMgdq36ninIHx685FUaoV86madt9NQdhr9IsuzUT5klSRYCtCSN7bdv
wdmjsum5yVBeQvLV3lv3ER+pO+985m6Hz3mUi7VecercoguRwKIaDZNwzwI1RoS4LsVdIKBkpevR
u5Xe02UiZb+o1NfK8OPfI98WEQjBsgD7XzQHj04cI0RNohzx1tci59IUroyUd0bOFoSZHd6iSY1s
7MlKqygK/i+AHCXRQ2IJEIQBC6ysRfMKBSD4EbIimv5Iy+KrD7RJsf3Z1RICI12UssagvbDdFMY5
EmGZ6fDslpGmSFu7Ti/zT55PKRoRvgLa6pVsgQi3AAXuJENuO/K/PrS+iR4E28EeI+YSsm8oYeaW
h3Sx2cb7NA89yHj4utyU6PveiBdh5NI88tJYGf3jP64Z0NGDho4LDcAaYoKgsYFOYBhXlaAKDCvp
g0WXQtaHPZXq4ganTAeUf04Dt0+ev+M2YKiA431xkSKbKjvfDSBJQ7JQhrCRAZlmNxTvI8Oxy477
CynSNYxAogE9dcq3WXx2K+HMvSaXyXl/T6wiHsmZOHvWTdBxeZT/tjBEJSlKIgHi/mSfd4Dmsu1b
bMldRZ4Cawjd2o0kfj2Yv0g+rblPyaUDmFWZv83oOiyP7cYzql2PFnFeFX5ke23AUWGcxHSc7rR/
5lJAdPwZJDrRx6Ys+s/oEETzITFKyPiKY5vnNfm0otVMLz+9FYqtWuQqsiy088LhZFe6bptX4Pt0
lbQOlE7gfnl2QFBmgUcg/HKc3D1C03Ieou+A3kwzrOKahGQRou4JnovQeZOaMUgPeTFpkhRgDIPn
0BVpfsKV3Ryl+HRpewkFL8yaxz0PccEw1vev3GggN7bfGSeV/lSjxqTf7QlQ6PnuXrXFxwQCT8ms
q9G3XW/kWsal4rkWl9TFY2PBRajBkKIZ/v7By6DcKAxepg2Yfnt9Ij7LwibiwYAEqFrNH+M0FWgs
OSkNLgbnTfJGPivkrWx9Tzs9f8ux0rrPA/5+WkDn7gWr24ac/Lk1E0nrqFTk09GgtS+JApQ+x+xb
r1LaeLkSuuKk4WbYuYQsKwias77YJ+onL9IY/VPiHmIPYyVF9L2TIMFKW9zQ+mli2edKM3omQsTz
FoFATXVDESNlHzTJQiyuYnI74hQqSCd9CVCuy45NXhe4IRDCs2unPlBXkC/ggCSrYr9bIoYZPbP7
unbGOgdnLVlmc/QuNfxgX8K4sbxT06RBKKvMtl261i1fV3IwMlWa1dcQFE51SO2xAxTNDpDRSrDC
IGoWXjlJjCStxC6QnpjMcx32klR3NAbE9EoZpQ6V3UkVCZUMJCOUEN2xsXcfYyNep/EkvxVjXabD
5LgcU1IiYaRMvFhRTBW9o8FSnvrEDbrFUuKuraHhfL/DDOK2sLoP/Dd3j3z05kM2npYdpxF07KTA
HfE3Zrfrx8rX6UVPblkxub7K9q5A2vKjTP1dwZo2f768I6a2XiKRmtN67gKfO4JvY9GJBA+sEZTK
wssQVtIzSuoi7RPCvFHBJIlF1iBo65MxHwu7YCxjX44oy48L+p1BhVHCWE9FhnPSvXtDTwTHJl9/
IYI/hj1hPRYuphzeo/cCjuJWiSMWS8DXaJnFvLm8FQgf70ipBa05hIYfg9hB7Gfy8koo8Dvk13xz
7fm4QdNQ+NDTHPhDn6/5mc4GrQUJe+/baN2nbPLjuhI6who+MUd2olup3XqajVr8DH6IvKHPVRtQ
QaTlaOE8nXrkdDrtyTaB/dJ7BXJtkHAfmqUNa4ET4CtYUhHYDTAMBHgSmJS9GOLa0cccuiyZS2BM
pfIoi/skIrdc8ofEc9KHfHEHH2zvYQBO+RX+3ANOrPpt+lAvHyai8xQ5oFgFDuQkBTHmTWH/6NMg
eI1MOj6/TO3+32du6u4+tZ+1GbvuAdSuN/cJd74xOLMqqzgL5o6/Zzb7Jx7gYrFS99aBqonmJZTT
Iz8itfp9gV2HKH1JIP7f6UIixHVTMJxPL4TMor288crmcD0G+4b5/IuCVHK4jxGjLhlLD4m/Dizv
qtD2eqoDfsQzIe+FOvH1VRuUuSLbA8Pqcj5iKYHW+Fm6R3+ZfKCVrGH+lDJTAeTsiRp0iKejq/cv
0uHTvclQSQWBN6CtdopMVjNl0AR1pPLQvApJre7LHzCOBQ+W+JydKI4bYOAP5dm3N4ly/7ahiGBR
T+aj8vwRUNiQiNBnSMBh82eqS/7K0F8Ah78o4wHykzei3WDzhKLyBF7cnJ+jRatSQWlR+Jaqqg5a
D+RCSLNjkMdjprLyuZl6Kll/ePCIXnAL4Ml7uh64MK/Liawa9LulMw6NKeOpQ2/Mqu+2iSZ9z3aM
gN3k5YKH10jqI36GmMJYrmMHW7rH8j6ENmHUvtm8Gp8YWbU5NwNHKfiREE5Kha69egaFUo/bMOR/
GIdS4crCiayUrD/Yf2OY9C2zSn1Yi0Dx3vGKJm3ixANL0ODrSim8DQe7eghomtZWzU0Ut1Lbc01q
gbM1KUWdyK3pykiOLTC3CTsGjMuJBqzAeGtnNL+Kcy6KgNCHrvQ7nedHT6SAcuSlApU1OgiTzeLb
z6KHiSKyF2jyEDym/whvNg7h2kgYGhBf3uA0N0rsjaS2hqT0HrNBt+V3DB5c6h+azN53gegemwHF
Pu2Wcw2KeosIq+aPwgF/Ds/4XAnc5bUFTMqC0xusXaIkwKtUDGwSXFa84PtWZjEbxZUlYGuz6u/w
H5we5dGz4VtuuHdse8whZtAHpJ1F6NrAYN3tHUXYMUOM9BKfPlYJl9irmnZrRhkEh7VTVI/bzFo6
ttZOjSECaVO+x/A1654LF5JZpzxs/QWpj5OUZQbYDWilk5Eug/kx0JB+yNJdxtBJjhKlL8EiHnlC
ltvPLd7qIpX6PqDKq8YPO17I3VcQP18YhksGiLKg7/uCtFSY+GRRGG8s6dSfT02vCmvf4OIk/Nj5
PK3vOoftKjKZoc7l/5MGnk/XZ+S4Juz1Ik0fau49YO7U8csDpryrylrfYZ/wjo6HCbSNGUNIjQWl
pO55h0N8ePaFZDOKpDun5mtWFnWT/uaT2ew3KuADRa9Hq2zBIQTAz3Z4fjm06x+OqEuu0gKQZ+9s
SGYG1cU7+dEV8dLr45brrnFCQiK0PxE823aCWdcrKXlGYVWuEPr+GGqpACnodChHbWOI88h0xjvo
MWXOqpyeCFIMDxbwmhRax6zyBs8/689PIOB3WliZ2UzR8+63gi77dTXZm5dDpCS6yDn3djjHCxPd
z3JypcQNB47IAvtVyR6H+TsXXAbCyfvT8il2RKKnrXz1h+AMqSCibAH6klYrllxJyFdhKu39bERc
Y9k15Cvfr6GTlg5IdeVyLqx1unVlSdhiaqNj+8m525R8NTuKi4iv7m1KbNISRj7OQ7MH5Sf+Ksg/
pCo6PY5xbNWCIFWxiVOUDIXh6bCPDwxgrQLtfFRKt6/MRNmnw2gOIluT+vJ1QCJhylPfQcLX7jc+
tYdSGrXzDxuTWYhNpbcNYRI5jckrE8YRUUtuNBL+bT6zFkEIbu7XbH4FOVbgfCq6rBCuZ/PqKDmW
95oB+IVrLUIaPOIfyDuyeiBh846QNDvmAEEILK5mgeKpRHzom3asUDt05ocJkk5Kw8OK5PnWQOGV
FHXJCC53fJeV0LABuwk0sy3WdmNioUZUQDGagqse6XwdVjEaPtZsaHRHAVcNE8k/qug0l4L6jS5F
of+Rh+DukogWyqlVvCIfPULPM1zmfm4T340hlocB+HHQWcSpxyCZsngyWylEYlhSUShwy5ojaetV
zmc4Kr5PaB7HDcOrOHcR4p3npgJ+Sul7KtBKk/qUVluIUTvJlfcCb7ph6quV+KiXJLrKEG9nc+fq
85Chqly43bi77FfCqu5kIoUYEVbEo6OWbZ4nZtNtM3SNcjqe3j9aEl97hzkZ9dMvsx6tCf/5OIBh
pxc5yTD5nOzQoAnWge4nDCjM1l+mtFM9GeG6AGd2mrLxxIFZLQBQquMZWrO8pWtp8AtHGUHjAy/g
c49HzotVXmCHHjKY66Gr/OIswUNWg1ynX+viGH2IKD5sS+09QvA+hzeBZZIiENJHan0dVEn9if3j
Eih3+14JA8X36XuE7kxLLuKOfAJhnQaQq39d7szk91u4uVYT+AAAZuu1Q52OZQCHaQCRx+eR5OxI
UrN8niLHuCUnLwtRxIh9qaj3iewrFBbBGO6KLIqUJgmjrfQOHU/NiZdB5M8Pjia3kGgTDbCYh24s
dK9NZY+4+isIhGeUVydAOChc0gYrCCzgERH/FSHHoMCJBYIYKH0aTUSJ/qn7Xts5ffBiibpoYRsG
LhN+Ol1JZ1hfK8XR+pjWcmlAzbTxS0jMg5JhkEpI7+9e4Edrxos/Zdgr7JjIyoqbVVG4lUG282Hf
uFIAtcCZAIekFxYw7rj3IszEOygewuF5ACHB9SLwf51umtWOxDyEJW/BBmgqZUJiHx5oVc5ZWWON
r/nVfeUOyu+T+dLlghmb8YNmnZ0e4lPEPfCjtftRzhFjY5ZVrOrXBk/jFn7V/rWH7w0nM5aX8MaR
bnT7tUbo9Ek55VZxpTY7BHVkPnfRpVNxhyjwBrehO9urcHjoVdQ6uHK/tL141DRTAk8v7CoDkEeY
0dyIRtYJgm3I/JWZtBYI/8e8hPlbc1E+7RblfiDEIf3+60O4bDtM27S657mdJzwgSj5oMPpnIx7F
ZQlBGWJMxM3RHlLVXm66l85N1uaxx5wfxIQ2/0SofS7ur7vxsAq3BCkGfvmLlcDhGHo16UmFQ6KH
dguomKt2bPfOrsZKK/qIzsVUu/P3kUS7mdUagWl/xdjiU57YaGmc6qqZ6bCBlnathhEHehPMrp01
prhELbhdaysZU2230v6KxzpH/yMMiFK+OfztuaPYBezGEzGSFD1AX/iYi5MaKhuzu++zVeawkAnA
2lZgHhuaaZGBljDgwcyJY2PqORrUXixvx/gWTpy7P/YKbUM5u7ByFyWLgZK0brz4WcGlkVhlMQZo
F7Wzr2BLKWSIe8NbHZZ7Nam+sT0R19RIYqMaDjIr8OuX8+BNdPXPbrUyoBZ8PSkr90I3lg9PPSfq
O6ALPsY/6TxFnTcghfVvKxlSuaq5bPKEQkHIzarcQGe6NVeon96Rnj38j7cEdkKFNhVNu6iCSFAJ
jG8D9ojf42CzH2BPi2JPE48urQMQkubv8ynBcGZRqZesUjimZls1sXl3aPl7QapbSNN6pyKPOtaU
13MFRILF6o3HVIXotQ3KlBq0Bw5YfR4jy0dThe8HsU9aQBAAlRS1V17y1whwzlR9NroG7DulN9nT
MCnXLnYEJGFotHHwVzwU8By4VWq6a/fwsP1R8swj1vN3glvsxd/KljAtnBQNkf6nt03yXrcdf72j
9iffdsejCF8LvxY4c4fHXw0hrV6EdltIPJKONMA7/Hhn2zfEKYFhkStKd7D6ChQEjI02R33stqpx
onEkIShLAMoV48NrFAvVKaPcWtKcfPts+0KhzsCnAghwUBpNxDc/w9d7U19Qa+n6JXBp5rsZIWze
UbXXg0Q8K9hUKs0pfQ9HAC38LY9zhMs19nyaWLr++pHEdPBf5NCns8Dl3srdIB38upUio59cMvFF
361rFPNtZ5c0vOn4LPDzekDU1h5SAv/ssqmIzU6e58TRBEFZt4ZTvgYdG6JBZkH4pjjTpVrNSQIT
yGFCbaY/yYes4b9v+jOTfGNDSA061Hu+UT82H2IZiQ/URK885KcnBj3Z1cSwcHcNoo6kHrYwRzn6
h7Cpd2G2RSRpa5ucCIjPEtsJUGMYkxcxG4DndSUJIBZJ1nX4T53dcHXDHVoMmJZZCCtJnFOM+Epf
4uz7VEe0lxNMro3DieSfcyJE9/zWGQJZzwrcVsIccx8GRPiVkbSmQJ4ZvL5QEdxsJoK9Z4+8jzJY
lMBE6AaHNF299mAf1BM3bj2z9mog62TOExGprwUUfxrMTLyQLyB1Po6kWePd03A10t8ACtqLsqMj
GT8GLg/E4kQxH/8uAuYfXpThA8eAnMcjUXCY0sCbfHihY5BAwWne91cygYg+Fh6n14Me+i6WMK5E
zTPOpM/omFAP6TEb8/OTOzwBPWkzPGCTALHcK/ztD7s6C8uoMGjDGY8qiLuV+bWec2DPrKEU1oXb
Ho/WdMXOa0nbye81jaFcCPPNn1oQB6wppVjkX8uBZC20lXNHyNZK0LDahC5NWwcaDaeJ/XY7G+Cl
mrB45hVt/Xo1poGLIiku99Y6u9GrXcrGQiNBT3dTJxZo7/1AdhtRNx6TrcECA+xJuxBYRZEid2yy
zNfNJQIaCsnKVWBVjMwiqrGAaffTEUJQ8xbIrSmVZZMLPJUi5/I9A8FkGeTwyyhvAM9jWOkr0dMY
RqjzUYWv5ViawQqAQ9xMyXTNLd76BFp+5qPgQQEdC53kpbIJ+xMvUYuXximSY9udmU7PlCyle3iM
nJgxqCgUPGrU1BmW7Ee9vK5QVsduBzsdjBBhQVcb7w8OAz/zAYFvwFqjX2XyWQV73kbjOOkSaFZc
R4ENX/b2i7I828uoYL9A0KyTOb0t8tb2mDxBiHBzN5J2YiMRjXsPrwN28qy0DDj6y7ndHKw0L/Dx
ytRICY4V6QRabJrY1EX3GkNI41vvXHN1WE407BmEh1C/BgF6+ZIvzGsE0u0mOT9PCweTei/cVzG2
UyaPPg8mmiTtTa7R7VKQwF61NXBaTiGyHToCI64+Lx6tZzzO+QtenC42U6qT9TAbdNzhrynnba8q
f86NoVVkC7eeGgvG5zZ6NihuOGLarsrk8WQ72+73ZP3fLjzjRPNMlOsoVLhYvJ8a6IDeWTgjcMss
1PVB/SxzNaDdifIEbxyjnliAsK3WFdnWjyUjII+xsCSw/zfwQJgvShQ8NHK5ZftbYtLR/DbQ3gwq
gqL+JV6VdM288WZBUKWX5glaJu+pXaDyWwEGWvvzFWYuhkn1G3/AMlLPfGFP2KzvG6Jai62p5Cb6
hnVWf8uUpjL7+jx06xFWkpzXIA/XVK3AyE8AhyWq/hn9Wx5NLt26c9aJhaPFuTo9sHT7gDUWCWRE
XG/U6Xe3o48wenwb85LaBMlGU8nksUM6dHk7CRmkJGwa2OCRIxwbKmD93nhXqGltlK5WVuomGJXd
Y5IbLcX1WfzfBu+A3OMjhe0cQuJzyG+58hVirC801+aFU4wYTU/ouKv5fvw/59VzGilwTXU/C0b0
OOeyPhVYvsSF8tggRlOaVAnhQ4Io4qgnVacsWC52GApR/gvrNBTcUzixHck031MxIHsCRNM7qn6B
dFCesFqI+EUN64K3/ZCl2kie/nQ3c9F14QL3OOs2tXhGLLoWk/bpw+/LwqJgsbRdM+vE82ipsKit
t+EwwT8yLgXYctXaQekpf6B4ISMnJLGP148uR2tnGlFRNi/yprjgFtdGQYr1Q1p45ETFFcT98qmq
Ph1frge4MykQFg9byWG1A2BO+cnzx8bAl6qDS6WiCLJ9jdN4PmnPm4o7EBo7OgkfyWCN6hzqLlkc
mRfKFAD109YOj5w0KVX1nXaX/YawgLmAHNwhs4NCLZ/B0PZep/TZaJ9jKyZjZQIjbGrPiNr0Bm5A
FOehQxwa1wVhk08wFhsdzCm7LsoZqIkvmccf0kT8KphxnWAv95yammLGS+g/Lw1SlerWCLvfQNeO
p++9nCv0jNlbOP8eS/db2rIfuAPBM34QnHUhJ1xYJdWqKXDbIAFYtJ9xDTk/vKrKTjCLao0kM8rK
6FNyZePuvygL0uqZiw6wq8z3pR00yqZveqZrc5JZwboOXKSKSflcXB9FbhCBY5pKCAqqUNYVnDtB
xUhtNMoLWeoQQywHDecWfcVBMPLzSwodsHsWuXBaITLPH7QP/wsbJC9s6Wv6g7BniuJBvJYpHPyP
NHpe+psHp5BGlEjuw93O72qsdh+ipv9KgdO8Q4NjNyfMzosGcnHm7CrU9vh3irdt6yGR1x+wKkxV
GAjtL+M5aBGWZWSVhYp4+LzHMYVLvZkWVVJ5FC8Nb+NM+CC6Jcj37qSdpG7vkMgn6SX/XVnGbbjk
BTz7eHg8ovmSBnRSpVvNKY2h5V1F+djMuDrlBbSK/d/Zg0pbK4k0YXbXDAiMU6ON59Zz3VhM+We2
8jGBuC3maDCdBG0BLm3rC9J2ntzJuC0pMiDcB9K8Y4Wrx+OFf5Ensd5BxokZkwspEDTG28Sk5QxG
5Ry2DR1kBDjLB1aqFWfLEZvFs+agbhC9zdSgBW1govmqPp910Q6Eo7alOvvtj6m8E627628hNNit
9o/qXd8FDUfgCrYX644+9LuywP9pxLoRJ3cjK5pE0kBvyqIdrVceKg+FIe0wLhE+ZC+qw9hdZ1h9
P2Se/S6fB8xAIuBCpgVgCZXE6A/INQseX5SiaK8gwhefupu3agHUbV4Tp1sTSSbX8K3igdNLsh6V
3plfmc1Dzuc3henpZ1CflmGq9n5Xz3ZwCCfC/aRzL/3l/3V1lVJ+3HsFD1WBQiadWO7bVd7hRPpL
aEaZF93LdPcOVzTxbsbKjvcgYkxnvT4sh/HLbpD6xNJY7sBu/Yltinv8Mu0eqw82920TNrNyMF7s
N5XpA3B2DpwkZ3AjJxVdjW1iJwijMKEs5M8rrlPYOCHZ34OpA3kDHhNRSaeS5g6PIxLXfpgnlT/A
EZXf2d/DPXJC4LMyQcOVlG1VbVvNp2xkq0Qz/eumoy1ClzlD5UH0LJrnHXzoakZ06HYUK0kKcnhH
LbSNVKerKH0gAjxQxgBJcYJt4lspAo+/8NZXygcnCsikcTtOjBWcuGnfz6TBFieCu/O4dehxG2R8
b5CUQf6S3BNgl/gWM4f0iUOoeRHPFiF/xFYxbffJB9KUYtEfTv7CCQpNw+qoxLlcv7L66OT6b6F2
0trUj8oHVvbqZjrqR/YOD9CjTqcYWG7mmDB2A81KGoVMDVKoF8Qg5X601rJiQwPG1t3Uh7cjI7ak
KPs5IuuRs8GDYVRAWRfxGph2z2xrXbdo7pOMtgGjzX/aV2RqpDOVUar8RyY+PMT8lbC2xG95XWXT
HGC3G09PHgJGREo4yGBj24czBN9tK5/PLaTkhXCXHRhyLhe+IZXfR75cqmd+RDv2i+XFdAEslOFh
KxprhoJzdcFMjisUNtnACfYyY2HOsoJ9nekcaXMPta7/+oSbgtGQ4ISQEnuzXWAphhkiNgJYnAHT
/BNKRMnXR6VamrfiabV6c7ZaI77hk5t8Ld+43k2A0UltP4QSMaPR/g/iO+SPVfnatSzcwjWTQf2X
mG9haoMtF2nzp95d1ZsaLsIKE9ELs5yXCPLEkfkro3GAlmJtC5QN7tDneL50DqSlbX6U6rF6L+R8
dSZn9x1cQPhFigne7+5bqujG1rURadV5T2V5uuqjHjMo4dCDCYPvUzXWLCWLufed/4PjP28rKcdD
MvP6oXkIDIqTsSyVusOMMDaTJfYZbmwv2catUwlITXZscgYvWB485hzXKZjpmSGIk2tc0QsYWwZ/
zAPfThlR/ZFyqMjVbagAqcEoW1xx096d3r47Ml+UhrhY8KM1q9UteU+nPwD8Roz4x8ntdNPY8428
oC/893KUhpZdNO0USbCBmFKgFemWu8xWunDkZikw6zx+bg3t8CJLjuezUF1kxwboiRqrSEM0Gkrg
YOAqPVfdv6aa7vdNOByFowDgbKnUNiQs4FOu4dfI1jTS3GMeIUHrjiYLvScUOUNIYgKWTxdZU245
Q55ngnai3zVosEVfbPoFgFIuzQm0idwr1ivNRZ1r20PgEz4wY5EfUGhW/8kcUj893um/v8oAhHlf
aezISB87G0HhOYpV6xbiR/tzbP47xa+ysnV6UaPw03f67VTCuOzkiOd1lFhqJFKWqxN/ArbQbDHr
IVitCsjSwfzm7hFGTArCrW6gbBjtRXQERQavXj0zZwMBXPxkXBZg3GLkFNK2BMubR9YUSuk5QaKM
PTd6BI7iWj4S5jR82ddFWGCbbCeC93QG/e5qNfXCZ+ozZvwmnIy/4enNCSMoail1S8QKSzyc4EU3
QwmnI17Sbe9+qVcMrLOq60nbwIBunP/COjUCAavYobZryBwLkroxXIOZqz+P8i2IdxPLRprEGM/D
J0leLCrYn7s0ZJCkmc1ExyJYqt0hODyWpQuCXIzgRoBtXzW5STtt3JUzg4d0KtFCPPlGAVGHFEPP
7ScUK6cO8ZnzVs1+5iw/UMVW4db54B4kuRFE95x8yAB5PCjm5XDd6nbDOmUO9/k4jYn4eAKMhfxr
p6JTu2L7jHywyX3TPc/S54m0DAkWiEE5Cf/Rt9pOyJMeXPk7LCBtYqwvSnGGzsc2Afgj59z7JmV/
kLR+SLUJrcqr6I2B6BzisFch1ts0VNgRR7YsJvveDleb50yxG2PVuQlmmAV8NHOK6V2lpCSRC4dv
y37B+OOGIT7cx6xBFkTajz24r/OflLtM09tUvnrZCATtnUeAZIK8NN294/P56wKrbi93zGDDmSYb
M3VCoLBCONj6FuCiNRKYF0GlZoGDAN5tBfnw2UmdT4n2Uxq2uSzf2lzYykuddego6UFEriSOxPRV
WPW37GewYoK7wHqb3zHXnNQvGI9Mc3+PawqRkkZMmo68QYWWB8tfu5Zaqr3aZfIrEUmD8qaSjDY1
b2+4G1RVo9RbLBC4bMklNTIexE6zSt98EdinH0EI7MLhfjwa4vEosEm5Zr7JXyz5V0x7+ndfN7bd
r0woiACwmPtpW6VsDn6BxlmzwTTWMQuJzKtqR5cHMfTp4sKGqnqviZmh3iSQ2g6xxhEiHarOHeKJ
nW0R3DPpe8nmfRgamwSEjmDeScPz4xXUDWM2ELtyzZF6VG/atWf0rT1V/pVlB/NK1/1O7JQNrGKN
hwqEMKh4tJi5yWm8s5OLbiYmgB0tERj84sLtv0ipnqosOFXL5C7mYRv9KhtL59Lymm5gjsbg5lNv
Tk2iP0SgF8Y+HkcKB+LU5/5nwWO8/lsSj5ZXIhTD5QCZ0aSHhJ1hTIVQLWr1xtEyDqqV9cgm2jFp
gIgZfeG6+o2cTbJc0BNTCDR+VeKnsOdPEWHogAc9AOwEhCQQ04rvL1132DtBHkG3gEn+YDmZfBZ0
/Jf95ojxwYCYgIdlx6Gni5U+Tv2dLOIwJcn5Ew0Zvst5Zz95c90RlANAeMelGvKbXC8uh1H8w3ea
DbkIsUD3AGHDJ1PSn2bDcJJ8zbkcTx2T/MlH8TmNb0CS5vQWdPQCC7B/eDysWTLPkdjsS1spyXVE
pg8j81eBoPjoG6nRseCrCrjrHOtEQNztAsnZP0mqil8h6W1pJvWWO1ubvERxB1D60I7/Cbg079v3
Q3O4ml+L/X37n4BhoT0GKp+zUCJXnndKII3kqZUhf4WaOlssTR2rlGWyVeksrKGT9bn3IH3tSukY
98fRGlN4oYaRq8knG+D3q0cy85SxbwUtAAZ3CzP7VdZhbH8ybLLjlzbMbqDy0dyJIml+zGr6Zoci
3G5sZxVX/azuVb4iwbmVvDIOuvzS92NH/4gqMpDN2AsW/HdA1XkELoUGLcdD18u4LMuA0pJXYb7b
/kxHoLM6/LanX1xumYPhuq2hnGIirQKbM2ebr+FbzWr0YxXcL71Nhfev/iS1GIrgiyRtGM+f5JP4
oJsqogG912k/Nz6fyWawiMPZS1AeiPpRz1lZ7vV2hDtJUYCVye67zGEqfaVYAyqhT8HCcP3T4vQo
2TyTEfCS8OY0RUAUM4eUCSdVurWkCF4VUNYTtMCXaOJgJEcQorshVGsRtZDLqUcP2yTxXs9IQn3T
81EgrVxEP/EESxRnGOujMsKglW+J0BscAT4q0NscXKpKzjDLs61le6bgcR1vpO83b2YU4z+u1Qb7
+lfm2baAxj92kfNV0GzQSTDU/WFyjdtX91ph87smcjbXS9o2kUEswXUPkhikc2nQHpKdiSFReIrz
io/lys7MxanjDYKNuSxbDv4RE+lHkAw2PqTlJ8ZOK3b9RcdfrPWZomcIqHhSwSd8otaFbJeej4/5
3OBJHqVh/LZm4O4fsmeby4DPlDtLcr8/lirIlaAlstRaZiqrO1xoPyqUyljXPPJaaUzPc0u5eZih
WBqYn0znOp9qlKBuzvIU1YPtZjn4FTNHuN6CHFLc8k1DbYAU2v/Ul5dpyQWgPJxhiiV2xwwT38E+
x+rgdNJhBAsy0pEpMh6AJdk6QcD3jYTrUuMYmDU73MVJqbdzpCxFGjjMqkT1Q5IURLehSfFCcBww
rb4yDoeVWRLSWMJOG/3ewFy1j5z6cKRMgKYyu6Lo4KnYj3MBZ0uIXlWzTqsETzBdUnmCbuOh2Lnw
Tk4EgnW4c5JjCxngCUhBuPO3kTJstERzZQhKZiwz4GJh6/ObWxvogaZqXJkuUPFG6RQ+K2oG+yC6
gUtw8hyE1BywY2b1Iv7AwoQxrlSNXN4d0XwfWJxaSAzeIL0PFRF9JGD2s9siTFxJSECFuFavJdXN
yNjhmjLl8qv4O2S4GuTaZpJ0tM/Z29ZqHSkkhAn6E+7UpCYaVCBJthXyeJ1qXDZ3JQXj39NXTjto
Hpt50LGZbTA4DvoVN3/F1vdkaX8nNowBTd4Ez6W06v0beoLCKzLhXnZym3RlzvF/+PB443nhgRrR
iyRusJFf2CQNAE6AiEljZ98XF+JiueRUoxWJdDFT5H50YItwYByjjdzodqLx1Ft7NPnL6r3AFRhl
WAotKZcIe9q9YphPSPT92nZP+cACyq6mZ9oKn06UBRR5wqaAjxmGslcfqnCZk4PFeld6RB6RjIQ1
dDU4+6oYtVuxWUxRSGyrtlmo23PBudJ0OI1MS8TYCIhBftt8diUP4G18HpvkPMEh1GF0I275IGm5
hpl4p8sKoUO2siThl79DZlSVO0WDglimQ1lu4AnXNsAk80vm77PlIhz3qvelOlYLH+22IkF7+PZu
KETty3o0mV73aqZhftLLXOya8c3NBoXWwze13Lk/nj/Y5yJAo2A36bO7rG/wfh9u5fqLQkNgSXrr
2yOZrupEptUkoPSuptSunwiTB7mM/VinCcIGd5fNHXDLWT9dWD4wzDAtQuy8iFP5/CtA4P528dpr
GMRkd/F+zXXVUrOeZVhnqJhHfjhJl27fnd98hClq5gNFycxUtlFvRzuglWX5+4Ctxq4vNZb1PcBS
zSzk3RmsxlbXqHz2i6B0kaRArZIiScmgaYvDTxOFB51zuNooY5NT3wVDpsK59luFkaWUVelIMmE+
jkZdjB8BV9d2RV/0FQ15K/bnh6r/7J6gKEwv7nzjdhPr0WeT6ciENR/PdfYOeV37arWul9PRPPML
ZUJky2Co+hJ81NRWZGTzOHlEc9hViKcwSYToSZRJNtICNflCMGHYZeyPBBnDPYM029ik5dzRg+k0
/to61N8nqCpbTERHh9cV2x/8tRpyQPISQWNNGD7+3mLXpSJC+4cqQx+JaiJX058dBtnRESXEsb6K
xlqArgDo05yUsDY8a39nxftsR5PdUZ5HM1gwyyP+FPGKhap69k0vzgDGx6Ukog85u7uEaugLtFC8
u52i23nO/HGBeB6cR/uYvaL9ZFrMIY55RHczNLJQ4pB7zFVBJNxAiot2J17yKTEeRgnC8IX88Ke7
e4ynEs5qYDeBvO0EG6/i/MCRHs9wvJVGvJniwDCDMrU7b33wO1sAXA3tpl9IzqkqDxNbGYnKiVfI
2Www+dSmaSxXCLzjtiCL88A7Q3/57A7h2ubfjQIdJ/qBgig/Lwettgr+/mFU9BhGlYLwADuLI1K9
4NC3ppYI77qnsuueui5QwFonW2qdgLzyjQxUpCO8rpSeMG4bZY+AwwqDiVVcJXceh0Df5h5qmYkL
pc2mqgEtG9Pi1UP20LRaTG8UYqBVGpnhwBNIINo0uG23ePMPqhZqzqT1X/vFyPuc7VDnjzfD1M4p
vZJAtuwv6AwiIiuxW/fC5DeiKBVjrUGtrxdIelAlldoPhT1c/wj7yt34CgOwfSsOqe8e3Fert3rZ
H7KFy6QXKuHZkTm5mAP0g5kBhONG3cbs8geq9ijXtdutElaI7LklDcE8YQ6lac0+GDF8JzGU/Mz4
cVZLJBPe5Elzsf4STuEEQgeOuIXzR6OdiigD39Z6WpOx/DRUCcyrAzN0I8dAbufGTJu6omAwb+mJ
4T9dDVGtXXp5U8CBPikf76tYEHt64tmNXcozJRKaYB6hXCfimJ07umhAzKYLPcPHvCYm39TOSaK0
v8U/jFNE0+bxUzm0fFbFeRuiXPn3zxwfu9Jepo12KL0fCRDf485ZV2Q5MGwMvZI8AsosRkgpXyNn
07qM+7awiusAz5eZKNopMeeYqM+CY2h+ygE/1M2GFxW6y8/phuGRDHmLkHAUmYYeNl2l4GeNp2V1
O5+o2Z3xFPqD4EfPOMiehe0Y5ODbDvqaTrSPWplDR8/p/Ozz8JJOOuNc3znfJnygvNXZGop3IzP2
Z2sCj+CxSPw15dmA9lYPaYgaqnrLMqTNLnbZUzlAun3RRWpFYe9TLYMw7f+H9pWbXgrv1cHNNiXa
Wgy/gjKvuYV3LW/vLcizF8Va28Mppo7+wOzrtbTBlf7HL979UurfiDYJTTvRGYg3Fh2TwY/L4tYn
hDb9prm01n0QP8i7e5DUfog5lWTbU7rjwBfWHyW8PTXxTyhDDytQ2Q3+uzSUd3p+O5OaxFd77W2c
nIVX46hDh9jJsGql1dTguXX8I8o7GycAlfegKL50VugJe9bmSuk1Q+djAo4WE9B+s4RrUo7IjO2H
81MAxfE/DPEgJsWXR4oA7dBxpxZu6jKLEK97RqozKTBcOCvsq0fz17WVfJp5TXC7+RC9ZuPaPnV8
db3HX8BgVEpLgpyh2UxRDVmRS/E/t2lopkixDu2OyH4SSWI0xeKHuos79u4zpLBJVKyfeH7jdj0T
VbW4sEc3stFDV9LBcRwCpOMs0vgzXRujbtHLjpnS+rQMOC99hPs6ApOGIL1bfYODughP9oViPTIl
v1AI3xsqdAfs0SlgEMQ4MmCaO6b1SFDHzGxURiP8fHJVI2dUwB6sCVyeBROujceKM4SqgMQY79+e
dKMBQrQIvtc9Qksmx962b06MBQPPcvWsLO2tUE4T0RbKT34urKJ1Z73uC4RN30N3UZtKPLr/N/eS
C/hNkJ14PiLaRD5LYr7wt3T3VNEVqdWH2eVTU3fSqvjoberEJBWOIkDpK5Fq7axylx8OzLoWek6j
qhVbr3JOvN0vXfnCBCjHIgfRjc8N8XQK65Ziwi8PcNXnD1T/V13TjuTj1qQxANWAJ+DuybNj9j/W
bcmcfMnQC7XmRyYDm+5vG4t6z2jT4nWZA9VcjsgYNMxe8GaCKRwkokNuJ2ahFdChhxDfSGfAMrBh
ni1Oa3cQKMrNSATbUHUEfCzc/jDLzzVG4GV4BWn4CE0d8f2KpkXnNX36BW4uznfImFsa8jNjL0Fn
pK4aEoKVDa3msG5mdwzKIgwGDY+XUDsExPD9oq10FL7gGxMZ1RK6lcgIwkpJ/8OI4dr465npQasf
QFQKIuJuEOi2KcfZynnv6ZCwePi3T/hzQ3Pc/8Rc8h99Gl16Pb9bXvOfr877ogTgvC4R+W45QVUc
JiScQUB//XpRfnILXJrkkfuA2Ih6EA4ZkeymwUp+Bnhchk6k4J48hhRgb/kTNmR2wsN0mYYZaP6R
TYKdUYgYFQCSJZ/P+hxl3NCdDSAqGMhk/2/Zdda4zk5ONdHIsUABbMgrPw1zo4xXoAOdA0C3AWYv
JR/HV5wWmiIYrL67yqJ9eoXeUw+C0H+unGf5wt9vVxTUf0UH5+h9NaVd5o+liteXxW4VMd5VuEdw
lQHwTeHfrL4H6++vk7a/g+EUgLoPRJ/Lh7YEb6M1C/gmDrZC0rPF6wC1cnwqRj0zRUZNwBwu/BVy
uyqVhlPB8v0gXGaOJ4SaTgHxIpClHehr0tvn9aqbPRX9uPuK/p6rm1ZTrUqFrZJmXhojT/VbC9qp
DfhYLbK8+1HN5BkKT3zVyaRG3+YwNHuKkOCnGKxp3O97kfdkYhXnkqq8dRJ2u++jrdfM+6EZ9A/4
mDQVZEI7el629Mna/WIYLJ0jWlmdz6t8pzZ65cAqnDdUaC69I9CKc3vE3jIdaR/I0iO11XGqotV0
5XssFD7TDJF611xR+qFvE9GEQKiA+fjNithzuE14djz8x0CAmhdevEyEqk0Z0umwjr3zSn9upcvS
w32M9ArlEnF/Ya3HtQMIkUNbVhcrYhBB3f32JrOCWMLnrT/SDgFXbt0fN0Gf3Z5L5C1w2d97yHSd
7Hd6EdJRiyMxj1rfDzmD8gwRhpjw6Z5diu9ZCJMuQyu+HM4859TgF2sh7ZUZHDeavPtRkPUGKhTf
0iCIlfAvOMblu8lIClFmvcLCAzaHYflLDtiRW7wxEhFrSl8jOpFKXtd5eBgnw2F/BDoxorl9ibe2
5CrFvVDFq2W5CsmM0NOfZZle0C5BPrt2da1g3RogqmeOuaeEDg2Y0Pj86Ewk7NTecQBFHgLkqMIT
ANOeh5rZ61+bnSUnjYdrrGd333khsXWUjrpiP+2mcgLlINGy2hfHGfcvbgALjy+zSlXoDzpw0LM0
PT/Ubs84o7OLVug/GIzblIy964heqjmcaAzdVEUeJgkjvN8xIY3t43tq0NF0YaQ/jQzH17tqdI8i
qv9zxqnj4E8Wycy6BOpnEiS9rCt0We3WjTAiJ7jnMOZl6dPFYX9daJkRs1Xo6mjsTTOQrw0utphm
dKbWKTkRJvCQBKsNPn+5OOrPr+RHXlJqZJmMu5OaSfznfX4jqqa4Y6X4JxaurLlQNMY9Q5end5bp
Du44VNoRAipxipjAh7FpNCYWhix51lVRY1UhOuOu22wxtTECwjjNL0Zp/9GiBXa6AauUl+JW850t
I8pw1P+noW6bi5avLIgG+tCosFQN85mh9toO//Ei+j+d/cryUVsDBaYEszunMS6V/Lpxjed3yqit
BqbdoA4liSpHON8l/OpWeWfDkPO/1ZMGxWSvookHVLGoYU8qxenvLcfBrSeHkUP3IF/z0+2MXjUj
YjcQhGFB6qGjEhYVUvfuYGxWZic/fw0xOQiyz23lerq40xNvu9sMTT+7sz8Hc+qCz6N1Tn8fZdvw
zuow6/Y512crLutN+7WBHEb2KJKOMTCpTPFfyHArmEQgt87ly2qzgduA3YMKsh2KmDjlz3oKasRR
a6rJ+Xn3h8I1Mx5MzPO+ptY52wVNzYBCmv4B/k7V36KHEr/5uUcDzVqXaCpMwlOuf7R8nfuAsmJ6
yfk3zvvIAe6qegqmqM2a3kyhfq7RCD2CFhXRlfRA3C/jFNzLEGM9rKTobm9Foxdr6hprvQ7N7pHM
q6olCqxdhBqm8nJAdugxDcO15IWPQAVDoNU8wIYdJvq9+YVXoRmck0rW5WgKoxrkBJ1LTe3xOMzy
1LjKtJM/qiuf0wExZ71Ie3AkE6WKgh3z3n+v1vqdw0SAvNonWNlYMZGg/THrI01GgLvAMJPu5smt
mfLq++Amgokfm9KwCqW/qgSxGTbrhIXLSwsHrCZ7HYOuoZUfLhs8uS+oLRUztcuXOxoMRW+xaxq3
WU3ULtYQNfkfSL8B8qSPt7ArhftgLK7KDsL1cLAjnV6R2qEn7B2Gn76jfEz9g4egUZmczCeKUTw+
NLZ9pb+zwxrhL4DhJkFdyrbOTVOaLs0pvBwwvEWplYGEsk7ItBple+qzjiqtZ68GRto6tPUjmiy3
w/Of1/a6TnvmNjdCkfAT/EhnD0dTWHoiUTOSxrjBhcTdyQYQ9Z7l3Cwh9u3Jf70MtBUO1rPlfXVb
IaSWbvtJqfYZf006nRA+UyqcNd17QI5OXicZQodYkCdDXzUMJXpdVY6yIuHQE+ORTHBQWYoTW6GY
tu3W/M0zNRuYfHfP4soKIUF7Sovugr6uvWZsLaW23O25Z2Y2nT6VkuU3Jz6fHY+I4lOwDY5GtUx8
HQLir0Ex1A9rHOMfH/CFU9DR/fC7xPKghd2veFAQwHLY/R93miTsgOP8aucLwY4DbQnOGhE0ME+5
qY+jHRxr+WQsJN5HCN4B7JfZLYPxiQErlbetyucpsvaiAK3sWgoxpdoeDgIhwlWH1MeicIRfPgIm
zk/nlb1vDwAHe3CBifsvaa7Rt6JyEtiSI3EKGCx0LZfxEL9FY12XROTzIu0mQLxOq8KWOEpDevQz
P2Tme1kgeUB+EvFAV1rFYhALYuHD4KNp4tNzJi8/CAc0vKfaFjsvjM6AYhqN7Dxy8lkuhezmCiN/
u7csjzgYrteO3y4UnqbhgRIQmMcfZXbfB3Ix08Xt6q9pJzsZx2NDuV3DhN6Fwdt7Svh2cqasPcj4
ncpn+70HJDUGmuwugfbyyo5iXPWPTGhdVJ57G8KdS/um0od8Phgre2F4jgoYc3DZZLB7opiTk0T+
De5VPej8K8aR86OdalCllRoERE9g1VKKsRpsRKBsk20rtca/8fvCE7gZcTzdDpUbKR4dBiyikJnJ
MTzhga7ua/SEnCWSNaS7IZDSkfxbW8KqusWDFy3Q1FBBA6u4vd4cEhFsBFBery1YY4bqwxb0wqJF
WlbvfOPJkP/kedi16ykkQOvcKyM+fgL6osiet6z1UqmGb1vwfQdcmDSqRP3yczsGES2L7amC882A
qysVm63Vf7GLqfIENwNbk2yTrMeSOagNB+e0EOKr4vaioyDEhMC9K9CI7w7jRMkIJwcbWmk+2U8O
NH0YSK6k0PdCG5VGcbU9+9WtyKXAA6xzrQE8TwFMYH2VCrozaoLK9YjyxyX49vRWCXLJeMfJJlUn
r6ZXMWK68b3U/4E+OZmrbBbPfBlBun/rNsIoQc4tUEqXkxFYWUTueQZb8/7e6ZNthuXZEz5bSdvF
DkttdgZzdcVODbpFxWYhSRQHhmszM3VXDAz5PxLpBhU48pu05C2+YSjjcmGAvEK9XGQnfuEEnRLL
3S6pcuYySVDTfg50irjfnwtIEdOdWFO1RQl6ZlgCEyWPl9jfLQSpRpBbu7c3vgaJd5JFIGWX2iEs
FkwMx0+lZY/OMioX01Ds7WIXraPJ4RFjp7CfSs/wv/WV9NfvI6/tqdYTQ8FFiB/TMaeHR3S2EiMN
HkGP3mvgxEiCPskdas/C89ZpqxU7QI4dFoL/NjvDwhfykFRPlgyfNoVE3tQtfa3PxmDjJh3/VqqO
PQvHD6+tN+yVlVePUNj5vkGE96G08aSpW1JmQV11wlVYVwF307Y+DvSGrLgH0wx4JAIXBFKyuGGQ
SAMu9ndGYt98J3WFjS7f0H7QvjS7OvQEUmbRkI8orxX/PAOoLfN7WsBJ8Dpg/oI45qloQDl2AxTt
INUpDLDfx9mn6zYpLC6TsOUYSnmeBcGIrlyzyGxGBspkgXVwQRlCT/lozlk8IqwqcuoUTdkvqbKp
HBsmgoqd4DCgCblMECPUhmouYCKwSQTAsMHcYedDJ0BbEFCcv6tZdN/SvUM8UqHnXsmozPCxusOJ
0TcDyzuUqK34bHCjTC8h+u+0hwGxwMz8cy1tIIw4ex/0h00mUN8WZ4N+SMA8g4I1ZGDJ+DIvpY4L
8q12veNbtk/PJP6/lolydYAWCKsNXRd//LI57W01AA5DpFScxb5289cSTYYtssm6n8s6DwzK5fQs
gfBVNv9u2bIzx+8dY6c3SmcOC2A/LzAOX/yOdkBXG/9it7Ybl9syTvprKmbv8LiNbVOZXWBfzrU/
V2HCeSoeS03aQQOORYRJlWsZmPhQW3JkQhsu097HjYsNm78BNTQjA9gXetcFbhjhf6oScGpFZ+c6
Uci0oQ7vUxMaNE8eoMIHsNrnDr0BhRneG/Q12Rl0z3911Oazx9c4MTpcUCFXAgU0luZUL4ALEwI5
jVdpnoX3hsI3ALMDpj4Ec+LoBkPsKoYndh/+3kM3JiSGAnLbOqZryq8yPAnvAwcKx6o0npd6Dran
2awmPBTQ5K23rraxxWusXntviykDNpcxEmkBVicVAfSodF0YNWAgvwd7JpTozSO4NQfDURNHAV+A
+aKsrHRYocW9n3BDu6SdV4prMAyqr/mf6LsGZA7OS1ciQ6wYOL6lJJmK78yCNQINJQgbW7TQ9L3F
9yYc6w55mdE9LRgjYMK5fwREDStZ/QCZ/bbFtLOVGigi7VSMZ8MCwFT0BBOk4754XWu9U9WHUWV7
c+MgbAsQyq9QIOIJ647gdwL6ftigONT3y+8INQUxVuJpaOsXYjD41WipPA5GxKPRutkHuyqqM5NM
HxZ29CMlIcBYpj7Qy1BAXRtAByAEcM64ln2AnJPCVjQmGaduycGkQcbdffa7eHMPmxzu0Bnel1sl
AH4hbTGJaHUHM5pKGM/AjPNE8jpJVObyflaHc8o8y9Fq+CSy63rwI+43ZPOsHoWNtUOVqvBHDJQ0
ozcbDMIlmxlL2AwcMa+hL9fwDEfKsCuPcXI7CSfX7/wqOkFq6MtPDj0lkLHmtX4hfIxEfd8gAmru
OOlyqRVGXeR21sJzfR/OMo9bXtJWYl11/kVmjbXTxEKM3AAH1RwDyvr1QB0CRmkFqbqNwGSCdasQ
wnPHR9bfKiViU4PFr8Bi8bUrDs3yP1a5S5RwjqvTDQnQaxrWNMJ/AtMLaCYX+L+FvquaN1G2bEqr
Du6ABSKad3JDp5ld9fUhMicUDGsVBqwsc5sMuoapjTpoYl1dX0gdLtWPaXPaZn0tKrhFfdfBcDgS
j2amxhbLxMZveaO225zCc5cX7MVSTVn6fdMp4UtuKn4wMS9HfQhAH5VK0DkNH1kgd19RNBii/+76
S7Az8Dn9C1vrSiVhoIR9C6g0kVxnD9lUbviRyq/J/Kg4TnevmZTSn5p5J9IPYTMnKaFehKINM6Tj
FZWCh/BBbf6UEf+CN46qcoCTCi0SrpwQmSzQ3+bbQThXlFY65sWyeHq8/T4YvpAsbNkFLW3oLIIR
6ktNKXqehYuibdRFczad4g7G8AiugKHqJzS1EMMsA4pSbVoo08JipYSkd/T/vINPz3O41qYBLLDN
ijNZwcoWJOcQ+MfUKBLHEZjbAJLh+Q1+p0VfctE9QmlHv6znXUfZIdS/5IzYYpd9LF6vZdzBcc6k
Lx9USp6JXTcdiWbLwuhwjSWbomEmw81D47L+6/E1AVp6Ly0hzFBHA0FpTiOIzJ6VHzenc0zI89h5
/E1XCUArOh7hRzAvp16ODaHKzZEBElAzr88v62xa5w6SnKtz/0/QrcLrzUe285AEvgqxGcMy9uAG
JYFz2TRqW7xwgIidXBlIjSM+1VATDBDuw6L2uyWIAubKbtK2w1BvN521CqUpY203AlzX2SXKA6Rq
xC7upNrQ5Gf64yIyoHlAmdAegIlIr1n8ZNc0j3XMuiH4vzGjgFqMCmg7KwlAanmZ925dWyw6/6v7
4wZQ6mQ/TmNpAWHdAzXP8TkRy33vyrmHZgHQdf9gA26Jx5SUstCi55wBRYjnVOWSOei5M1vEHsCh
wA5vKdbhPaSS7k16qK2Vy+Nct4jnIhxB5C3FZmLxtHU2AMwS8lisVjxndrv7Z4F3Pp1/LlCE34tL
cIxuq44ikxjB/JA2F7efNOfcAicLGhUXh5wFucgZ6n7y5x89mTockhnjLJpzW8tbGycQ/1QiXqdS
x8LYIp3zD+FVDkkWb7hT7MwZ3hgdKeyDIBGQ/Zf5Legy+UNvZeitsgGX4Rr6DSHuB+eXx+hsyhxP
HVw96VEVcQFKD+RfjCf6Vcvt1d9qvxvYHmPCZq300EGsJJwkr8ignzJjPVSzJAbI7bXNJ6OxiVBP
wq2PfQRkN9uOntLoSGjUsmWdyne+fFM3zLRBXVXxZc8i0vDgfyQ0OUA4Dsm8FimgtZehYAx2VuZr
BcAVfmPWpI2Mbgs/8YMI4RGZ60AFzUBQrj+B6mH1qg+L0jX2oC+/hgl6jRIFYhOBRCrACgnLEWMo
k1jmf26Cz0ePBGQRnRSc5tEDIQxbALapGelL2d4w6ujxs9iZWoDbyCSSD3Yqj64CA2z/Yv23nplr
1Vf61ggYoNdX4SMJjOb2GwyO5nVzO2xpDjvT5PxI4gTos4VwYbcV+/E11LGtZDqwdG5JjmtaSy7x
w/f8AGCn/3E/efqOwxph6iePvHC9Dz2tVLfo75E03f0xClAuArpCfjns6KBfb8TAUR9Ag7WeUU+B
MZjqcpQ/qQSQ8pXGhDbZM3tOFLI74n6yeRxEmmeEaiAxc0AJaJec9hmZ90VM2kRUjIhhUyRzX6yI
MbEPM6Ob+OaGbmFgNX/OqhancU2F1vbWyw5N+xqChBbHjG5/hmv4JadU5IMsBzocY7TnsxFP27tg
sW3MiuCGE6xTdzhmy+gHyoAq5qVKGXqAnfD6AqcYKIacm8ek5ovWQU5UYGzool6kfgtB4WNjZC0o
KXXko9ToMEY2+6iorVtH6/H/0NAUbAhxTlEmG1/i/Kkw/sVn/0DDVt74d9csFnaa6XDK8Wgr1TKb
KGQmWEjU+YO4KirrrMnb1HFo3c7Ee1SRycdDSsO1qNpy5y8GcV75eYU+TLTCLV2hMA1W/RgGPCgd
A2Dopa9EujpuZUagHOnK+yoDiNoD2qm0RZyjwc/akOcxnqll//LfNghNZTjh0oVSVHp4uloxV9TM
9IWbroSHb5FwiabvxWCPDqYNSzXUnl/4O4FAzuMPgyzyoXUCGhZRpfJ5GFaXd5WNXWQay8pJpEJy
lyFhYHI9EeRRkGQSN3jFDAKtEpPpAjCoahIeKrgftqA5Oos64Z/KrVqArz0NFArN5JbbQ0UOhuA+
PPiKFyfrPZXLKqrOppWcY03uhd0PmYj+GdKMbuBs/xKOspCyabyAr1Lys2vqPWGuyLl7mBBOvNoH
uQ/PW9PbZtjzirK25wKxJAAvUaPr4wXpACoGbuZLwgfoiTBLSsuEIFsrGadhcmJGrRRExAl+Uj/W
6bnS9rqsYuS2BjCkM3GvEEYn18GPjOfj6ZOsAb9zUdcq0bDc+5yT1EbSfqNEO8yMsZC05MnejK9v
YgxH4eYZIuVl6l/0Li1lVbmK8WiVL7kd4w6Fxs1GuMYEJ6/tW78pmNmQgWkNpVcrK6KmUAmgLzMD
L5C4a3f40ej6LJbmJ1RY26XtryICD8jlXGyltZO9KUlAXh1K3sib0XriTke6DOZLAjZATHvYD9FQ
AfXhdUL9D9+a/+lQifERlH8mXTBPoA7Kk9VukVtOmnkS3FElb6akj+HU/B17vjzRMJ3Xs+/QyWfm
L01hN+pGFPduxsFxpxcLDgci5QpRo3BdyjkbC6b3gSbn1i13/QE6QU8vwZrql0KJtwFM+lJL1kX9
8Wjh9K4uOMGeJuCgIqeZ8vKgM/VaNm28xS7j8NulbnAZd4OzI9ISdSKJD5+FuSI6oO7xZwmDAms/
P6RAWa7ohJVvk7RelRVLs5DYCzCFFUFuVxAWOp1rgjCdMQ19OiBI50i762O0QX8ICVKdYnz/N4kI
bxX+ByAgUp6XC49KEhpD+lU5SF65L/tQc8bnPXdkU2Bs4IF608xljFXGQcED0EEiuYrxqnRGnBmy
w2LzRtFcp9yTo35e3Xlehv5y8sjj9GxOQ81DqVj1FhDCMnyc6PPLHAkqlAsfnIdPB32dUXMm28DD
blJzu3KT72LE+OrA+Ofldnucny0T0eqehHIPFJFzVFOQK06QjHSdJ67/U4hcEYLpJstEYyGTqnMI
sQO/rbEEUlnK+YUXiC/6alrUT03M6QLxSw8/xkK1eWfyPMZjx6301unqJetRod3rmlRsxXOsagyT
VWdpfk3M0GHiAR+UnXA7p7LOZBypDDnj37QrtMO2lZYe8oJyZT1A4NQKvj0j+AcEDmeKsI/jvMgE
Eo1tn3cERCrLlg8X8MG2HjPixTp8Pfqq2irMFQWMPEgn9KEmGM1mOx8onGuB6DbhO9gP4zpDiVoE
jJUkIEi0nKAmgX05qbJs/3N8WV7xjmZgXlSHCXnCtBl0VZopNLge/JLemTPgoSblvKrAswQ025Bs
fFXFzQG1UwycFuUCUTMnQD51Zpdb1DL3DzpBwE/6LKtkYbWOgClnLgNgVrz138LZbwOP34lKt6gY
BYAGFttQr+Tekd2qhauYjrJsymAB0Z0VONN/FEP5+5LkfhepP4GX/PkwOlvgeOYv9+hGSka2h8H5
9G/T4CZVyiiFrSMF5zdptKQOXQ+AJM0tR3jxQNi1Hb4fVV8MJZf3hhNXoHDqBEuZ7+6Zi05uwATP
vJPltS+HhedmfRFRyMzgniEXFaG9HlhQ589OdjxlpQoUek02+JJf2S6NcTY38UwGPrmpke2e2HYm
v1PlfogtqaGXhfn83Bl13BuaWtfxjt7Vuv1wAhTG1Ks+X76Pwy49AL+zJfXkI7/8kBXrGSiILSH3
8rUfLFuypOuvXLiDiXdI27MaKWiZxKZlA9fyiXR36JnZ1iWLOPuOWj0xm9Aj1YevH+H8DIDO3RjD
gNYivELaYzL21rRbN+axkjtUbPoyCP2sw+m8rn9BA5jlqL3cOi8YkeRmJXQB/nhAet7iFQRHsQ08
AtEXIyjbpHisQTKDUxS7KemzxookDzCbRxQU69sZBuR1I57qjvXjK1ZfxvV0dq14gJDcUMKIytro
oNzNcfloiLSimN8qNijzbimAEAi+b+qtWRw+rqFIoyoVZo7PgUU6bqCEI8q5KgEfLrUhFm1xvP6H
8cQlsa28QoRA0SUPv5VCx8OMyzw5195nSiZQTeUOPgYPnnRTsbKykoMG7y0pIV8pF1ygfLY0R3Pb
DNKQcowXnOXhPoBg+BB2ZLPAOWL+2fcPRwO+qVF8/dUX28v7alvB6irgLlFTbOl9mrnc4Ip5fFem
fzDYi5xkx6sj8mtYatKwM0JRp2/K6PM71zm1oV47tRwml+E9JuHznFUVcNGSlRncB8+Y1rSjvcBT
VxT374L0uP05wFdzJ8uaN4t/1qOeSXWbB7PEcOKS++0jOTsAWytQ7f4YmN2xblSwJGSqSXtGW8Fl
fducHNOt+/q7jDUHuZkv6CJwb+WNpPOZA9Rt7rSPk1fb2VL9gQmT6ul0jPf/KnsPRxAqMiT8Bws0
7QhHMFrwi7tYKgeJYT9/QAX1PUYfm59vi1OkF04565UewKKneB3SrsEEdG2BGXldm7Pe1FVN1IG/
9w1E1MEinxzwUwKvdOJDBjgEpfvlj95y6ttsTWt999cNQT/H9fvwMvpKx/0TEocX3g881JUXHOQ7
gXRN+SjiygtaO9Q5ijtxx8EzW1tG+VyhqXHdfJ+m7j43j1GYq9h5ywnpQbEU5rw9gA+R6vOZWXuJ
fRKOWoX7u5E0YDm+83nO47WvjqtTku2AqMqMINyRuPWIpZNDxEv5MZESuwSQd8W8SKDjN52KtWh4
jVH3v9qI/lxaoZR+R6CTstM7kqJ1jBfFG7Tlb+eNz1nRKiEhlSFPHdJrOO5a33SEnrWqkN/0pxAQ
+iHq6O8o4c1RkTDNdq8RXLRr6xMTqGGP6cqMVxnvl/e6X6sairgmncMYF5rOa3H0YBjkr1RGEJgR
yVa7QBPM2UnBvbekVdI2duaPZnu1R4q9aN1eA3vSspIFc9PRDE5Mz3pbncTIBcor4keg/+34mdgv
VCFMuxLA+KGqJjmLgvk8/o31d5PeZjJtJk5T/K/haR6lfrKRBflKqr7Q3DcYSLUvUs4gsx6eg7i2
4Zn+IAPzikaW1vhB7lkNHI/j12APftxq7pD+zuneOF6D0hm2922bRi8Hz7SUcn8iDYdU2btzWq3B
6+XiAL0K8mbx6E8phmP0nRZ8sOe029ukSaEGf1lhqAuQ+FNJEMhRFYte4aPPVhHTbvvGDUH0SRwH
XNynx+QVjGTVJ37g8uF6i2WbWkHu1sLvS+yrjTUpQppijrcPY9xkQusJ7UKGWui5QxHhFC7YhiD8
zSd1z8AWuR0X167Xs4mmTL7TZRN/W1XiFL5PAuZ5WuFFsflji6h0CSJjPRbsY/B/Wk9zveWzX9AF
AtS6Cuulj/DQ9Zo/TyhWgPc7DMMrlG76WOngpNEhva8QyrpP54bLjOtQmajgaLCkd7QhfiWs6OyX
J7GClAINzq3qTH30cV1w1ecLaDdcGqup/vuGIyHUq4LRUXL22P86jdK/KYNx/pMFEOAXg0nv7hIX
j3As80dITqLCS8Z/el63OSbK5n7WQeXsv6W1F7z4YnHAey0qv/ev1YnKLHAN4q/wGUcf3I838Pwe
zfLhpDi2udrxnbQ730quKWo+xjQ1P/NupWjPRnrSReA7PB7OTRBcuRAPPIBnqB3BG19MkfhAw6Gh
WD8MqTwCRO7C0GM39Facz7jcsZdG7y4DXeKNdD0+OD8zCKu1t8Ai8nsMdEXlFycOTHPmBwl5pGEi
YyPTpbS4doOB+1J7RtT21Opj2RTcZQxQ8ZXJoJ2h0X0+N6FkXPVdR8e14i2uJQLGVcRNjsd5RCSY
QVKcy27Ne1Wb6VKB4QmlOKWieVjarLmLon7GJo5Z65XIzRAmocV6c7p6E7ecVCdRK1bCVIfEYafd
abafpnnbxeeKuDVu27LYQaVjLc23LoWMaXxQ5BeWSKt2RpPkhID6HaQen+h86GVppARFPVNx/F4m
obRNdkPaOfwjEzzLEp7ubhKYm3ZNa+pVbfkyDpbHQfvnyMedf9RnoIIFobieH9LXFAWr//5t7gX4
BEKCoK4thbdPB4rRHK8dKzbo4P0WHoqW8QP2JaThARexgiHL64scZrF/jNO3FUS+mKlYsbdnp7zN
qg2wAEgxg54I8ABv7+JYyJOJ9cJwwQ8KYrattEayHR9XqAxLjJSdsfOicAe6wi1gqpNSy1cbGCN8
iLUQ+38LdtE0jdjELaFhL9jssDqOpFN+i60/yJ356Js4DqhAssOpbxnjVR1AW9Qt1ooyWsivZSwg
A1UYZZZRL2vUGC6dA8Db59V+eLGGXmHs/iJMsdKOw1BDXIsPLvFlu2lBx2HwBe04TzimnD5NpZEq
cZ1SxjuftOgMa7oaH/HuO86+d2qVqrbLMFXxljsTKoOvIMC8NjeOXxZ9EndBaAjgc9UWxb6RtVvz
9C9DrXJ+xYqkew54AuaAGFQ2QQguKSJeY8t0MNeiKh9xUDKa9TDJTcXP+gWWUO+6LjzxUjEJt1wk
T/NCP2J2iMsOQbWL6AogH1m4Sb3MhN1F5kCC4GVunZ3dXzyHFXjq7SgpFAG+VcaOXTt+afN8Jkqv
/y/ilmtcy/3BfuDIYIFjE9yzXWRaori45MOol7WqPGLbm7fXOUWnzd//L0pI6tNmhmD5D4nyk+V3
xCEJn0/0hJd/l6j+UwAoq5gxFgUDIgRhJFKjWU4vMZhYpDtVZJ+vvpnbozfRMLgNPzUxynjbOMtl
4b4j3zhvM3dWqrKAvb5l7EMDjE2KXtr+QEqWRRUuMyZQl4+tD/OtB+iarX1XzTSzimOff5xZthp1
bjdpmYRVuGGxxeKp07FvQtu3ZeE+NpGUvMnN2rrzkjO131lEV1G81gISRwPFSfrOC9/mmweB46St
4W0+qoNFxizSai+GMxUvqWxR0R/OObxWtbRrs14XtD2Eb/W9ejedm9tdfS5uq6gCwrqTOBMWTB2i
C4ya9Kmn4o6GkGhZDtP0QMtPdCGKKcPp8DzkYL2OoLenBqdeWi4S4th0hdkVcXrXrae0bqU69rna
3ZwUiPCByVBLTOE5BeC/HpDxADm6tg3SVq5POdM+zqo70TtGIf6sysHW2w/aOVi/53iAHvNl5ZDs
zyTRX4jCKr1YmnjPcqk1z5fs5GOD+IqtjdB9PVFumDiRQjLr8uuF2sdcoM884UnRZvERa+uaIMNq
JX1KKocYae8ZIQR0W8ATqiqz5FQZOPFZWK/00UBDGs6Ia4ZAQqjT7MLBRikjtSnoP1AL4xA6oK3T
QAvPagsCuSojFj21raxkKHDCoBmGI7DNv3Pt71ho7MBdFJxLiV8y/Ug2rO55cBBJOAN0TuF2q9bB
d4HGaj1zxDS6jOqmio7zE0VWCqC86ZCRNSeWVm9fkwI/yzHn9kNdrfbCg3ePFp1QgHY02Cf/mGE7
Dz+Dl6wtz81cCHTOr8D8VkBwUFjCGwK3+oE71uXtRCc23Lr4oQJEOMQV1f87XaSgdacMawl52ZJB
IEQFY7yUqEa3S84uUAfl0b+3nmfPrvYtUGyPAfq1FYCOl0jOAgGMcQIbivRmtIwXNNAaWZsAv5LR
hWH8YKq/4UEeHDuBEIhxob4j/TajzHsvRa6XTlGecHCh0zeekFnc66804GTnG1eHyd5j6ZtPlME6
TLTGPnayLED9mdmMtERp4qrhR7i7AUDnhEvRRbZCl0uR8fN61bL+Kkmqo4xexAF3VUbl0Dc7N0Gu
5ilzB4Ueeqaso5o5ycc2aK5uQ50BWsQqgwQsBOhtjeW6V2fHF5NoWbR6rztqAiG7zKKp6C4pyjvB
732VT7exZ5Fkv0KPpUnoNHDzZOPO52lNte2V9AjskNBZdnF43U1Bi6WlVdzLu0WWZJbEpGpkOYi1
fAvBZVrbB1Xccexyfukrm6fA5uwfW1SRZBo+PM5+FubNm6Cg8GgeT1VwbcyWjsj4V+PQFLCd5K6n
w746oonUfd3nqZjvU2CIMhlPL/4g6SpSnAoZRm9vuLRP+skJ11uLKueW2v7BZJb23jYfrGcW5qy9
NnYB9373rv3/3vjGSBHpfOpZgLlIhpfJE/aIJNcC2a1aWBJie1xcadHuNmjjUn2NcCst3nqAr8NI
ZLBIeDWT4ReySQ7Wj6lw6YvnsyVqyHrSfJYRPlYLdPMeKue2HQRuaQiZARPPZ3eEZ/mPeMNtgetG
AcDi7rAhsa56HaYV1/C+X+ixXfsOtBBBs1PkgpoWmGP7RwH5ZrKz0y4oCJK3cn3OyI1682Ar9B+9
j2CxZtgvEVilaU0n62+uxlwnB1zPEL8qFejIvPf+rRpGITIgc4i73CSxUW5srsEM0Q04nvCT63Sq
qhEzVkg7+igJ2oV9YgSNPk0OipE22Mgf+LKkyI0oEa+Hul78z4kdPmlzz9CzhsBwGw32BwdQsXxV
KBWn+B0mdTdWWQTmfzCw+nYaxPvlNYFcWjx6LEPBSkFnO3pVJ40pIpQyTbqgOqZ7XSx8BvwCoIsj
Grh+G5dcRP79xrpEbgdDeaVf7qC+O1XxKpKKbKZk7+pVrrEYBihiFSEXb3W+rawSssANd984VMpl
DaMNWC9InI1NXB41qyQmz0tKKTlSEz/PHo4+tKskkGiQrUpj7faaZAMzqWVqp9nNkJ0lZoWB4DQx
IqlCGsa/JOxGjNMlT4CyVnAvLCPw0rXzoR3/lfbGMWJuvNa0gm9HIBjiJ/acJYaBNdIcNmBDttmK
FEIDE2cqSPzqCNMQApt+ivN0kR4GntTPdAVAAkN2ZrjxTNUEwbb6jBHTm0gkdeyry2nqW/vzcrTt
TvTxUVJcTxaQRzI22lCCPOLOkUn2ePlRZRbE4QetZvLoF4a5XYDLREr3xBsvWWcjwSFUqQ4H/sf9
G9jlpo9Dv04H9AooQsnzKPLec9mZxL7SGEO/HJGqCyXz+c1ikIPilAbjBZHUB/OZMZvXKwhh+yUY
ZH5grbGl+aaHAltI84plzD3G9iCPopib2iEV1/APxouHNF2KPEIITRZZRLvs6ztyc4ylAjUTR5bO
/vN+M+HLCZ+Jgk5BQrYeJy/voen/yjEfRGLsr5nyhmKPFp8tpEwH+YMPoYVZRHMhzQoeMHEp0pD/
YYmSIVdMKqe9csTLcgAoWgFIaW5IRzWhliXvjtgM8PtJrQtnEIvbXEnKNoF+C5orLygKbj5jygWP
IB80ORPX7w6GkL8dsssVquwnBBw0r1zr+lhGlxCbZsFdltj+rXtXlFP8YmQEKuFK6QnG2Xyr4+G9
lwh5cGptnQTh1wO99J87LhNdXyRhJ1azrng9A/pXVA3toLG3sAA+fplYJRfvv712+PhRXLcLWSYg
dWYH768eKYPJWZy5ssQuXaJ9+4L5UNU3dBwTD/w49dh5Pm4+gKXgOM85NZMEwKBB3GtRzmxVvQyE
zRqySu/ug7mneQbqVCQG9Kx7N4iHiMtyuXHsKbaCq+hVg0TL7XascUd9e2rf2+96hXpCadMV99de
HSdZcWyeP+zTL0R0LmcAFul7DW1VTs9W/fd9kV0eXCUcbwwkpAgTkM4djUwygPdr2p7VSxLYbKRm
iCzzy13/7LI29Ej8OIDBzKWYuCD/9JO3j9m3B7zMv31K86yk5CWRJZ4EIcjNIN4V/lr7G+7SViPS
zmJD+qcmCJ1Rt9VBapyOV+1NTYOj44wROEDg0IibWbYSATCSW8ymwae4QtbiiSDvYzZkELGmWp4M
Aaj/ZRW2xd8KzWHC34WT/lQw80bDj3rRBnvafdT8+LLbMOF3GATdVWFK8dv3zugzeVareWS/siVr
tUvO4HxQSkZH5NkgisQ4M27/vRzPQDzAF4QfAdvPJGJibMX3o9AvB4+1xBwYmN2OkqwLo2uE30Ml
RH+Z1jW4XX5CnopIeeNg58bp5zImhQpdYF5/TzUpKf0YniotlZ0FN64ZCrZjpfY+o2oyKax51UCx
SZcYcmJeSFq2zBt3/Z8fAn8Rl7NJO/y+q9wXOU8A2COg1CkmdqDokngdfkKRFRMImHuHvvvI6Szr
KvMrAKqIQvSyzxslt/vNgBTnUqkkKJYYqA8s7q2ta3+dwR6bOw/dSp1qd+EP2NSf+wV3cGNbIWse
i8ZimbnxZd/uegJvjEGuRYi7NEyqusfEufsabSapL9tJ4EpBYW58NeHmS70rIfT07iFusUb9PAC4
yTVPr9ztNfXJNmqHqtdRiJO4YVBjr2BOifR7zHoYQTEZMs0xDMZHKNxokIgeyjVSs+A/pcZlreE2
I0uMW8pcLH59hGpyqF0fBFrNUUj7mXNuMsaUQuqNMIL+QvFkihGoC/hrezNa/1hlEweLqR8qVZaT
oZ+Aey6Ihte8mjdBm6sdNSelkKxQ0v9z/dx5VW+ZNdJIWyXP5pFXhL57L/fFD7cu9iF76BGSDs6g
8q7ht4weDeS34/btBwm3imbfKozK4CjMi1/fZi9Y919A9AFq5H+RuBwDxgUDABScShHykVfL4x8U
YEUql47Id4MNUmGPfqe72Yscoo3X1mbehcq37o7dSUv1XSI9e7Qmy1OtyuRYLmi1Wh4bhvrcGAAp
fWmKyjMtux+c5QIV92W5PmPo4wc/AaCvqKYrVF9uDbYIWgSUCmKL+ofWXx4iVmVrDXqFDsLEZFw7
8TcMWlKICzH+AXdR6oMzvHNcOFLipi6cgKYXNsTkd09E/qWSRsyiNn8NSqYGXLC7+ZpQDu2CBh6f
TAety00ReXUH3cCd8+XKI23Wae4MI/fT2/dsaD44nyZsgqSglUsyz0SrDt4MwSTQs+3JRoObCUD8
wD+df11d8MeXbiOhJQZ+oD+GAzEoz2qVTiuQLBsiARe3R87CsIaOIrMvu0u5UoajvLDQrxwsBGmK
5AjLqUiBQYkMQlHA5u3Gwc7FvJQqBhLKoVymZe3O7lifWrLiqhO8MxtYqANAAUsHy9gPnUy2lgZP
G+DrZgWy+mTOMUY+jpsqJmQ1fNU8+pvEjJPZ24sH4C4xtOjhqhyv/LnhfElPQ0KdlbLaSPSP8CQc
fRJbTO3WebVLZaugJ2gEC9TFApwGA6X296a9j1WMUGCOnzHp1auzu1tpcRl9XmQE5rqL577zcYOn
K56IhW0juJhuprMFuhezoVAduEGJa4kd2sZR2qLCMKOShHSL1JOiWF7wbsaQnTX6Asgyw1at1057
R2Ux3ulGVAWj00i6ZNPEhB9iUKMQavViIsdrqwHlqQHkR7lyWRgagCaC7TH81FwWXa9l21ybg+HI
TWAir0IWwXs+2VOcIhXSmyAAetkplHx+2orSULR6IR/qoDuXS/n69VKY0n5cQkeEryF4Lq00ZoW8
OPzpmBPEwOwb0KBWOd9D/EXV6nb/j5y2ijsRo/gN0BtKfDkC6sX70FWWqvBwr3R1bDCxJq1OUkwW
Pxf48KBmmjBvdKwMrmWH9QCQQDozbYnSw8zFhMU+n07+oTKEhmLT1E5ccPYv4IYQMEqL2dFnDlr+
9EBejxiz2pqWb0m7lrEw48z3vLxkYcoEq8rVn9pLC4XRRwuq+aIMJGJD5RnQbKN3BdW/tD50ebRL
TurGtWs+K89YcU2cucjmRqSctcgNeJAbYYfOb1LHs6xn7hdSj11qhoiT2gyQZkHhsJxt3hei0MJx
S6SWatmv6XhE79UfVsHceb58Slxx0TJ0cBd6mp+d/xeJwzIhGeTEdsF5vko49QwYM5WHzpKaELqd
jvErFkpGFy6sx6R/G3l6/VBYYoaIvq6HmIecT/LBOdaYvbdRqrZn7O1aeOAd8VTI+FP1DBro3UwP
rJiY6h97iA0zKgmtChy57j3l5LQViB5DefNE+Ol1FRylApzU7g/1s6g0UbO7awDTOr9nCkyWp4Uf
pOD8p9uVXZcuqu/r/afVOGRpykxw8B1gOxFTJgbM6kyaHg0p8GQzVQP3uJzaYp2CWNQ8CwpPezek
IAYTbecfDyyYz3kx68W5UDbAxFBKLsChOGA2JRjzxVXQh1v3SbqOnXzQQNgVegt6E9N1rDngVjV3
ivjb1UWF8s/0Utn8QU6KXEaIRF3hom2JBSaR/VLZxjn2ZFRBOSxZ28VuqsDwEYa3ZwEjJz9Fhb+4
IkahWo7curTd1elYMF5YBIbAw0ajAoyrokESNwUrrwFZzQ6gCLNCP30PWqV7YjDwoc+21IIIKNMk
UaMEipXiwN6OKijPePou6rMoJu6Rvh2Xj8kW+UCkpMUIcvDNfie7YYU3KdLE6ZkZ+ywNxwVyKx+s
04pJmwx0/j6ETbd1p3s7qznC0WKcFUiE2FUa0zC5wRK8Htnyf3utZ+7/6gqsrVpKFT1jJaaOEPaa
GE7zwgRJWOvzEKT6mFLGh5WKqncsZJoBG/QqNOnH69O425SSaDcMNFTed7jNt9wrLjpf8wv3GD7N
XTc2XbY2sp1oowQxrPvb6jYJXuikD+PfIO6nrjNfhuOvEWjyE5DeLP3MeT1d4MFoHKw5mErKDn+H
Ay3p4e605THN2zHjiK2moAbF0w5bQS7B/MFT+89r6lB6M1R/FJihnT6K6pNKD0R8B5nt+ofLqqea
4AK7mf2eUc+JQokXKBngtnxwN3+PmhXxBRDn79+3LS3IQsGvOkDO5Mv+r+09EdrQyemPyPhoUYVc
Dq2Mc6g3VOrxERdR/KmdOXSww0UBEguG/U2vbxP3mg/CD3SYe7KoEw4sYUnvs7w5Ysjiawib4imZ
4aoFhC/ugbC1cDzoP2v305BWwaIeUUCbY4p3Yb1h5F+VOA2UXPvn10MIwDZsvJBWSJ2J0DYQDfL9
I7bVwmnLp7kTdlJZRNQmjhZ2EPkuYP0+/P2+xfeSgbamJsKYJ+ZiZwRy7XZzhhjkrQIWtH0Xt6/s
+ecJI0pV1touwsrjH8Zgp5CqnRx6ENjFNknclmJGb48uCZRoK9P9iAc13CgsXbo2ViNWW/sWxPB5
Pa9QHjsrUaNJ2t2mHQ7Y9rHlqQHyQCXqgn7bttut8aBE527JwpoE8mO1I8uNw2N0dM/T8shStMUM
yo7jMJIHLUWz/Na+9UQzvbee48q5ovlqSMQEDjGTWQtx6wqnc5zGzW/B8kK04TxJRpSW/cNY33Dx
BMdvUSXaAURDbWmF5cXKJ5fZDBQdqWkGu/av1WuyL+NWUOog+nSGF/MRVSGcM33AqPaF4JEnft1n
MFbmULcJgTWI1sJOUU2DOGiaFeRWNGAbJhGxK26DlgOh4kBlzKAs+vnrXC1gpriQxJNJd3SAs3dt
Xr4WG8YfJDcOIoTA19FriUJaXlppDiTXMopgi2HuP/tQJFpl7uw8I9KV1MEgh0skdJT+pwZOmmNO
zR7WwVSHS6lhkVTCE0r76tz0aqfVpc5eToTLxrDqAX3+Bn6jg2FhiFfDTK5ADlygpmLN6nh0aXEf
LRmeXUnvB8/qw77RYC+Ewcs1SLqoTnAjh6LVbEG5OQpQwzZoIP9RTMiqtj3H2eWwW6DexFswRRmf
ygYj0oNKEscf/2JWoBruBYR+T6xJvvfrywyAMVzDLG3Whr+KWGYVs+ZhIwBTgyChl25kjpr0qeR/
m8kvHGOK3NC+Ois/xXAaDLQCYjezrZHuI+uxsVaH/pxvE3HY0EGy+TftCDweu+dvfDtpbrDmM/Yl
MLpnPauY/PawabCnRn2ZWPqYe8XJOme68F5uFfT8OPp3Hxp/wXEHjNAG+Ekm9OL+InSzLTBMt5RH
9JAXLlI+HuGeklRDnSIjqXtVD5BGaspzBGYw9Wk4TlPkVkTlRrb8PRCBprzhBmG7ssQFiJRVrcq5
vYuCwjFTf6wzn8HnrtkEbLeI8Cn9a1tIwDCOsIeeXxZ8+fKOZ0leDbKLEl+T3SRg/6bEheBsDmUb
r1llElxoOo7gm6xY/tsibwY3CHCXmZb2DEf2iSQFuIOyQ9r3LPHfo6BknJxA85L1MP3lNjiU5ApJ
Vy7SinCJKK+DX8GbgzYEEfOEyq637OnDplTfmdsrP7jsrr3/FV+grGfjjpoJjzzpfp5ZgJ+63OfI
gu/9T05jLM80EfHX6mxmh0W+wq+7zkZrvrkEC19FTLwj87v9u7q3dRRX9sHwcoOZqm4yP894/Lpf
n8O1aOhfBK8gNSgZTtawRaEPDfdYZFXQOoReJ1LjaBixBAsDs0WzmaM7Dg++40Qz//Cz3k8Bioso
fX3xw9ukmB0fPNJ57Mol3qoSUiatK/uv933Ik+vzGJjsQEDXcIzG0kvPUZVVXa92ryPA8YvYHX+I
1wMRghibx4iRtdNEODmQfaNcfLS7mOTMWssKhmwN9EaJcgsx2qPagkCAQ42BXmCPeWt2PGQQffKr
On5x4EFVB5jHFOgwa/CT68Oly5ZuqL4Znr/ywcI49opEAvkQAXJNGfZU9GM9ssSZQgh6UesHioju
IDN/UN8SZk54KrTbw5brNO2nZZdoH5lO5xqMj4R8llnbsQDG4eyQ1oU2xF30I8djjrWo1c/paQfM
3RMuX6Zi8pPjlho9wVKrcOSM1thOsiTxNgBRaZVbLPTJaZGnVcax31dBc4dxCW9tG+c4jC02aBfT
Ejt2w1rpczNGHKAyGjoFTg/xfS1pRXK07znBApGu3BS8zOyVkkcpZm+Z3u/na0pX3NpcSR8hIwUk
qOK8jgpUPXR4k2ExXvcbOrGYjcN7VXMiYleCVMTQvZ5J3DtojKIv00YgdpfxsRRuZ3RkNRU1DHPN
NmqO5u+qfh/Wc5KM0UC5+lhIOkFJE/v4AAbTgX6cZje4J4Hx88t7t0WcDnaPjgIrpD4rcBeeDoKp
AR8wo/qEvS1kJlPVFEIufnZLkqKeyxznVutzkf93FVTHTGkwOpDY23SUi1XhDE3aZGLDJ73jfFeJ
EGjdtOz5/a49UiW7H1n+YXSff1dny9slSJ74ya3foQpn/nB5ygvtBc01IlKSNQfik2m4yOXN87IV
zrhJirB7B2mR3hiAwdq2siVVqFxPEPi8dBTTgSR9jvQ09zwJwmSmjyOn9+BBTt2Eu+zSP1qc7IAt
azaPWkNEMNwqq4zcf5yaI5SWeB4EUqCT0dJY5w0tqWel5RZUuiQRLiTCtueYhe3YJBJRzR8a++0l
RHGEQnclaPaWc+62E01vt/qsbMHKrBsLAK43locAKDhApk2kz+/WkLEzf4M87jH94lWNb5CqAn6m
Z9TGoUPSlgRc1wUQBy6q9LpWYKzgmdsOKrkHaVp92Q8diyj/imoXzHbbjMTU2FDRDzk3Fj8X/OSl
ThRfgc2hSVfP6iJCTzKRCmVgsFGkxLqWVkf+lcip0yjdAwQNxkFDaiqsnC3FFJqYq4xdDrpiIrCf
MkqKxXs2pmeNW47LW2Zqi4NiVB+vLedlQZk2fLx+9wsRuvoY5gcpq07k3/7zwXPtfZajK8+S9yDU
xzCLmud/csHyqXDok7x8cWIt8mSEmTLr9hAy03/Br1WwX40Al+r2ydpMfpXdrh2ZX7ePoY5kiGGF
qrFT4FmVet7ZTRVOfAYXzj1wBYGVateSO1cm9uqeysi0XdiKzX8AMFWunakRMKh+QSnY9R2MZzSU
kd0eRKqf/ztPw7ZHi45MZ3Vr1x2QNO7AC9r9GiU0UJy1I+Wxr9ea+hci+SCMPPidCKny0sN/1rSc
oG9m4/B47EJFYQoceNE8keu9AnorB4w2n2zz1vkX2tCq6iieeaqAfSMpkFrz8fSNi7uCjKUOmts1
FvL7V3QNd35RWkGty+laf37sM3hEVmYLvKjXwVAg9ieERdJUZVfJORg5rdvcT9CBw0m8QZ+H2Pdd
4EHr51rdl/uixmQEMGTGSfvWMQbLCynFQGsXooX7v+HjjR5MI1vGaefBg6ZPv1+ulvBUySUEe0QQ
wlUDl2ytfowuKRAWavD0P2O0DFP0FLyM7QvT3HzU2U3R11cILxBn4ydhEDPwgypF/xC6str3mZVm
XG/lnJSlEmcfli33x0tth3xxvE3l2tM6qAFf4hl9eYlwb2j1fDlvmEkA/upTzRQmuUYws5KEQDBI
etU/XUXvx9bdA9YcnvRIS2il1hH4wTNhfHwfRuMBPQk79+kkEfwKJeL0KEUN0taPsn39aMC6maQ3
bOgXc1XLMxOZUod69fU34yQRcDePWUc+6SUSIomDbIGliFDIPVpshOhccASCiVEummjgOUwKfBGh
KmpryKW/DttcwtP329uzl9Aydc8neZmppbxqFS1RtTtr50sgFm46U6tpIthgNFEL0HPLvZhQAOsZ
aTkI8F0yVp8/X0ZvKAuuOt+ROY24S6I6WQGF+EOL2iidrif4m7akaOhqdodomuRKHRG9SH4OL8ny
M0e8Yj81uVvrphjBBfeYPSXtVlYgpvkyQwiuCQ8FT7Fy0cyMtNXv4ITf2yUY61AqpmpogpwgjOwA
oegRTTn70w/6n4lqdhv9IfyoNWityqn9DlxmgrAHPTzo0EEw7rhRb+nr1xEXYieTmWFvwx21xEYy
pJuFztL+wBUkUIP1vKwCwhw6f1w5CwDkFfvjccNKnszsIhpLzeffDavPvJVRykfp0+AmwvcFGBji
76CN0X498LU24W2gD3ucDOejZPFF8cSClY3Bvzf2saTWdq8KgZwc8MD42mPXe0ZC6IT06ZmKJ/ad
ShZjUhcD9nT8Cadq+hKBSRTlQDW8iYvarTInQe59qqBteAeu1P2++HCp1XJQ4gUx4Kwg+3SYIkyh
FO/h2SZQHM9prckybL7iRHr29O4Fw15Gv6BblAW7FS8KeiqOamWMa+1pn/8O/aAJ/mYpoKHHen1V
32fAOfWxZoiPNswRbbD/62koTgsEly6jY1l2THC5fUrwe8tiLaWx0xbxyWV7j+p4b00K60SuG3v9
uJxxmXXFfgmRaHME/LbkbkVpkIcHNceSczC7TK5QsYLp/5/Mc2s5RB63OykPeu04qc5J8cLZTKjv
ASexsx6XEJNFBg22uC83LKYjyOCIYJHfWOxw6YrBOe2w/fOoMjCJ+YhDoQtZ/50qSf9DOvVSIJYk
aNNtcdN1hTV8lGBuWynNYTjYkPJByz0ImQIb536pfjmuqrEsr2IeIayK+/8TXDrDFks13DsFVMNV
6C0CCltYwxLDRyDEd4+OgfxhbuKxfThP0Fir6wjXWo4vZT23q2lDWZyjfnPTtRuhfqzph0g+iLyX
n+/mtocwfaoMWd5iVcTS2GLWsCxJNGlaA1gGxQYkLv2/xfc/j9aeNgW9JDLGiFZ5Si/F2eKlpQX+
Ad990GmK0LTEiPBymaFnP+aVCNuLLhy6eJ/Ds67+I49XxS9tG5wsxmtXz5N6KUUJxj1udnSiP9Rj
m4YM+ECB6acPkA+8L1GXcVE5IEodAPg5s1X80friWK/hFvIWkmhiZBwGj/rMtF3OH6XkhJfFeaV3
O5WQypyYxa3qHuZh3MHBlo22EMYqYhQNNcygQyZFtexqX6gjWgj0L91T3EMpII/62t7TbziLWuGC
fTyaWXqbMaadmP4XrAjNTgsRu+p01j4zONtRfuWkKR/K8lpiJXmaQwoTn+Amxb10XQiLa/6wiAEv
fPWmkCIZsPOckeJeTvzFjcspzLld8vUQXwrmqFBPZBstKRTFAVSjLe+s3AIdqI6rYFcWBviv3MxP
vYzU8YO7/+0h7SK5pOrz3OAtQz6QiMunrgsKPR8iRSC4i4VPxw64AHrrFhU1HmG/ncII1DqESlCF
PnvMcTpylhjWW7dN7/iZQ1ZUJsNF2GFso+IVZOiTEigV0Q8gNOdFCfsRrv7CkLWJ1Ln0ubeaplHC
j/zm1W4EjCu677qtkcvUoMqJG1iWNGyz5z5V0nvqJig5pyf+A3id+OvucPAUjHuOGHGkcD3QCe3W
HJ7i92wAA08kLqBgXIhwMdlp808G8gLzLZ/yiFWDMtAi8nktoJWlCQvFniA63hm4rH9gYXU+nAhy
rPxOZWH0hszyIJrUvsgCutDSXxjexkPyqfmEW/hoQ79a/N2xdjEy88BFjc7F18cVV0Z82yL4hZhz
rB6j/UkP8uIX/PmaH48e7z+UEx2p1ZzmwmVsQpAkglMtki+kFt2BWTjoRhwKgIl03Mc4iWywzl+H
MaRfqQ4lhWPL2t3ZOmjW4S6aqwFWvK/n5IpMEZNc/5ADNB+ultop9mAxvz8djo/Bx6fJHR8wqCf8
XnycKD7U+d7t2QM4MGpKWB55LAMJZltMPB20tbBPUiOTCyPN2b+JRKQUsWGPfAB9bhoeZsSlz+0e
Eij13H2E6wusNkqfyIWrbp5V6n/NvJFPfCh1dbgBIJ4S6bcOcfxGbuzg4v/BQnoXhMt5kTVzgpvi
mod+EYRdQ7EOJvR0n2XFngj6RyekyOYQy2aAHcRmFBHnQiBf1J40GIOw0eB6NmaSTbhpDMTu6UOD
AAHXNdYDG43LAvvkOGx7YyUNHzr4J7K1MLFXWX3q7EtBobTaxBtetIEGkiCQmihSuYt/3F9JJuqi
mqeRrw7FusW6XpgIhULqdH4vmusaMcV1S4GFyOWKNgbwcH2/v6f0/8X3du6KPtakf1x81y5QATQ7
2cSoY6ZFVBbt97yyQtvneLRNkAp57VT3ggv5r7q/s3SWsEj1xe1S36wdO5+FLupdwL4VapqUAPlg
Y4gS9TPZsGRMnofHISQ3CaeH/bSktZYInK9O7SXMQz38lQUY+SzPNHzqSZXOPEjfLmFYyk8dYae9
lD9ouKTZf7g5OlrvZs0tT1HPM8RttxF9f7Zx7P9/1Ynkuquf8hHnDysxQwqd1p9JrRjvbfXCvH3c
uWuDpU0X1vtpiUVebP45ZuRaV6DHSjXZRXogRx8FxA4P/BLNAPKG6tlJPH4pcQq6Z4EIt0EXODbh
fzCC54bRueVZLA7x11jyLnZoSj6/Dr2JNN48m1mN/jVzI0FTgTqNWu6uwZ+2BZ6Vsn8jGvGU8s7n
fwGzE7z2C3GQa+kk1UeueKMTZRAMQ4JvqA/0iTs49YwZ38cRf37KnJzXNnXlOkAAQUIrvip+GYDC
SFi0DtN5J82NTUXDYGtydkmhD+qTwqcm0m1K6BHNuThTD1kWs7uslU0a0J2lzdadVKfiKOzx0Opq
eaoZO65PmXman5Oy3DiyYedwX1vgZDnehj9ujg76LvLm58p+PrAihWMEsKxr65hvZDfCEmmwG9G9
payAsgwZ0CBkcvQuR0PjQSHu7b4Phs1wED6wEnWxzM08L/glWuLMEH7ZtKTb9zOhR0sstFRA4EWI
n094SHGwq6b7vzTl+ZONELtRSJBu2ncMtM/pdjawfZ0p44zlo4EQwEbunnlPQAYmln+GA19zS/gd
7I5CL5f8tsGCq5VlgnZmAkNv/R60TYaxJR4pdS2hVSG8OzGA5gwq8Bg6NkU48p/ABwtPdGABiiFj
itc88q9DhHjPPEyOS56p+zVwEF9S9ZaPqBpcrNcyvYOUoubQZ6zPEhCy6c/G07/JD0X03LfAFM3w
qDZfs+/i3KujAqlGYgm+G4Hz8rkl59xDgczkYOKn8PUjsC/O6jacUNU/UBgFTQU4CRb5qYu45WFw
umcAB3hO8X/ow2W+g9sRxCXNvAOBtaIHWr13FgId7pnX1W1nvHTEsU/SH4YkjeXsPmvWREOD9IQM
Fpm+3gBspkRHS9OgHUA1BumRoHLaYRP4nMZLEMIMAHhvpOSkiSWneCkVjrQzxclWH3ixJDDWXL9h
jKEAQeaA1dgQ4PDAShpWddMy3QrcA7n1+2Fk8QICf5AKvx3qtd4YdK02dn71sVHfwcVD36rTrTRt
OKn9WnwjOTrMT1RubQRpUMlS/NdovVcMfOxD7VqVg809fI/I0fh+MpyrbsTdk5ZxGWOIbno7OGNq
mCnjBGEC/juvhQYaSz1Ov47ckbF+622yi1RwXVMuJ61Q32fRPFT6EHJQvkGHjybFS0AQGBe9iNHn
lygH82l+Jm5dR4Mgjjz51W8AduyUNHzUSeEfZDWs5P648HguNhIIJadXzt7lJXj31ZKpXCbacYbC
nqDZIvuQNr6z29fXToE2/wpIMeJmluO9qOf5itr2lV9lVFzxISpbT83TIzN5mcLCWT2aY7b9zx26
FqpvzJx5CYlzWlOhtW7ZnU1JOnsYVM24q4c2yTqw/xcCu2juXKsrKTnUANDM8sEgNThWjzkMiBDb
hXw8KykyDse1MHaSrJarS8HdHpCudiyKiJfCqPfKhmgE2far1yIQQ+gn0dQISoYxXOK52qhSDgSF
3BYItLB5PzRlojiH6ZNx/nFpiVt5GFoM7AAdj1Hqk3ohXKX921G8/xXROoI3YRvSpzRB+jYDRdP3
kzcQu7GJmpElwiNLJ1vUnbk1qBYM8013cap2W0FEG6Gk6wRK0N22kPAXoeHsxCydHYnSnfFZVaIH
O2Lvttgam62mE+3l6KF+U/dIYsCeP4MupsIP+Az9KlE3N6c3kb3Usoxf4+1/FL5YH8jMXX6SddCB
KUACjjNFGi4gv1PqDfvNJvc6YkCUo+GAMRUhWjTvAbf0QGQXis4wUiu9g4S3sbQUzaWe4OLB+iP/
ULUSu0TCMSdpvN7vbogH7TQnKifO3oXWcec6F5nqbAUcttjlwyQpIxkuHxwxsJ/CA8jEf7e0pM+d
aU1emPvxBU1Lv8caVL/cYsH0B2c+QDHeMFVyqsa5g0iKrpZYOACzpTfUi12Lbc0Vw2DQSOlxY63H
2uveMADR7WwePUz4UnY7kGBO7o3LvO5csElgtBP85QE1/AWbnKYWnYsUfvitw1XZYJ33/taY/je+
zPZpSOeZzFg9AxUSbgkF9HVs+hik/BJxhffdzcNcALlzJ6gPxzh1yioSJJifBKRQ1REDa9jTQ+Ar
yZRzFR8mPT/3l6UVGSFF2HVh1N0BOfgeCwAspiII99oke2feAzKcLoh+TyDU7qmlyJmmkad+gKGP
2H6ylOCI9ADRb+N3GdFjai9WfmSzkG3f9e/DXPy3Mtu1nY2lB4/pTY9rPmwkOU1hkg4D/mnPGWGp
uUfAoiegbGztVMlj57blpAqdUBei4ZreflD3m8y2xCIUvNQ7IH3adjoieBw8Tw+t0yduzYk6J1rM
Yc5bU8oaL5Pra3+noljg1krB1wIi4raKnMa7+EMQwJ4WSC5lze6GBBEgT54yaHP2zNdZ1246b8Nq
tnR5oWqoc7IZ7F2znUnMZgtsfqjXKNtOJN/tgoB096a7bNz3bCfbRJIrvD+eN47JPOZsRDej62z9
IAdhQLP1ThaCY8kn3LFYa5wzR6rUQSIHZSCRDHJ7hEtWk8s2Jrx/Wd31zwdck37UdxJi84rraY89
F0Fd63w3UwjtY9As2SO1A2SfO5OVjG14+kKEjyXuflrjZ/utymElmMxUW5uYR6ymHvV+TNAFw/ne
ZHfWxAQFtoaxf7eWv5+n+DYac2qYcotJqRIu9Kpbc8vaFVCoyorAHocS9hGQrCRXU326PiydQUlw
ALjVoaeaxiTXT3sq1Fr6hisLaC3eiJ/mN8jB6Yvu4clCZge4YVdeeyCiQECL7nqIazylD00G9R7L
6kIBggkRNh7SoSJ9MPZ0cbDWyxxX5f/oWucYZK81hlxgT7CYWziH7G2LdUZuu2zCCiAR7DRxQOzV
5RCkDRRRRt/tn3DzFjljcfMnf7ZJnuz+hfL/Qbw4d7wd0Y2JWZQPXyDfFTE6O/cSc19KCj9Y/7ly
3TQ7Y6WLu25q67O2Ve+ci67096jOBj9jADxRp2jWV1iI1ilSqSspL9HFKDMQ39Os4Dzi0vdOE1wq
CWMd02X+GsULMpyEHpsdCQWp8hfKYHGv9zgtDulUHCRJ819JcWGM+GPINMmrcbFq9vjjvL7K4W0h
DmfCHEwJtqejmxB9CFCRajnmlZwtLlshvjm8dN+8twUykUp4U9q4hRVFnOUg3a8qSpIlbGcHsLH9
5SS+73OGkgP+Y33h+caspDAW2lyo54Z/a+G+7Pp3k7LWNbTt0bOp8wZqDMgsG8elnG0SlCUQy94b
CwhBZXALSf5pnz4VKRh/EeXQVAEp41/9xBVlLuq8FseCyf6iPAffDsT0Xs1R1rWl80NVurxRik2z
ttJBPahmAKzQvMWy8a0rdk7tn3/Uvcf3cLZHOeuw9R6h24iKVUNFPvxW6T8WwnX+ti5RZ/38Bwe5
N3eSwfsD59vTUHyPszGS58v8dWt/fhPWm1ztp2SUX/oqLPPcA8io7iWZ4TZxUYidF0EyaUbbRO0u
tC2p3CqfVXpKEctGmLjZ5N2aDGPLHcZU5hsVIU9AZE39qT+W/ekjeR9WWsC+hJWc7o8TpKq9fJpA
jR/7s/xsn2HO+RziifghuW3aHt2x6hduGRYzMrCxusxxyj6Fl07H1oMutGuDYIkGBNmn7tyfMvBG
rQNMAqD/kMauzUrxMjRdLtOH1Ghkyyf/iIMETuEVqy2F2HuOr2ft04pPlpW4osO28s42mhbnhqxR
+VPAS+Piy5+Ocd2g7O/xPZ9PVAJIUq+yE102mtatH9WXJE5KgnMccJApDqwIeFUT78gQH0cYlAwQ
pG0PLf43wGi4ZC0vDid87EvkAs8bAJU99Emfg/aoKZwQX8HOrvTl3R9iwxQ0KfteCTvAjwV4cPbK
7/g5iQGtNXJ7NfV+KcAhxaH8+jvj9LBBHSuFDvrUj64C9eBFM7g5JNkv4X6qdhLYU5fQAAfqMl2i
ZiXn5AM7HUarghVZ7A+t6O7NifePI+AGyt//9UBh4HVb8A2UplgcFiVroHLI3gX5CnkVaaw0QQGw
3892mGiifYEivvdrZfdIqj57HHQWfVcJCEe/rzm9EJpmZqlW+21HO4ZEIZJgbM9Fx8gsymuTc9p7
7swzeluovJ+pKGxhse4KXA5XwAG7FySCm3OUKPrvVinbQZ3YgQ1pZ/XWsrxdS7pneQb5ak9u+C8Y
DJYDgOlnvjJYxv33zR/tQDi8Vcqbyikl1RYlxk1KOMSf3JfgiRuNXKNa/qZaTb9ZbKAJzcAV97sG
E8UxXeunCPBKVFL2jTfdefhHkzNXpjJcW+M/qekatvDuCOQ3D2PO667tGIAjUqIfdFm7aLgM/nil
g8D0Uc/ppXoOBftz4AZDt7uyGsm/tRtzrPLXUulpwEWF15fynMYPPcVZQy5KvmZJQ4hcSmUMS5ey
vxEIZgyYSWpI43vh99SL12Ho7/wFn70FcjyKn6r8IVnKHC2ZOTOg1xqBuEPmwzLGkda8tHwhnr5D
umbr4rUtlYqfmcH6sFnGS61SB1mTG38hcqW85zSnd3eyKGgLZQrzlAhxW+G7ZARrfTW5LSC4vFAZ
aX4ANzsIA9SyUzkGXIJeZdJEAqOpC12QYoCoQ1Cwsn4tSg6DWbeOz/cs1YmaFhOdCACqtT/Kptz6
jvUQS6L4+YlPp6bfm43dcpzW0e13cONFmrvzwdr8G2SV/x6/Je2FAtbJilqRd8RPrr1lD/jG3/Xx
qyVZXHpo9AQn/O3cd5rDOGuaRb1055AaaV59PigYfkeDxdZRhz//HzbIGSsHTKFDLojh5ZwzI3mM
0lo1+Sa5sJMKTdInMfmgNI6BiCTKTgeB+OYAdveD4M37+2/PUm9xOe2fIGodeMyIWOITOJn2mX0r
61DrlSJ6Ao5qfGtGng5/w34QBb4qkPnFHtGm5tU7HOWTPq9SEACLH8K1/8+JluLUp+MuQvo5aca9
wxz5U9DDcaZiaI9YRI7XyAU2QGd6eBi2/WaL7ZNmgqGYxdb+1rWlIgDoZsDwq5jlgm6BO0PSpnl8
IOPyCK6aYnZiV1pQ/2fwfPZ3M7yz97hiA9a7KfetTFYWW2uMB2Gb2WYVYwP5VgVshX74e+GgWKGM
KE3nJ0WUZSODthQNq4wQ2fLGDQYBRUPebySq//SNszKwK9jMa6L2X91xDvre+ysQ9FwYYL50l3t8
l6mhEXngJAzdx2/1ix1smr5Vb+iiYmF1ZGczyzluBPxkSWvQ7diVgw8Mrf8PO/HRydK9xMWc8ris
qwqHpYtpR4KMAIEoEs2wlOYk3+F92dHT2wHYGuEiRPaHDXpTXeC3mdTKzAgrT1pdCsvhPqdJBUbB
AgEvEGQveNLdrK8BSkbAnbOJ2ZTIda8X2s3hUFG2iYQ+/yXiBand86LPar6/P+2xBeSmDkSVwv3Z
UI/iAPOOBkQSf1jzum1K0r80vyktkufEU3Ne/l8yb6OlpdiafnbkcNz4cC8e0+KNeWCzzOtY7Ljw
ZHaW5NWKn7hgn5SwkOLdEB7erR4tVajk5tTLw98EDUcWeSYnVLd1Dr5a/QHY0bztocEGq1gQoyD4
xRi+XWvy2SvinaSBVXCOFWtlKvD9EGcomqbb8Pea70E9L73eP+BHINyxm4wDagcBgqdj4bdddoZy
QLePbta22VQDry631/0vQhwkdA2YpmVf5qPNMwnfTaNVqwARxO71UqxdqatsN1pOoWpDeaP0Rhcd
PWBSIsuQHqtmnPGvOWJqkHSx0hfz3sHsLzKwE4wR2TAzHEgSjXeemZbg2Y5GshVlg0Z5GDV1Sg55
G86RmT0Ow41zYXa9BR4mj1hum90RujFU27BjvgpAhPu15f6p5Wo1Pj19X2EkVslIH0Tf/IzYB/vI
2j8MSAIYaB/fpLf/9n/r5KtNDcTOGp0bawMxHFfKZBhJFQ9cr/CxPLpbdYjdGU2aUUonMe+8yCWB
spLMNd2GotOwsBPJGAnQTxRPC4V7ZbQvdHoUjBxIHAZHZBB26iVGnxWumVvfWwmcyPSrlzGYEtkB
k7XsaY+NEE9/JWQu3ihKJB+j6rM6N7rQMQhQRbxhsvfBLyMu+x8dsXmV4BVQ0yRDojUGfZ2lWIcf
7EPNIR0FdfE9STJ5cJE2emllO0tocWWtseMoBsmJSB6SE22E4q4clh1Vqarkbk0eHTAWH67LQq7M
wmcIahUeYrXARCrD3DHYruO95g0daRkDbC4gPx49lt+rNXZSGc6d/6MUIOvNsA2Tt6agYjLZmha8
HpMZ3niB3Yzq5YYWeh85G5IUpXy3Qq8VI0MDpyEknDnAANuYPcbN49OWXYJxELo4d0Hv5oc3sAqM
0CIKDO1RycKZGsxVsNn8dzDhTsypQqjTfYMF8oK10gSJlstGGCwszHk6gSGQDyq6rA3tL4ACqu4m
Fz50ir2n3EOB6YNPpwmDfsOSo1ctNdss7XaZgXGAi5mPOz+tRVT0YafYIr7bMupW+2nXqOw4P5eu
iGJ0YTBtKgucSyRY8b8uCbvyHTtAJsHOgi8UkYNf45zlzMBlLApIi/s6zlKhBybCx99A+y7d1lov
Ms6qvlEwcBMrGs1yHeqkNke5Q+QID6nxPzveD+J7srts/N1GqE8jo7akksmkic0wtPmW+u5h2KG9
tCYzgWgrpObrzebg0FJ2eFmUOYGqjQnqi1ikgmFlWejXt+M+DjHiKcIItuUyHl3gpPJfLjv14CQT
+RO29Ef1jISq2jvUUNsJ4xX/X0fWbEBqy0bcxfUz983JZ9OsgZPB457qupn5zwZGvwwXKLAmEAN0
kjqIXSTpGnOv36xHSFNjhwL/VJCZjanr/yJEp48YTUlJLiTXUrOWeMEqU+tcRJYEp9psDR98YhQ/
Q8PmRmyEFNg9kveToqVk+4XD1NBAtl8bpfcBWiwrTcZUjFDckvrP9NPSGimSIImK8VgYs0Sx5I5V
Znp/6e6sSICtfi97XO/+SMzZqHusvTx0xEmuwfDCqt9jYWkTcMvwSvM4eY8n7Y63w4QysgWC59rs
zwGJvmETak6OsRwN1bYlh8GohM1yQMBPENI47Qrae/0+UIew3CPQci7V/vEvjLU2I+iiwXNlCMFy
aNC4HdSbkDpazm5x1Fme7yvF0AJ7wF2wRvc5GG8ABBDZgajPrSgIxAtZ5OJVfRxONYicCJYIvEOQ
vFiZTzTYc3NbpWQ21J76X9oPVyqJosTdqIW5pTWKK1YRT2hREJ9pSRljfKDGCD+SR+cCzUVo7lto
BgrudRwssiYTm15qKYjSb4iS/suFwKwXOx7dZ4k8Zy/YrpH64D4j72yCPREbma59z701oIj3c2cc
jEPI6Zbi7jhYQkgbZ47iEftpgn6+asdf0Ko3t485w0m0322l7lczx3REBXmE41ajHc7wzkpbRGHo
qoaCCjY5E5pZIZ3/urOFC5wkL8ec9Dx5+KnK9+8xPLNNmt4OXM3WAUot1SZWJB1g7cJEENlirW2w
vz5jlhuevtmwHyN8CmvaoE4O6sdILZK477b1F42I6Qp1nwakAiwT8wkVw6J8iDIJllO7aKA+I8KI
c36L0a0plXeERMNuTkW5sBRpzMkflhCxjrtt7k59sCC+x1peOIbNihElCdkwhKu9NAT8K+CNVOwq
RiC6lWjz+V4lbl3KhM0DgCjkmyLtmgNlGSgEWSkxNr0r2y2BsFgXPLpqKvVafnzF5A0FfhvhsXCW
OKcKeffEHA/clXr5HggEMuLw8HPHYXGzCd0D44fnIMn9dZOBy3OJ6W4nxEe3fm67sfDn7g5AQajt
soEhrf8ACi9fjHbwHIjzEYyLQOympOM356lUSpj+AmGm4pK+pEyL/Pu8mjaQijHMtFjnp964A5Bt
80pqfUrlw8wh7f1XCiWc+radA0HgNhSIl+zLNeuwbh4YUYb/9R7nvr6p0RfOsZ3Fq8PcPn2U1oSk
OeJ31sl4gHfqYZRbHLtB90Otxv4snGvOhpDJJLIO4hPcxocJqEXXnAbZhdE/q2bs8aaCLoniy8xr
lnezoXlUPucgCunXdGvqQK1ag8wOvVw+N0ASkt8ybNpX4HSiVyZcBDY7G6NEu3M1A3mjX2jnH7P1
anMSkg3OFnmkkzDIiXjIMkuzYRE3RbFchJbo21yo19oEZsyp0a77yKWEfCYRmJxphH5EghRRL/kp
kzHtw/z//WbKo9Sm4+Kw5u22hVUMVs+MdNT3PnnomBoWsrlClKNxpwfCBaGB2Je5iuRABIxT8iy0
5E3DMFi/Iz9EHedD3MXlEmT+pqd6SHbUQSXeUNHhptDDjIC/Si30nUxDa9b5xzRQ4+ChixJwp3wR
rnOROEKDiD/o27lrgu8EI8L7Fvs414pr75qgq/tgZR31tehnQPM0ayvygAZLm7zMKogCCOVVKu+A
9WsZ8SjZqodfArUA+4I5+fyqPeT7+NGdf6x11+GLdwGYT519g+d+9N09OZojXtnwksizHkhY9rD5
YnBZ6gNdtXVOeAgiG91AULX3tm8KkkjKYGiJSc1gAUI+zB7H3Ut3VyXpOGekrlniqVKWa37Kcjh5
fp/SKQMmUbRhjE/58cMCKTaqr3Kl2HIb5VS5vk6o6G6V0UgKmVa2md/h5o9bBF828Y0U2mBGhlOb
/75hsgI/TwTXqoGZSFDIAVqBiikNkpFLsbYUw8xMiUJgOIAByr8Gmcka9XyyLOtqluT631ew757g
bavw308dD6rEx8/7uYewTWfaXAbn8dP3xMBPBzfpbICeI1Cb2t863HtGCrhmF1UgABhXRgkVv7cI
yWAkRpbI/8pNpCV8Gr7wjq3GdNTVNrbUcbyrIRZwDVqsux5Q4OcTbvSg3kua5pzfeQLtwCVwwr27
SbshrSf+nai+sEMFL4/2WbRZSuyEq5eOWYFHpHh81tG7JbUP2+I533otoVnhN8GS5kzOH9OVsI1X
l7mc7R2ALtpuN64Wn2MWoDohaqlrwniLT0vGWsPuEZymuZxylOa1JeLbzJB89VYsnjWiUw1nPgMy
zSL9o8Hocll6eGwEK/2ataVmlIhZt3DPy6rX4Mq6/tMZdNKEQ2wcDPowd4eh+iYCCfQDeBuLFMjG
nyCi3acoC2I3+qYlUMFweuQNCxFhXqMsZIfxb0/E7U9E8op1u6XFDuc3+YASb7eoTLYO6fvafuSW
zWNf0Aqy5W4RqQx0NoKMWkO/ap3ZK/+5n1GMda/KGurd+KdZKIhHBJ84qAxNqbBZ3DN63h4g/hEy
K3XxLm0ZFuBaUSnuRq4YsitFJLSwAjjoszrmoyIZ4OG7D7iEmKY8eLhqzIj3ij4xP9INGD1TLFFx
+eTwXlSnFWfnzmNEQYE5dsUygM2ZUnxsnAQg6iD84SiRdkbhpYMmo/J3GhRo9Vo4yQuhvF49EfMb
B7jaP758gwUKlp8oCXKoCSZCcqDTUcXsSfFsYo7Oromqy8wPOhlxrt7s0uPolLV/XNyCQ63O5/YF
BEQ2paFRCQpv8Ur1E80gdp+S7Yj+c4TrAOOpjKSuMgoAQRrE/4tLoKOxgjFkw7bka5NYNCo79vGo
dLkaJJ62W9on/J/yg63J5sl7lxHUCjBbJ1VZ5k+/eiXRKE1+hkVu5IHECTrtmK6YhyPqb66VjqMK
/4V0V9Tr43RWE/Z9eF9+Nhp+mus1w+hUhE0MbhT5ZGU9SL7lS6fsXxP5OtTKH3rQBdMLCSAJK302
vj+UcoRxLVc0tO5VVlLjnb4Tdj0op8yJpLzyO40f45+YhwhbM/xZMncdCNa8fT53ZLI+wRsERM/p
JwxXzxB4lI5Z22Z5PpEANjao2GLEZC2+811liCXBYX4wg2ZoTT3bakOX/YCranoNjKSLaGacn+al
UiY1JC/Vr5d9+05xAdLvBMjn01vIGCu0xPfywkptf8/h29nyMOxnbVr7uGuFnyEb6RT3pjCzuY6i
O/+Ws2J7KSUzfM0v9abSMbinZIXKIIee4IKuQ8ym7ITLs5tBSTLEvkdp0eC+HyogQBiVf3PKUT3U
QT1eSKCeTOA7/ZHBmTB7FPshQPcG7om+RIt9oJLUrWzZUSV/C4SPcnn+stYTA8cvzaHHQ2f/dx2M
O4C5lJUFrNA65xwklh/CrrBymiAm2dkNxwIA2Wnc65F07CtEhm+rsgDl/NFsU0Hv3GRLWCup5U0G
7ZEWC+ftAQ8dm7JrGUbRVy0qWaTz+eAl0eKHWGHU0U58VsntP5m8loRpCStzpr06whvWizzvnjBS
IZG54fINm3YpE0lq6DYyoXSH20cjIxqQhpHU6ZFdWRK2Iuc1S2bRDJ++LX0UpU855PSguCqz87cW
9yPjvYBkZBXsyAHg04HNCbFNDoSk4p/DKinHDcj4If+qce/EWoA1C7J7TMcg6NtD2ET5k+iJTgtk
rJjUtw3bNusz88dD5utTsgdLB6IcO6GlaIo2sq2Bg9OQU0wyDwbkqRlQyq42KS5d9l8qQpqva/Uo
eIvA41Ecy63eAREvV399hUW72WiynGwhX+WI0c0kFlWWpgr+YmKTEQHFWIn/Lf4NQCoHOoManbgJ
Ezlf216v+8Ib1Zfw3qBr/LoAVZiKbF8YSF3sgsptvpKlU+qCQ1fc8hmyh+qEIpTkhfbU4BpjuIHS
UQtLCqSf39mC9Z9+9F8eZL13ZjXB6J0PiBoB8c7aAFEZdKG9ejC02hEUE4f+PZk/XkVdngHhnDTc
pRnOZ1AtfcZAr9ZJuDZwwRGCHFw+yyLuRqtB7ZVQvEFqVrCxIEfDMWXakc+UtiH3D44Er2VDxnCa
IWPpFpwDzv6MsViBLOoE3jOwoX3IRqLbdWnN7cMXi+hJksWGB44iYmNMpMfKS8wGoo5TXiRieIUM
SgyEGCZRaXASoiM/jnPy31UexUGu6tDuo4/Q4m3b73ilFZw/xn4TAmg6byBoQT3H4D5JkRtS0bX1
eo0WIsWVdRIrPICWB4WBQHrR/7VCtzDbpsBq/OvMZ4vIjs0ElhD3p0CjqsBajE8gz18VajJZR6P2
b5oOsxsumMJqvYQwh6gTKS+X+dNUaVU66R2kidWmqjuPMicY2bm1lv6j6/HwSsMlYptQc3ogVVb1
PE65vmNTB3btIz/ko5vDbQmNnzmFO7TY1NIe7bUA6c7fLfXq4YNl038OG+P77cW8e2O09Q95411c
TsvXKRdlIqeuU+N0f9sjT5gZgEwFUOsXSX6jy8i2awnlqXnwGFpKN79emJf6MOFaMykEzvx1yrC8
zVIivsgrkBX30QfUk/J+O+ARQFhsT93wlNyv/wlfvTq/rrO3w4lyPTmgToXmiIBMQ5kkceXWKpGu
1tDnSa0tt4ERBt6zhuJt4KowWITQy7S301EwD8t7ia4cAGfGAUPSiNiQyIuvu3yg7Ja6a0QRaUj+
Zc0T8oiBKft5lZrDVGvjaXzs6eWtoLEri2KQEwL/sydEfdzahgvfQOO04+ugYeUmi0PJSoY8sEhh
SdbUkJrRU818yBrRS1o8Kch6DkSNfjI9ljDpObQnWRO11QJvysKJ2cac4dC3XsDVrSBsZ9z5FZZS
W6RxiNDv6U3jxeH6F1Qk+HUmbn8umoFu8Xrv7FFee1ADLFOhh/zm0OFxipQ2EryyGTO4uzaMQTz6
Qa73O7JKuc8pEO5eSnauAJPPhqz4ZFIFIPeIjR6vu3RPvmYEwA+zf2QmyZgoptXB4Jn/Y1EH/5ay
/WD0DV0Ooid3Hk9zDP81lKalklYJMyMitsXRZKqWJST92AMqhKplPWqTZlsK7q4ECx6AMv5vfeMy
nPqxTA0TvzsUWSYBM8OBVyNTAQMIRQbT/OyPCHvMwqwWcXEComanIdB6mQfPq4YjqmQPuCINQbcV
l6AzLkklKOfFA5luYkBbP/3myKHn/vgvKsjg1lymj8/xKtzwhN7jCEbWjjNyUVz+QzxJn5ARUmJn
iLJ/Smq4eEmkNQZ6Xbb3C25oabxFgJ7H9DwrBl4GoJOo6mz0XWSfS/jQrdfxzbXQW2TCnaYjCDHB
/wFFYFR6Nj81IRyyCkU1A9AkMHvrEP2XFbFs/N8F7UXK5gzPVOgwRdc1ETTqvTnq7SlBOCbAn8eb
j++12l3LLsql8WG1pOgVRlc6PskB0iqXqq261RtErm7n0zkTbhv1wv1u4inU7xxl74NMmLFJjZg+
mSk2mwRfC5uNLFyDosgISUVdFG9x0N16xGjs+P/krC5fCt7Xd5aQYVPfLZgJtyMMrPI2hKLwF+LK
8f+mt9MqSnCgSrdSqiD2RB1BejciRsaZZ/1zH/kuxXjCNMEYsM9kJ54I9zCc2EctS/nnxT9QOdPf
Xa5xpGod/hcHHFq5gCrinRM56H6P1/lLuu6uTpwVNGKayp7t5jPZB1WCpgi+2bADwLYRxtyojgp9
K7QNN8HxBWaVYbIGMCjDgSemBDYjxLweD2wLydFlzLCkherSiQhdcdA1308l0clNWDGCGWtDIVhQ
nmN7vw3Z2oD/pX+Ugeqyqg3vFVxYG456GX8exvIaHFVJlfgWDmXlzKgf5W57Us2D0T1UK6+cKbGb
OY7l1qnF88sEfBz5ejmpxGfjyqcxpBodQLY52b8kdh8HzhGrNbd4HncWzfPKgvwBzBuANJ6dezfO
cpT1wi5P93YyQkboWCHoyjX41dJn576dgQ3RTwZ5V8w6t1Wapyl4mcrsm9fA1nFSCt5y+oASdrTm
eNuhPdgyd+dplVGkcaZ3kDZT7B79G5pQEpsnRWX1JydzHEieSsJxKILL7NZkaXICJ6PwgTkW5ifN
rJ1qch2IU35xWZJ6pi1yt00ira8zfXofYddWnESier3Sh82OOWpbIou2ZrnYaD6pi90geDLHPQU9
6w9RsPmHt6oiTxHmqgXo2WiuklWZH4oEkfT7il5JLsQDPLuJ1Y762j+JjTCExNB6fyd7EJDsNgnx
JSkh8iVQq893FUa3/BR5eL1Brob79tvbmviZj6ZoKF9OXmgA60X+wZRousxGR1bax9MLPHI6sYs/
r4IbE9N50t6TLefr+G+VVT0iJVem08ZiEOeyVTPc/08bOX+U6guxoIpHmMmXmt0VHBkLk51yALcI
DsU4/Mpb249dUQfk2y3CWzPrlaAS05P5TaLoNiy+97X4JztHgqkK1SJLSrQiIFHlGYQ5BJrDwDbB
BqK8DTPkUsSo1nMo8aOUNkoZowg4jnRmfC/TRSQiL9BInOj7XJA3N2eZWaMsEOXIgi5b31SCQGzL
RMgQ3qnbmkf5cFeHYxiULDZBXkVdtTaajJPlvRy15LLCLVgHaUEmXdhG72RTgGV+a2Zy3P47ny/m
BN3tJBdqs1Evo657NpgWyQw3mySKb6U0zMjJ+XWZFZ8LvIVS8zaPTPGAwQw9MutircpZbWa/nyvX
bS8Dm23sKoaXsEZw2IP8UhFbDsqGR08gvnrAOZ+e0J6ZEG7OiDd8muk8ZFm3ONqytyEZDIzzuLeu
RgysvBxj29hxz847t9No+EY3UoL0p9slTIrJeMmtDo2+pHsVMjAE2kJiR286tFrAk7esD1xSzoxs
F+YNKiwHmyebzTEpPa6PMsQZXBfV6oMom5Fsl8XgyFibPnSgZo3xAZzTPiZYo55MV30C7e8QuVk4
VAKS9fqPmc/bcRrRflQmlvlettbJrhGloKSsVLcJnh6I8noQOmgckuXoZ4aeT3ebwldE2ZsUTBaV
EAnpIaV46j8m31MEagerwjxVGqgscfnNR0jkUxwFpbPkC4QOEEbWPnwFLs+YOGW6Z8yLkdldYJUV
4fJz3C4TeC6Eiw0ocOsjbKz2qyjhxpgu2SE9lj1/S9aUJAi0z44sRIULmqKsdI67wYQrRD1oXmOU
U0bADl33TdLwQJ1Y5u2itxOrDYvqLfeWbRe8RmIAxkxzGrgOeNzgOPiLbSl6gPII0KVdhwc+kaOH
oF4PQmZxdGzjBYv00TCyKI4xIiicNogsvnWvPFQPlhxOtS3ClhOrg4padFYK/UzmxdOkdgnDN4xm
k0t3yhHEocvNzlZpzhbHpmHJd1UgEfXJB4RhWFtQJC1icK04NnnGUG2J6GU+0zSNwzqzuzMuvQ+T
8JaCnwNfxKJIZZqNUeC4S65MGs39PCiQ2C7fvNkuX4j3Ru5pk6Lx+tyXsES0CouIuuOi9Xeb6FwP
nqySnz36QJzFfaWhijBP4+UELtLgl8Q9rcUS5jCVO6gRkPbOmqreVnu4Tms2F8sNZT9couhT76O8
xrD3HmgWPUKFDVGcftQlTDAPgrxiGQZe5BqS9OQotPE936+cvwF7BaZwkOpkeu1J8ZEtRaBhqzIt
Y5SVCDinycbV7UdgyXduXZ6hMJDf9Ls0Ui3MCk+XRLy5qKO6nmwOopPFKRx2GCrqJ6R/WS8Fqhgy
Brj+I/V3SoLg7MdSi01UoKFxGFpUwG23AZGue7Oy1lvcD0kur7gy9xA5DqjaqW2XLNNbV9j62+o9
hE8tKQ8+RoWmJCw1eORhO+/G+yZREES/QoUWfwjJCeRgUgRAmKmhBAlfonk02c2LSVvto1MB2aIG
WyJmYm3vtOYeMbp/Ci8v8aPWh1kCFOeP0FCgXUQLy5eZolgWdkruMy6g2TKz63vgwUxb1eLeitcR
KclFOzwfvECtp/Qir7Ok3wB49UFUAFhE3U0NHAOdGFKb1anLgu7s49dhvgk92Q10m1hXqNQaQbxR
AyqGc3bTTFAkUL3gJOr6Dlh6vZB8+/B6GfZicXEbRVIiDYR8S2tJQDTUuBUkpAz7cGQXwo5IfwBF
iSdGrdRl5rFl3dLR5bjkn/AyeXRYChP7STmL3RQqJ/BsE8dCTqsCCWV5U4TI2/Qz1XnFao2FZLy4
G//4jBytqe4RJx9upE/mllmFq3DecBHTlfg3kuVNnSedoar6KQDqgrSmGr/EsJdQ/40A7t7VHIBt
436pa3KLbbTZvHL34XxRkAHaoO0nDKvcYvba0/eAAQjbCoaTNI4QJCPJsXrcqbvmz6NPy4hkj6ze
4WgH/MpEn0wBUSg5sjqo/T4GRH6B0OF0uCd5+Py0K2kd44iuFtAOBIxj4pHoS3u69SNFTP60QYqv
h77/RmH5dDp+f4x4N8YcdAFI/J+Ng4VZVBmvXDzPZ6zTSVaTKOaEhTKjh+/w3weAXmlMEw24jSTX
2vwePLCP6HYRD0is0sobAEpJeSS+3b1kNjBLWTOV7ZDr86FX3KLZevXNUmef9jk4Pit55NxPevSU
HlHFZFYvEBshIMvBZAt1Xu/dfFFlQnjlWheDrcsWY7CIOX8IrvNxrXxkCyhp7pqM8FS7nxIbqZ4t
5PT0y1G5kXhaV7uwzFI4g+1S0ytgtfmXH9CXYSCXg116hirCSxjPDI7iFqc2Gs32ZWErWIdJ8cGA
PK37sOqE4x0j3ZDsUIQvmUminJE5lBMKhu5ji6OpUD7CvQSE8vuanLyUBY1LIKfvF/S9a41y6FkG
WzCJ7y/JnkIsAEODdQef37Zf4WMqRjuyyrdeUiOzZyz7KrW99HETg4xa6qW5EHoIgPNShSi39e7f
etKmwQFacbVlWaYzSeUM4ZdIR3oB6PsHRXExZAORxYn+4cuGCpj1oKRHumf3mcUoeveh74EpBRkQ
2KTrmjZdYDJrgeXDY+w74Ve57H1pLgpGFTQO6B3AOsGR6uv80L+5Its2IeqH3W4QlknA/4zd0a+K
XrsqdQlfhJLsNvPSOFM87zfUzyysVZmKCOWrP43s5+KgJjTSvj3TihHs3uSEp7l5HJ8EWye+3dP2
3EbcPlfQFf1htnE0CkIQDOlHUY59n0790TS5JzGJWEBM/x5jzXQ4497fnYK3+N9o1uLNKdwATsFy
rUskmF6Ba0owrXm6XjkxngWb53CsrvL8A9mUhrjOs/wt1ChP2XppoW8c9QgOvOp/qV+6FHxHzj62
oesfj+ZHk1U73nr3i+q9ms+jgsJoarmLYiXEpzciYtkbz7NbXpb6PxUrvys8vBND+l0UA9c5UyIE
QeYrgCsyfghQN/pliaUSgpu/E9yMjjZ0wcttsjAwQAoKOlGfJvVoq4oqOMYyJT7FU3EnV6jtBdDh
9s88dSS1yreg7ZkDajiQeFK5phy82I2w6yxMlGo9kZh+SLUTtG6menR8hciDZBqgWbacjR9hR5v4
ZNfzljK/qgFCPNVblStS4UhyNloqpXngaGsTkYm/VoAmJ+sceoY5nUFTfQeS8n2urjwzJdI+uju6
q/UUxmjacHa4ZXSC3HkTV8CcF6ypKabKEsRzdYnQ+L9i4cDxQZscXSvkvGiSucmQzdTtqYJ7vzxo
pngp7gluoijNEik/xDiO9zUhsnte4bka8xE4Bwsrxm5KnYwAuSUjiAtIMfgfqUgoaJL2kz9q1wFg
CIgYzseJoX/gqfagkZesNefBgVfaoPnzZe4tq+qY7uCE/uC07TG/oUVtLC3ACFW/Eiz6jgiwj2d3
T4gjazV1ckVZdAxpra4/sp+jv+eEmX8aEj6zYorinUwqdhqdwl2/e/MNidGVzEEBZViAjBHlcVkN
fIwvAKC6tKSox5yzrB+01I9ey7X1TuhKaXMKh8mUdg+HOQk+kQz1OqPP5u7cflzrv1wQDJtSnPd0
OSCLx4l/AivW8W+mB9GGExrTQj+MHzjLSrit1iAM467Fs0K0hfDcu/aAQ4az9pZqycOPENq85ueL
myRWkTmd9KynfLGYFzGUf+lz+8Mp+LYUWNB0Y6Ai5yOBwXWAVz+3e3iQ2+Fae5OmwpLjhQR6C0rY
IhPXQlAA56Y2UHekwyo2zWdGsi5ePTgeADFOZSpKP4KlXGjPo6LYZIUEm7u+UsoZdn73LdyKEQya
EeEEGSusmQD+hJ9td/ETubhQiOWSoigc59w5MWGSZGiyZAS8ywxno43FdglXTVSiAkcHnlwaNihA
xXqQAu+53RPxzHPXrFyL7YNfATYp8FBxvy+ll47Ayj/+LlU3RFk5XvQQOqYUz924eNN/Lyj8mVdy
BLqg9TvEqPf+dBsn6gtTFK0H6VguB0m4ILRawjtRgzdr5+96kOAfODESNs+UPSSquVhlqmN5Q+Z6
qEHS6q3oP6IUhZdTcopRUeIn+nn5JOdVXyAzPGTDo5TUZw3j0nByex6A6039mznKFyU8rsNx+ha8
RoIAERbh7qfEyy07AeZpma0374s4+mvWM2ZTRgIp8YWeIZZ7NuDVlhK/To0oDXfdtOBqyMx5/vsH
slw2KXZU4CjNv7Fy+qQ101EYiB7HUyfGB8xXQTz+l2RAPwi80kNB1kvzmv6W7t1BxiCX1bdAQJW7
s3PzogxaH1rWk8xFmzOjJkdwdpntqbB+AthaUUglwaxnF+B/B6roA15PGTnic5f9QE2CdETrOByh
PcdGMoWV4eDo36ry1EwZKsU8RaUwfi0jkmgrBvZRTiTxzzGd+KY7Xz9A1Hejd3UWoYYgQa0Xm+Jm
6NqjlJo7/n8Xilx6528/gj2DQ9Sml6ay1DNM98AByaDhTjvuP8aTLbcV+rvYD8gcjrqTj705pcmP
6npBqax7CaAZBY96RHV6yoOPzOfSywefZN6pA3JpjK0Nf/rZR3S9QW0UOi7qHbTQcIlKkT5OBJwW
XC6uvCav/bTha6V1dzCQAFVpPh+/YmYt3KhwQN2tDIoVawuc5AP9/hHwE7DMU7A371klXZfFajtt
B2HFG+l1NyKvUzTdBzEKvGRzfjgBWAsvQHmMzBafVrdOL+4gCy4p1OvHRIFvuwH+a5CarcFSrIox
FcCwQNaBIbjVJKBeUvv6/sg3W4QwvhLXbd0Dn5tp1pv2YABq/Z5krBt/SCHnc0wyTa/KLwDkg+Uz
MnumjIcwa+ZXoNgrP/GyBBl8CiGiGKYvj/KLFwbaHzzFFsgkmo8Sg9OqJ1KS3KAMOtfVJZ2FKhbb
Vs8+Ec/SHSS2xaOmiDAZNI0u+vV36ZBu6hURWdVdHcW6yE4A/PuzS61KXgA0uQdeVq/otZd4jmhR
uoiWJOFsnEX4dNoRUeg7KEW8vnRUsG3ZVASST7O3/HG1ybg3D2FC05fPtyDkOctWAxAMhYC1HHsf
S2mvUeMWXAJEsWHFnPInDCzuYceD+edreCX1nvnZ5a0OJ63vMJ3BwwqvwbVsw/hVnX5Zjw6iZcC9
zkbXlI5qL+kdsbIvj7IYHHHHk+JWav7RdabQYvodysDEqXQCnjHbfFr2+TtKVu5OR20c86HU6AYT
n5XH/ZIls1d8ET61y1jFwLX6ZelInwSHrsmB4pLM/0ep+FdS84ab66Mu8OSoh9LhBwlTvlq4qvJz
KHWXxgE0ilzA+Bw2GjcS74VR7igDfyIzVdIzh2MWVQ6/9VMakvV38345/4kz2kCpscA34IbejZuy
HNxjYTNRd7NwDuYZLUjhkIIjCCBhZK2gMMRWVWGTUYAMaEFL0nUQATj7LdbcYYtJiSIp0KHfADwX
83ms++1SakPBTiCFFSb7ZxCja2t62SkBghRfVzKxrW12laKn8n/HS2hnZgxjVXiftdK8b+LFr65h
8ypg5+M0Tp0kF2AARlMgeGpmBgzk2v9QaiqxOV1JuoDlurc3MkNLfcF+8nBSEozWWJJ15SAintjN
CLgyR4zYxL3tyPOdnu+9LgSVsJLo9039VAb2CJpc3wlpMXNzpXYBxmLSgLN62QPiwEq9nSVkghFX
4AnjS0jHxSenaJNbctn+Yh+JlrUxYHwPzZ6OzQjn/j7n02rMdpaqsCBNQGc/OXfQ3bWpFgkMiBwf
QXmT1GcLtN22XJCXsbclEuw9AcQkH56RYs3MYr+hOhX2+NA3qEobtrhnr20Z3OiDZNE19UFu3Uve
9Lt7fms2QChGvHHhmLl8x73WKXcsyROPwXYP6cKcyhctCClCQXhtOT+lfr73fc/ezmXx500xQQHk
by3zuqtYb+0cvksYgnch2lmBctayoqFpzpzyYHWEMMLGLpkUrS7G5fiOZYxiL1smpbIuBdgIY9kB
9KXY3ImNmz+KQpZ9Vcp0Jq5HLGqZxKgldnM2AtqwhenMBh7JIaJ9+E0hEOR8MSWVHcuOdOB87f0C
ZjgkWBOnTJAAFN2E33oFBIRItKedJUXecY0Yq20pDrpXNmeZC8IZWfjfQoMWQ4zHBZDyWXk1ZwmU
TgPL/IMEy/El8bOdX8RTXOy3qrcoM9bv1CITdoSxRp42s6+MrWTxmU1qJGkpetuhdw/nYk5jInRC
tRtfCwxPWTps7N82pZkffPMzodXEM/39czppUfkmFfTP5FDgak9Fz1/KV6owmZQfAfK0M2eDHHnY
0Rml4v5HF+uI254hH9zeoWv+tVPQYbBXu9yudGHx875Aql3ecPdkRct+7wYhsSRy7Uph9SSvHDKx
bXpzuYtkobpSt2M1VE3PfsntQI+7LRyqBq3K3J1/MxL6OzVmNiHoLXEZHPGz0VNNyu/BemC7XxCa
H0M2KZ0AAQE4kHw9lgAnXRO8iJ+WIXU0MtfKtJLrTijtnpXceKvOi8tn40YVG5DLNrRsGIbk7HHS
pKKHllmHP785c4+Zn2i9/JbDWi3VIBKy0JqxJ2oR4/O8YR/minW3qAR4qC0tJgedmPscchnb7whG
K++GSMPqMxUJuetF5oifqCDyb7fanukTsDqtR7YCgV6ghHzT5ihG275L7OdmTQDfdDOcOIuDApwO
OGpxmL9anaXxrENigme0/teLF22zQGKs9HYFw4xvp9u8iBwY/VdSynV/P813eIG2cgRsu2h8KTUE
Ojp9xkVfpEfajf+9K7Nx2x+1OmWZQoQCG+8Cg2/ntJFzO8tnZtTXMs8Dh8tbo4aINpL4j+g4OmJX
/NhILtJ8ayC+tYPReRKueuJsFEwkt02R+38aQAxzogeu6AkinZUKYqLpfzgO/HU5pA9rXfeHp06C
e6dpo5DNL+6UWjjyd5TPMaXDxAJnk+p23MKBYB5eH5ME/ZuR6k942o01RG+0C61rb75vmeoILTI+
9uK1XEkYWRrQNYbOC8mjXkspVMChc/pJamWJAxrm9FHTvVpHNjdq170+hLXHi2oPAXhuXtrJx3qd
BO3UN+Gf1OGAHWzY9lDmcypANjbrpwBDyYAcX4P6CoeQBnV4CEP/Np4VJX2wRaGL046bLMfJNY0e
F+e4MmcQMtEDQ/5nn2vXlR5pduW9KTEo5gds3vqRUJnhux7dLwt9LsFtpFT+HPIB7uTKGm2OOY63
LSDfKMoVPgLi51D3S4H05fSMYxbN54b48RpmYmUxcZ/VA5Ho1V2ijXjojz4F38RHPnmX6V+w4CSM
tdGRxJWlr6LRAYX64cOIDAoDjFzCX62lPyy+hvFvu4FXtD6Rfj1QOEydcayFi2T4K9Jwp2Zsr1FW
uELW81dPiAZqu0qDeLQt36GO9YBCwvaDnnNS2l6ny/slZ8bTSjSnwpBrJIFr1N6ZsJzBkTB5mLsv
cTtGlNRDbZl891GHPcIhz7iGThJEQscejUvPV88YRNzE4lj5OFK+VFn5Q/mS7eeoxISf3008K4M5
BjYR8LaM8MSBFBO+HV/wr0uWNKXvdo2rM9DEPnN/XNJKYcurU4qvL0KkymK4IV4/RZ0XxXbroshl
IM1wwfavx+Cz4rr0iA3S3ueeRzcHmszvUDHYNxUHwOf5yV/OKMneX4RVKGIFPf9EDl2Kgihx5qKw
P+zfNH3tbH0pLyJUuyTg+yAS2RZ8B6ZF2Lnvb6nZBEpIsLnr5Kw4gCagbnqRJkTt2/wRkHqcX6hx
WLnypab/zNGRSamiBswG3g+2u29dYyyltUrR4sA9yv4BYw6Cq/5a+lXXZ+gtqvO9+WlfopL2mKme
tdh/NBAP6frSecqTFeRNH6knDruWn34JPNgP+RLdVzU7IDsTRLxUYLgvFV53vJUfMHcoF/V7QONA
8B0+YoSBYYq7h907fgzV3w2+dZP0s7wvlkavN+Zl3tiyqqTpbaKLj1yPkyEEWIGl0reYQdJtvYHO
I5KpAKNu5CK80maQSpZOjchGUcjdNSmee8zZtDipIMFGvGv8niaQXLBDi7nzMBUJh4ni2IKxGv7l
vV2udYFTyFnWFXf4OHLc7HH2hT/TdBx1CYeLm10bzG+JVJFQAVg1YbgRbLh+RgJGnJLUr6nzzUVs
8WPmfOqVlf6mfIgAXXhoRSwXceXgiBlmxnLzkW6gCzcxQFKJ0JM1m4/aS441M9l6Mz2UIn/eWL9V
5AJnsWQmJ/fZgcodkEZftfVwGuLT1hbfQcdTAYg+L0k1QPCJ3MZ5S0AbD/Q4jpoVRlM3znRg73Qh
oysQYR+LK/1pouIZVnhzXNzJEtdK1/hvQsIdzmn+BRBevLPAfddYmK0VqiYE2q5EMObfT+1daD8K
wrpgTpnMASgGbIjvPHTOcMUgN8MDNQJYKACQKkpBbVCeMP9OMmhxyTdyrxOrO4gJ6JII+adc07CK
Mr6ThdWrkRu+pBgZQRDeZNXYvby+cebUXmteDg8df3YG/l2yvjwQjgwCZphgI6sflh2biWGrqI1l
kd2EYu7jHOgAPMkMR0zAaFZAP656BEU2PYltfcvJB5QDJLjJgP5ES5SrKwKAo7LWnniJx2NCr0rM
YqbRWATKBD8TGcuADwae5q7WpJXV/ljURa2vavnxteRDIDpnbGyzLIaYyEMW+egGIjPobfc+h4Nx
4KsipAJpe+YDLwjQgc5MzJlpRrX3XwVumrVcTUVJwpHyPCNqvseXozdOXwvi4puYNj8OLskVygOy
H377/MmJ+a1pGCYuudkd7NsG5nGsS9YZX/9p6M1ImRfp8BlalxyJm/2ZlEEoTEBSr1x9E/YYMAjn
KIVi7v4ClQHqEiwVZWQ5JiEk/h8F4f7HximEnWspx3vUCABh+1tNuYUqn65kxqjRVOoqEg3WGAOc
s8boFU87qjJMZf0uwwF/MZICQKrr1blBTl/lmMuyWwsYxveRaZ73VIdoZfgEKjNK1vMiQS8AP2Us
enuexoNSdPhDAgy+HA5/8l0Fqa5vaNckTxRy51LOWGpo/BnH0s0Kj43kIKuOmjtmmI9huP4GDdlx
FXOfWT7t90GQkZNkENNzKHqTEvTIw/JhPI760UCPq7YOQat5g4DZ86oizxJ/yjCDe0E3kyS5qH7Y
ERbgxCzKv87S0LPk185Ij0iblHvSPpyXTz+KSA9CTwX++ceTIU0EEUmcljGMd6BGYPoJ6NiXaxo8
3gbsBLr+uIGWSGHwWH7BG7lMVaRV04a/vrew0INc7Z6Qx83KIy6vTDBMdbk36MLR2oaFbKTFbFG1
XyMEr4LP3QJ0s0L2WR+lif+Mb9oGdlcNa1/jWVEwNWLEcfKJSapfGKC/3bltmgafpqtZR65E6+qu
Nz3iwrx49JCKB/JMcHjqhNUYwsj6+5KigZklH+dICTpYVoAHknud7iCeEfBksXUGEW5q9s8gaL02
8DrhI200pbLhoMKO6yOUdW06aQSvPiLHTVRI1R9ugyBj3CIKyAK9UsGOFtUHgXetfweDppArmsft
pxfH4I6La77PkKQYEC7Uf9H+oITgvFMc/LvSK1tJxgu41K5xzgedSaHKLjO11RYrRWeUqhr7vSct
DuWeb9iQl4SyxJb68YR6AO7wE2Ws0tHOZBb8vW7zAynI5f7vNPyU8vJdokBk/kGwBrdtM1GH5+Oe
LKYttNx7lO4mYtKEds4GBM1Idvuf7O3bhugoga6zCwlnqmbChVlAyZL0R1k52DEwu/6wxbZE8X2d
KnvufOqOM7zeGCiYMN4QZ/iQ1BvG/4THQn3e0/s33yvs5HFyR0pE4CpD9qfj4duXavCykK61nkJf
aXYTl6juSQq1dCmqHSfd/a/8bbiDnnysnop/RJmGqL4Swnv3+SJfQzOBq/SE0EPdut40Gk9esue5
NUPd8X7qmgrMlNHwSEKsknv6MtHyLzxCVBE5tk+g8QVMSBJzo7NGBNEeNpIGA3oqavhTbb/woVqk
JKh5nVCdFK/7JRNm0fWsqZJatpyWgLs/QhdStvtDn9FGgR71VtothBHiyxtsf3Eq1KZ5KVG36BU9
m8Cm9DUsdx733/wTPNJF11JaKFZz2FwLmpYBzNh310+1BK/KsRWqkSI/UkxzKdYzIW0BGkHgsTw0
0Nr/q0aNUaDLSzbP/kt/N4DC0uarYDPTGAVccCKTgeWDb0ZAzOV67aiGTV5dK9kgILdhG6eFk+E8
7tGC8HFA+pJhVfntmYNSZBnaqmQGCR0QpLSimyqpAMjp2WrQF3c6Pcy50N1Djm61E9qcY4tSrzZs
KytE4j/LOPZQ+oi9i5kdsV97HLqgHPnx5jdpisYteSVetyxKDclc+R/NM+loxQSxn8Ptrkt6jJ2B
iAzbWYZvaHggqKvDR515rEm2MdbwryCrmmWUMlzxDQ7M9sTLg/88mzw7zEWd6E+xr3uv698Zfx/P
SuSnthVGIpvYtbeoAmogmdtH54vDexh2k+SbwRfToo5DX8TC9oyyn+eeTr+/EKbfD/VzSvc9mmWy
Lr03Widx0O/b5bG9I4vvoqfU0B10VKob7GvQ4cfqlka7+MybSL/5m4UFBQi3BE5fvKma0kiCdoYO
zkv3m+Sn4yMHzCjUE7ryFjS2FggZb7U+rgbGKU4m0l0GeAn7U3yoU0JvPku/etfXwV4YHCFQt0Bb
i/WKGfXl+eLdNz3dL8DlJKrk+tTkHI8DTpeVezyN0c4Zvq7/My3gAA4HgKN6pdK6PzMGwJhKYrLD
PJDyFVgtE18rA9K7/+g2gMlIYhO2Y8+8XDMEXh0V9md/7sdDCNVtlUO5lFaAW1auIumzZCbXIlZt
zimBDyE6MohIEJyONva06yQ//MYrIduyH+KHeCm1l9PnD96LkYd68mgK1vN1CSiovBgLaMyJmNRW
418IB2C4Fdy2Izl0PZeK2FZV9Uf89tGJD8RQBsoCZ6ACvi1FzyYGq7Zlw2Juq15T7nmDS1Cb+Epd
bDWKc0FALW+t9UKCRTnsMu6OQ6JoASeG6oVYNsh+LG3tajC+o8tGr+PABMCZ13jGr7iEdWCcnv08
y2cqIFh4Dmqr/I7D9E9s5J8L+qMQ8fBjVLb2kwqPkVuh5gg/jWTIpgYlS3th1Ddywylbw6S346TI
ImVoI+Vsk8xQpf9e0W9br5T4hIO/r2cyWaK3pbajtzmdGgcmak4zVtzYVOAiee0YfICrSbpM4oW0
ET8JDGWFDs93PckCx899vauj+yP4gmpSCTl+dd0VOiWjcwpL7p0pHmuyeGCLrshD2U1+VFE8zT1E
DPfL449HjBaZD2aXk7v+zvJgITozHgAeti7EjCxN3rSUT6pMsF72hpjJvETuxJAfcxqlnNr+ds5p
c2GG4R+IkzPeL5R2fEZ3ZqCLh/rFAUcfCKmMTOYYSdBEps9xscFzudPqA2+odROnJLh41jhzwlld
3P5rD6i+KpBvY3WJywsX0blzh8Hln3XIQSbx6iClkxqf2v58a53119ijwU6kZy+WCHpr1MeKKDU+
MOTtc53goZqJItQplOqqR6zhKTXQPccbXEPJKvjIJEe95qcdZZ1oeIEHnRlh2IeGU7a0sy5cAtaK
b525TN48eVfVdSbbuPGbSjyVqrAJ7MO+yxsXUUgeSWWTDqJxekfHyk2Ji99Uw364vLp61amzmxgL
ohVW5uwGNYSzJTmsNjcSyepfQoEHKPwh7Y4+RArVpJTSfat3zv9DeToEz98WLufKSmc4LyWpS1Ky
xkzdrK2p84T4ZbRYB3Lm7+uvKcFIrjuEz74gALViZuAEJiLg4MpsAMp8YkogWaNI9qdrnw+e6XJB
v4R/suPlX8xSQHpwumFavYRA/IjmLDa530edLogu1ey9/KwW/zXf0l9zT5UQ2ti1E809g/lwgMzs
1lYFi1jkHnfUYrvOAEyh3GVC7m5OLyAHhJZjTgcFue4yTEaM41Iy8ULhk9Su8/0XnIMdsj+xzE98
GADrqKzZscQ4mcOvJ1WFNzyxSq8e4vFr7AfRKOtS0IE8qWglPQ5aXCSr579G4k8p+clYowLLXKbx
6Yq3fKmfnPPOJkZ6YZAWrWMYF32nwlnzTg8HOup4fbLTf0g8NH6fxXMWYwroxGl8emNluDAk5ziO
AG3kqSZJps9VqmEyQ/HA1eS9A6bjQTIRRBdCFdJD8uNfUn5W+eR+CtGZNG+LqPXdbY0svlixt0nw
m9FNf214aysPpNRy6NxBcTYMf8Bmew9GDFeamo1CX0KA3roLqWq5FusUFoKzjj6iXq5ebfFRHRiM
LTm2GaM1UrHJCB9H5BfsyEzmFGgCUrtIPdkQa0lkWvo/TVz5e+LPjWCfDC5i5NUPGteoHmluR+in
3TLkKeaICN0kVsrlktFASl3yqOHr3Ga2fb9gh1dIwIxTH20OMAL5gaSwz8sQt8d9YFL4wacKBpPH
ls936W9jC9XO0AKmMkdbGavOhYP+sq/yPJdShXvzh4MJA+jGedZ28Gin7ipahLhzGwR297mPytO3
vRcLBpZ4hjtPOwQlwXhTYcTchXbt3WVyH8R0ngH0qHngUsk4Nrcs8Lkk/xJ3QpVHM96vflhJ5fsP
AkocC8RXSL1TscS0dLj4g9PJiP1d9gM2R4/S703a+CHHau0Wybo3Tl5BwnvM3sjWjKBmv+qaLo4F
tKNk5JdFd1sRPeOnBoOoZt/CPjlplJkiG7VsR7I6DCnS3DhJnDOxJtyCiOdrUzi5YdFGc3pVZK/R
yEbEvBXB30pCachhjTIiPRBM6mnyovssdeEZiySf9BfG9Btk64nS0+IeM2SVzLRXiu9Xwt0t5Sr0
urTNBMoH0SCHxrbMJCwR7RY7BlKLQgGlo+x9PrW7V/Cdr4TBH3h0OF6+GR/+DpwB92rTrM9FOR6S
J0U+u0o+/HfIvv0kYyglykJiCYWfVW0XfycbzfNHZlmLu7zpAifHPYo9VPRzTlAixY7TpvRk8tiN
z12iQARISNVSH8PVQWiayEYEkurCZOCcPzwgk63sYea8Vf8IkMN4/9JzNSwUpDDLpgYXIPLV1KMF
QsFBmPg7JygIWsOR//S909c9WNlw9usEDPwWCMw4rvBsw+eF8AulPcdKTRg4MKY3IeVf2+utR+cH
mCaTZTSgK3pHXxlHpJQQ8ypAvYiNh2XrnDW9wyQhMbWkBaAPFu6iEiwjjX/VPv+Vbpn7qBgxmpi0
BHH78GwBWeTZzbEAZfjoZxcmC9y4qvghKSgqSp9+oZY+Hp8aUQ0iFfvnOANxFaqg2hiuMXrm0ZkL
JlfpBZ6JVe8yRq2jPu7574jLYFYxhZqPNPhaJgc5gncNFq5PeAL4JBxEcug3kC1RFoMFgfNjn4o/
vL3pUrFTt46i0cAV7D04JDPFpRGRrGUsJTOk/SEumynQSe/iASbqoVyyD6llys4iQppzeDNWxzAD
mw2P5edcPhG/+qA++atkQdMxhRMPGqqPt5dbCSBia+/toDSiFi+OEypGiUwpO8N5PePtnhLolQ8M
PM3BR0fCqC/PTWx+jgqp73QGvKxrX7mV63v2NXhk6AwVcHOLOVmaDJY+q+1tntt4oDjIWMV0SRjE
Q2A43kdan77PoSeg9dQ13BNagTKkeNxhfzvSY9xmB2teKt72t8dUCkWJVSpc5e2jY3VzY5T6rk5s
h3y8KaGvEM3MOCHMOZ9olaN5U+KSVb4wT5axYERq3+Y8rvr1RvN+8SgYmIcc1pEtxsoSDvwaReMW
DcADkL5rbp4mtwYdoJ7VtoLjSM2nGxE0P34CBQXDSp0U74H0RLVzqjU4JKGEvZW4rwvOYtvdqEYD
3C3fM0BXTLdI1uTKPKWtKZ23zegu5hgj7wA6sj+zjLiceWAcj1/FQbP72LWT53hGGbrjqfvGxDzm
ZYD7PduIIkFOH3ryrS1o2waAkOS2bvy9nkhk73ZuVsxRjqEmgY+TKJspZfg2DbBfZaheJQD+/Xff
9YM/7AhM4yT97Lvv8ACAvDubSUeiF4u550cPd8e/rcCdlvSdkKnp02ktVtALMpsNxJGjbkd7ak2C
VDNWY7TE/a/2XCkFoAq9JqM5oNuGLBs4PCxLftCxFXEK6kwBS2pMSEsmU6yftz8/HYP++kdG0vTA
abK4Wz3dzoX0P6K6XWvOjg7yapzp6RKtWk3+0Z60FJ/12ukYVphdYIBtTFmplmbPPSyPIDyS8mpP
Sap5Jku8LWr5tpTbmFFcFbDl0gBVMawFa5y8PEEIzVfNP1yn8CWEL6KKA4uCRaNRqJtb6wrR0ii1
NN+dnt06Q+D15lFJOGr7QdRKxHpm37acLM/yAm34CJgGQLz0wWFX3xq6YXsZzn8kV3GjTWA5JRGy
3eO6AdmRb46DGgkSkkcRjNMalop/y+2v2dQIWMZABBdIM6DKDbWljJwEP0xMnb8+P+d9DLtsGRlr
J44kHvsulkiT68ta3upAARp60fpBtLdqBUnfJtiTg9r3DU2z0Xl5CU3PDfW19PPxwW8+0VS72zGz
Tv+p76ZjBpl/VzyA2lSmFGKUyT/SqXy4Wkn9KavXU0BpSgRUZ0kVcotZn+TkiRTaUp8MXn/lLo3n
j/OVWU7Hk+Aih2TnPCDiw33TjNmryhtWAuZt9u/1fdOR9oOmfke+y2NN5SsrbNjpgwfa3xRZM5Qh
LLHwiFoNalQWJxv5qB6fRnTZht+cdSMmTe/VT19H7+J0nVZ33uIuSz1/nq00kTWH6GuAkYEyJCXd
xFBtIPCvMy+54OuYBGVjpZvr7G7LXmbfx1WURn6vA7E5nUGFJKuHpdT9FjuM1nYzlvMQ0Y5qalu4
OXDjwUsZ1AsR+msaSSrYwTdXPWhQb2JKZVQxtBSxvcM1rzNK0n5MvW8gc4BicsuciplY7m49l1DQ
SSXJCsUWpvbZM8LacuAehdWy2CBQh7HcV8QdbS2RMh3b30spZ8XfBoMGvbmguB1dl/uZdGwjcEf9
ecRkU6oC75t+LGskZ7En1hAWrRww+k27ay440KWT8JWEecjEFOGpDXT8BtZz8j4uKNQZWCiF4jJQ
diV1xmpPR+lO0Usod9DPmHhk03TW2apomvFU7VnrDXR8jA2uQ3G3gbDztG6LePeE4H5wpy65ZTem
y/jXwFpMUOBvY2Y2LeVVIOFMvstRIhWdSwNxrAHfMxycmpZnzher1FKf+1Tlat6gu0k32pZfXLmk
upXd7I2jtNtP4F35x4zuS82wd4OY836QczbF6ltOo9mpuWAAq+0U/LJ1T5+XMdyQiMpn/MFIMDxB
sDXIOxXBGjeTc2sYPYRDeu/6l4qMGv4ab39B3/SWnUdbvzlcBeRAIT7VCa07zHGc8liblTnIgAel
fYEO76lf2bB14z0OFPAPGyBzMWB4ZuqRx04HM/wXqDXv8WrM/9vzVXxsGqsdNOI12gG4UhWFoSy9
+3NoSxIAKm36lPSytetblDoYygA3ecHUjX8DmAFxpLcvBsQFq1zl8YW947oktiXE9K7+ZcmdhfXE
U03MNBG8g+Se1vfyW4GySLKHWUkHUGuj3WQBxufuMVZyRv7efoVdRBXcsy0SIl6Zu36qjpalD3q0
AnDJcugXe6ySYWaO0btuffzIDIYwMu459iAsHcQ1WSOmNjNYJRU19OqhPWVOJpB8d4sgo71vh2x0
GRyNEoUE7/1OlUK9jRAJqoN3qZYryMklc3WVuD2T3UM+2G3LxS8m0mM5V/sM5BUMIxOSPtJcow22
CD4f+/wDHMaGaZ2vR9ujIxt3Ozy0dZ1rTSPKB3CbRGItz6qc1zKNatNuRA8LY8QfwvTn8g5P2nIU
2Jtf2ARn8ypioP5t3UDor0cENCq4GhfEr9uRUTkWwwMFVqIjruECeuo2GiEjQ8sljoJ5zATJECTa
zVV0lrdT6KkD/bs8Qc1UP3lok6xoa6RrGK4cBKerOy5XZOV180SAE+hfPmLc26dseRfUbA5fGCZh
0xRZsEmDJZ/Y4R9Vm/MucWTs9uWzvpEaNUcBJGB6f82Fw7hOwyG2uak7bqrD7sFDxq/4eWO7AtO7
fgqtDRjyyQa1qZMwjBPyzys+NSdFSBvj9NM7SPBqTZFQPa5m6SepG/wYwVNJWpBW1yq74PVa9tm2
Jk4HzDyt4TyKIfvYdOd9kEimFdXk19SiqAuyvbBnxaacy0pMlV/GzakhxWdXr3uNf3KebDjd6nWe
292dAhFd4ilIqS90US7BZE3DwMNLhrZ7RDQaPMQNQ/kFyNx12fWYlogSpe7shaTVQBBZSo2NF01Z
e6GnYnFFGXAIFnMtNOl+V65l3xlW8+ls64ZZq05TjUZ9LSaSCDCaBYAOb7ym0lcP6pWe97Jsnizg
dRgV44pkC06uppV+aQTJzXIeg5xBgoTJQ5XRuf0T9kaZvj/dlkRaSLn499lF3nTuQU+iaB576qqL
a3xFHmaIvBkDjQeAh9uerp/BbYf4p2/89tFp1jU8VSQowdDXeGWBb2J93S4rbRMHL6PcbIjwskru
OwgtHEIKFM3fvWqH4pktC/hKKNnqWarRoLqeX2YFAnaW/P16jWdV64Rpmwtm/91c4lTd4oirpSd+
z3LZ4LmLbZw3KqHm5NnB5VfDcUQj1yw9zYsjnzpSZ9vDWqdDJdLDhxJ07aTxlrQ6MYsXH7qbz38X
+sroMp68mAJknqM4+v6TuOyQFqrK1sVveneYgwM1pjH8MBgOCJ+5xj6h+iFA+OS1uwwKdXJzdouV
B5OOncMfzQin2N7cPZ3eDZgL4rLzciRJJwGyjAh8uKfn991x1PFAef5ouUrt6sisZ8fe4/0Ljjjt
8UTBA414rb7v7KXntXGCEIixk4CG0Wxup9kMNUjjDvk+n5wkZVb7OVsiXpYi6dDMPVDaw1F2YlGx
yuPq2VqC6LUhEyKOY6IlKqne2wTRJXjDa27b7CaSipPk8/ufwt+j831ICPfWlaGAlwT62t4ubs6J
kA/RKKZSsd+2LTAId9Z5C7ijmcwv4hu158+hSoIlmha+5C4ODtRjJ5kUuDSALoiWvlkR/g8pHB9T
cGcpdM9BrPKwyrGhct9SCL7p72UWKVq2nBTFN4xExGaWtdD/bDSm88XuTCD9nmDGYQKcQll6PjcL
Y0oLyjjhRuJHuu/CPueIxQIm7yGHn98jAfw+LwzKtsL3t62QjPfFZUXYOswFbpBqkNTBhd9OsEvb
YoSfpI9LH2PzUdBUz8ktgCNZyTwRBo86IZyctlKvsIHPz0W3Yd2uC03ecVquf2bqCTV0Dz7DA+H4
eOxUTTDL52atUwmubJxFjDXOj1GR2Zdot42A6O9XuONlJMH6mT0Y7CW4V3JiPFZ8FRf5CBhkvuA4
k8oRLp3Lgt+eFOG28tAbYbQQwY68nB3Rn+2DW3oRiuiOi0ZsBhWRPe+4oPQJ8ieXs1uH5WAqv1Sb
IGTy9zO7Zdgjg0etNBfMAislSxsoA7BO69AvFzRX/p+csCbk94tBK9ExvpX4oKRxrDydfPNm4QeG
YlVG09Y/iZXWm6EXsQwmTbZbNfEcwfs5U/iUSzYdK6qiskUhg9fcH+tllv/4gm/di/ZzACjORV0o
AXncG/SrI6QnsxSEypJ8x9af6MbYoJPbIEwxW3jn7h0vNc0a6qcZ5FmOXbAT1KMb51W2Rj7nudPD
xfsuP9rqrfl29MRGzs4ZnRi28L1IRtTX3exuljWKyx2KEfId8zGTXf1aAaK2MUiJct7y2OddeNG8
bYRQxG8bQ3SCLqful+J0V5U/3ULT+E5Vd2jeB9DmdMF/31jF/3qivujyAQNqYpgCfeyR++2IN5TG
idmOs8zc3eHeK6xIuq5KDskEUM2DgpORCVvNWu2bGe6rUWNVamH/5QzS5+y0toKBizJ4kyLQ8ALZ
0uYG4njb5bx46ZUrRB7UzYA7p3uLyegN34lVzUOUq0D7XJS7kw+AqZKRFc+ZEVDIotBstTByH8QM
gs7yaeNaW8yD31vuz1Jmxc4skJfY586Qrg6NSbZttiqv1CsUCp5tVd6Q6o+lxhT2ztS7YpOXzMB3
gexWpvpNU5xTtfQdpdeR/hCbsuv4zgE6xfkf3snIiBbXL0Vk6HI80DoHPSHuC6EV0UPnfFdyIG8D
qX8+McsimEdrB8gNJING5QsjXssJh2aGRLDUkTVsq9OEN+JD+vGk5PGObxLREEg1QKvFJKCoruN8
XlxBlYJU8P2XL2lGmr4KmbKJJB8LvkMqblOprU4YPDX5zGkMfd25rSp4T9pwk5rhxIJgTazs3KPU
N3/cXnxI542fqT7rPYya0UcJ/omh4rtTj20+xCOvHwlAMPeEN5IUJ/HcadXw62vk1/OdMdeD3PVX
2Bf5ws5ulik5OHdU+lJz32FBX0gtTMmaHHESzRWk/swAQ7srIxHn8sWLnF9OF96Hc3C1fub/64Gc
qQ9/JZ+LLvnTtdnzJUBzvVvCCHD5uRBZxR0kqUrT9UW8+MxI6H+h1mREkAE+GQlzu2fOI29IRTcq
qmqh6l0HqsZ7mfdpPme8pElc77BfcaJ/yL7Pq2AMwy3aWstKI1LBO6nWnoNAHX6J5NdsEWlk8cpV
iGf4KDa3dT8FzbynJHfFM6vcbAU5ZqHGKvs3vHFJ95ay1KwUMOMJFfK6yncdod9CUmWhAbLh59wT
T5Pf2zfyeZTHw6rdvGyyYzooWd3hbgXV7dHTHFhpFn0Ht86lOHcLcRcOAm/6Wf2sx/8cRMQ6/Irr
ptacUfKg5Q/YH8zmxl0hrfaUX8tfDjqKI429H+Hl9cLImDsTYJAKde4aDpwlvRcUNzXQvmZ3k1UP
St/LRhwLGwDgucTdBe6KaK6UTdlMXAML4IVq441hrsopbHFDmQLjMhYzrCzD82lAZj9bbBJI8fco
QxaGgv3sE8Bj9k7iRQY/9DGHTfTIGwu2XPoh+KbP5FW8gHvDLOrmFZwYzM7huXtalyQCl+iiAVt2
GvAia+7xHHotqhv7Ouf5Q0AMKf2y4ts4rFP/BrrFpPA49HQm/lxSrzpZGdIZmNp8S0KwbEYuR8nx
6cuRwhLRKjqnVjgENEZyZ74t7Zx7YOHpC/ckVP1Q1QN6xlnBTQgSivALDAJObMmvP2tdYQcf7sTg
LLx28HLw679eguQfZ3ki7xjn8qbXkIQYzIFUjxwnlpXWDsv6N0z2aqDcQq8U1qqG4E22fEbflU6w
HkeZGJedGqpB/aWqYJjkQCMcihGBbagEiEyh20j7yvdcXinsImJ01WezO/JnjRv/jw3FEvt3hhxc
+hj9Eos1s+QB0+Kykl/xVEgQdO+ET13v5leAkGjswIyFQjzkqsUkJ+bbXIyIGeQxTAv9WMfYt3PN
iTAEtsA7xgy/uiCuMAZkKXxXYdw1kVwsGxiEKpL0/LI2wnQtJsX4NcdTmecnzZjFGfZnNClbPCzW
eFc5U19nyfOFVxTpkMa0TGxrInOS48xNCrWNgXU5lE79uDo/YNjDuk7y25KVUAPHdk0e8w0HbFq+
gFyYQK2Pa1AFDNcHQm6xyO3W62yvQ9xG2qOORbeWWTHq6eZRlDhotEzC0ZCRT5QZ2Jm3QySdTHwz
Y5X7futqsFWXJiKXO3TuK9yPqEYNPJqyU9POvYsqH9QcNWkUoezjzUImLXiJ4HJUv6r6Bth7+ZJX
pUI6gaq99xy/BIUpc1ctP8g4Xj1hSokLH67aMQgZI0qBl3fuaqovFR7relJCfbP2j/5HBGVw6M6b
jdB1U/9KySGjPUScnGvJDUe+1KIcrEl6Na5O+ogNLv49d7dLf6Br8RzJnoMVG3vSZ0Z7NPpkoxde
UCB0KbSqkZD/VQCanVRs1xfaTJG7QwrNCgqwSZcbzuHZQQsO7v85IpyNDatGzgXwF5FNmoV2FJp7
ZoS42e2lvChj2ldtU391cytlUcVIbmsvsi4F2PY74ksMwOqssKX/ix4pfVsDLUdO6PH5oe1ngYqC
oqVkFO+QfE5y7GXVP+dE5trQdGG//++1eagK2tkGRRvWev5E9jYpQGBmxSEeLFtGs0bJ88I0Mm+i
O1V39F1f3SVX7CbmXWKvdoolIMv7AMRNPU3rFZh4Vc0azDyOXLZP/L0lNuu4B5eDKHeSoufOzejS
o5Y+J+BciP2xghIxM6PpzQ3cc+0QcJsmi6MffAdIYVA44R0W790OlrpIgG1kwtpJCVrPSXvs6yPt
mZAPUerFlydCQtUXKtmEzQjFDERX7TDFwPERzSAQm3wScF9QTEz/dawuJlle/pd3z2iDTMOPlI7p
19hn71izZp0HTQqfPw3JPJZ/5RxMylX1h1wFi77k+2U+WAiR5a6NE1vfud0gXoY2q/qU2UK4SJPG
a7mATXVbuyRhyfB/VHl9ykhCLKJdpEuwQyDuyi//eUSWFy+vKU/9rHKLe5VZG3GokDKDfiqj67LU
S7rQrOmgkDyIm7kH+QBMPkgbzOfPJns2geb99OTGb3qySd3jwLXnMkpvY1KfeROXoXHHFqiGmRMZ
BaJ7sXypLnciASTTisLBDisfSntNDZoXcmtSpBS8degmszkm4aTQwGHkamLOXzFsmYL51ZO77i4X
AqGGlavByoxEGbuPAqyxBhO37R2oC/MyfviqNKzf6UUzjDRtfqOg9IA8NwLSh5srdoTpWTH+Q8+c
HnRFRBCqxHyeJw+1FCDEKorqky4Oj8IIqAWi4NcrT4BO7BAgo44dUQZzgmJjfzOGDOESeZNyY1MB
XHsGTPj1Lv9ELBFG8+avpL+Nhw3C5W8seEfL5oMCQtwz7jQ8jfaQIm3np7LBO5jum4Ljp1XzVhEy
N7qddzvInut8Ma2nFaqh71VX4arH8NJX4VeZcaLxcPzkfSoaIAG6h9z1ar8x9/4MBtFyQ897rGe6
Lb/NxmmUqw42e9LfmAzRfUgtP5Fzph169bHKECzMmkpR8UnguuYiPBChQyHhuJ+n04fls3mwwORK
V4smibkIMve1ZOJlp69iXtqIR8dx0FnLGbHHRCRgpvLT+/NQ16f7xRhznCfGb010eqshI7E8PKan
RPW8al77NlfUuF3D0L7e8w0aLbPWa6rMsgMcTxtP+zZ5rAHQnXl57j/z8MYKg6uwPOvWGu4UlL8I
wWKqAzBIcrJdJxJ9FyrUI14K+gvR/75Bq1hrGygHQ49X/5lBx/4gpPpxHESY44kw4sTtX/F5Eias
o/IkHoN4COxh6tQ7Hc3s8d03x3/KP06ENQuJTu4CcwcAVlA5IamouiAyG2yVdTkGKJ9JEzSL+Rqq
mLFlDaHf9lf8TnyUvsaKCuzNsrHZC1OUfYEkgHoqrCBw2VUAmHusCN8jxDxdvudAZ9rcMhFD01/M
s2M7mCYHZDuFdUUYq46oth+c6GFRSnOy/K1me3ahjzq/Cr57aR9xoYvBYv+dYdwJbpP9TtXzLrLH
yEr3UuEnAw0dmD2tqnMHPoMYJ7OBZjH15g/wLwzc2X5CIV72t3P8etM1YuXJCTPRI07IWzTuPydx
9r5NHMI8hgdnbzZo4NaDlIG5zcS/jnQXjNUI57VVYW/Ogo4sQQvDVxLdzt7eOFDNuzg59WuqLiHl
jAlECTxM8NoWjquH9isrGZauxGyNU9mETR7XHfa+6AZ2h+ARnUI+RyuM220WDF+/gRUjzWQIMSC6
icO2eK4mbsTVI98bE2g0iOLsGTcPzxO/aBqqM2lcGCCs0Pv1xm2wn3FryxP7dApBo2dr+RFBVe/8
JDCRojqBrG0aSXkzeNyPbAkDL0ZvN4auypN+04GawpeH2BtllQGbLCJM4e+l7pNjKRhGOAWd3zuo
7s36ZwcG0ph6u740NJ4OuWx554hjHDX+Xhk2JXS6TnLp0DEU3v4gccXya4Nio0qXX5Qz1UNOu94E
JK7b3PApaq3sQ20VBFhgwB9Mkq6/7ufpSZJcuYAv+4LHdVLqajkJaU6VApoOUNu3SEdd6U7sGV5s
K1nY6etIkxy45U0kmUtq7C+LQ9yMsXwHXNovTnFvpSremszEbAvwp33incaV7C5zddybTj7IjUbq
utOR282XdLBpA9bGXXtltYqZVwP7T5qkuviHAXbNhHa2Mi1R/JpaLGWubvaPxSl9VkudM3nTqWdK
dLCfkRHRzad2EngzzdT9HS9kN9a9xQiRqIStd5i+oXtK6RjWULT4/SCogWjlmW7mGVi+mz6VL15S
rzcu3cMBsYpFVp9m3BChSjd14cucsPduZs4GzCtyYIcXhc60lPNBzZlIrXTMEX5iqi4u5jni2uKc
mB6pFWrgwGfvf5xw7vy46+pXluPCPUOOHsG1ZvYeFWoN8Dp6CcQyBXZ/YNj34auY+j+WKGXrR2un
pWJnYSBSrtKhK06SPPJ/dx+a1LlH9qO7rrAku4OY00fvnqGCoUr+9nTILlZ+42yHYtCOd4+uMuqT
YkLP0W8zJyC6bsBiA1REKW0CVoN+5DAAuHqHKCHoVurHZhHT/jTi82yMrgu4hMgONSM1B+IJWQOB
4cg3Kkhhm2ygd5tdSwAr7Gq9OxgG+B0qJzii8UgP36ZdlVf2cjk6hLKRi+Z2y4RQXI9FR0pPhYRk
khbTBuu4RUZXoJQEu3A02OvnZv2gLN0poEoHJOPj8tDxYmuTYFGQXs56Lcu0NbnvnyBmdDVvrGVc
isL2muJhtNQPSTclCGpnMwU3IycMQ68UYFxkN1pGElcb7d91o+32E+YXC1eGaC4/gAxJpISybr3L
61Gx7q4IA86Fzj780laC3yBCx3Zf1s658CtJaDz9eMr+mi5sjC2AJWdqYdMo36r4FrIzsk2LCtEx
5Pr0T3zfBbFmRnKH/hE7KA+IrsCHnbrJiM0y3WQW+DBW1M0/2uNot6GhJzVIVgusSzOyZqPPjQst
nAP7kZg1fgZG+SzhtoH/M2FZH1ITnyb776mNMyX0p50RZSkwRET+sY/nLHi6/dUpchoeNw4731n8
5hM9oROzTREao91JuMXOo9hG+t73GylwDA8C95sxN7U1TsQv2f2aXYCMg9m1k8lHFS5Hi6+JPcIt
0hK8Y7Y5OMAJ4yPEk8BTfIP5gMGfGKy8R5btQymmTB+GqOuja7Xt7z1WFI/xokU+p3+lUrfdEiRW
hMYjx6gdiWnRS72yFfjUForSzxc5fpjk5O4I+/AHDZEhGBuJryunCCunZrCd6Gurj5n4/kYi5hzb
Ew3zGBo61GLXwSrFNe23gUwP5OFahYXV8+ODTSq33tDI9ri6BhAl7Rh+GhysHk27hXBiwrC9YRLt
+iBhw5VyhlY1eOMcR7ybQcS1sWDQlutQYuqu6VnRs4F9era9UlEriWNbrEk7WfZE3UuGejTDyLUH
ahbVXv4e2IZhnHuLBpwwsQ6nDKzdtw1X6ebiFQm8pV0kIWZ8hdDkNezohW88+QVzlF42ymppbXJE
Pr9OU/gaFaRv0GTuGPo6ajPNObVhy0PLuY+SRCp21VkJUrObycLtb97mAmeyQaS7ydqODtdpm75n
1hg6a6DA8FvMfqh8qx+ow+pxwHQQt1uO1k+L9o2Tx8iD2npobNUdzL15nSgA0epP0thMYEMT0/Ki
5qSfbLfzsRg3hqNJRvVh3RJ2voTfRJkYJ5s2ZvSHEQ9FThBAeglF6xJ/ZYo0pm+CkzyZFpVEBQWN
Sgvk3WNoHPnU8cZ1xoDXgfgQoD7/9pei7F+DSHfm4maFTlv8caCyiCQIJ/7iR5FJbwo/vDI8jTLD
iide++HqSBDLM2h5ViG2gnhTwKrKYj3dtRS01HIdBI3i3pIAHNqlqOagBBc6tAIsg9cek+wP6LWO
XWuRbm20dBxNCtIXf6wNB6mBRSPPs5TLB8CrF7co7OEedhkNSKlYva+0prMsB1Ay13Hvf9z17Dnf
NoBYRxHxhp6If2QG0nvWcefIg+m4LTRbZBr1sYyl4L+/Vz0WqHhS5MkANfAcoS95A/20x7XoAC7z
PzbWBSljmTEzfCYiKLY2stbNgTRtZ2JBhqQMQmRNooZigRLCl8klxgmJyyGFBqDL43Ca6SFO2wdL
9au6n47orFnETAMgk2ogd3tTVpxZOsQwGH/muON1Wfgp7a1wXW23ocXsya3Eh6MDO3wxe4j06d8/
Ejos98AHDyp0Iy7zYWEMzMY5cvoAFujWAfRjnp9oTwrZjxmm8eJNKAMX/l8QVFYB/TTRTwLAtlZZ
t+sRzTvVvRzmk55O7VhlF4f8nrrvEItgw/crBTdL2FISA6YnFOqS3uJFsaDLFi8X4XJUUbSWiz30
69pQVHTk7neDcXGwGjbdYtxAfxKUItQnGJhqLXoAZ+Q2ZZUJ63gUDx2WRliQao4pVi3fJsDmtbTU
G9U8sUUrEh1JBUWy1Crx7VGA/XrLOv4GwKELA6k83MxiKI4x4BdkTzlA7518s91phwUFyT8o8dHb
fv20rDRf6TtUNvJFirezJpJ+dHReWtrXrqfV7MnavSg86XFskKj6P5E7j0aZzoVZxGFc9FexC5xX
EIjfTFfIjMUtX7VNOtXKXeA8OPHU4erN956axGaGuJTLzUddIy82kIkB+/QhqxXmGvEIcLjzyaAz
zjr2MT1Zd+Lf7fr82Qy+jQpvlQBDDsU3KW7lzp1qmA7Qd4jhJbaw88QJlSLUzXz2a8jjjgXWYYS9
10f6hdjCvioadiIemuHpyM5UBzsHmLUwiKwJ+INdt6hNGD61EnmD/g5rhZWBX0gJbfO5dZPQnHvU
UiUi6CzdTif238UMwwB+Bd6wo37hXrR4W12MHoGMkaUYdv15KM9sY7DWktmdfroXja/KQPZ6GpCk
RbqbWxUyf5o6r6dTZyg7cmchpLN4UBnFKiklwWbyM9YfMc7ztHVEuIPHG+1LT6N9SZJTodPOidps
ePyhui4ODjREikOITMgWmCEEKJfh/vPLXZUwjw78l/0WpXi0+162KkuVohJvRnbZ8W0F/yrXLHb0
UC97sPdPQkNt5lsWznaeT/GUyM+tB3lNMFGCLiiqwOjiwkE5fyiINkBCNZOVFg8srjkKHzFlx3IJ
ifwi31EDCZ5sGJJs5hyASeWaP4R7yoWMULOUNkez3FgiB+sxa9ptUujyqrecpfDmUZu9bX+uJVa3
81U2gGHJMD7F7kmeqwiGIdnkn72KNnpAGi7xp57frjM+CpZ1dDhAW12uwD80hP5618wwti22Bk97
J+mWk2Q4RVOKTo2DqtyRcUfnu7uJjeNYH69wXn9Swh7lQEenvd8gGzOPyPzXmYUSFcHurnVuxky9
1f5EemB8wfqaS3mdbur07RqecAI4uKzaiyqDEN1M2QRD8rTzS/aSRtm/i1lgLuwH36+Xb8pJRHmP
ylswV7SLXLM8PNV7dnBTGEjMNKl2yCz5MXEfC0q9YWR65DFo+tfFs/osHTnR0B9F9x8UE0ZybLF1
TghzK30HzQIbJewOMcRQlOPXLCNrvPNXqJ3mAKgTyHrmT8nTVjVKuPJclNNby1Vgud6SE3LlJn9C
x/ywV1WIvSLtYuTd1q5MAXx1aCai3Z5XL+gv0ZE4LG03AZTExwalIsT+UZXXo5nGRvlO3C0UwpLx
AheqEtRl0+wTmjbHSZWwpQWnmM3cBuWcJGYjGmx2baT7/HhEtTRMGQw7b5v1Vu3EFDVfDdIgzLLX
D36vk16Mo4Ikl46ZiGMTPx9HsP0Zu6Vi965Is8fSr0yHRWP6IPEA4glVflJe4TYthNcrD+tptAvg
gYL/JOteN85Lf0BWKyCAXu4yvLVOPFJPp6lXocDEE5785I6Xb6+lzU5xyc0xOVoVHpCkaKCZ3AMu
77SYKL1zIOT3bYMbKN6Zuf/gZSDsws4Ewn7WCEHMPMCPucOm+ExgS8KRIF4gMxrmw8ycYMzXt00G
kfdTF8/liKt1tBJqArM4gCLxJXYJUncBGk7swLVscmqu44B+dU3SkrbmoODOYKNpJs1+QzINEWxa
3X1i+9NwBMOLM40Nm49ju/Ox0fkDgp3o4UM63l4AWUwAhJPCkw9urjDWTmviULSrcLzXuFd2cACa
yvAEz0sVH0rQ/NTbN5hMq8BdMmPZvIp2avAaJuCxgviHE156N2alWQFgzL3yVcqeYOc44isv1VMK
xZg0foXm+gXhdYH+wze65bDLIgDbah1xf0CtBH38xByiXueGWUis640U4vHQr6XSINevYNYoBxtO
SgY/XcAl7Y7N8s9XY1Eijxap41W7eqqrRz+uIRsKfSs872X6RvRCj6q647TeaNzQYp+/StKhJ1Au
j2/6cgClv1x77txc4W/nYjAOxMBdzCpvbu0VVBL9sQcFP3BkT0QlO1iv0Y72h3adNwQ3RxjX429N
eqTaoBJCZrX8judWy7lIpM3XOTyIjSaNzk18JKyrCjvbjbBQEIl5Mz7EQImf69gOqecll/QRWAne
AgB5G4vBXQrFRy9dkw4gJrSCkVg+sguaU9lgJnJkVYSa9CLw1SINsJu5wZwMB3KpFR3SlBLStly3
7LERVLwLpIMjLnuIelxJholeIa+HNbcKgrQEMVYxdRCbgmOwZGqqf43vgU4sdnpMlbaWOgx09xwh
kO3+t2O1czEAdhF0CGXogNFD8NSxIyWjlYhIiy5cqCyAdCICe61iy+oZu9hCS/UlE3As7oisUp0J
y1giqSOInZ/KmSGsjBsGSv6g7gCp1qbpu3W+HQ87a77MiNQoSsQXA75AmgsQp1AjI2zf+aF5s2Vk
Fc4POvJejgZIg/NB1AdKodLyLdAqCdVQoAal4MNlGOTf3IrDkWQovLx6b38sm/SPWTRclGkD6V8G
WkC0FAOB89+l1Wi7jCjyK5a0sjkchuzeEzaTpP2qHZK0YQQiTW13otPgSPj/ex+46MJRzdxu6o5u
Eu7SvEi7nfwDdoilQer1TQaNkNOX/NEDcx4INYg5qbytPBFmV2p7AxomiuQsrUTra5segCJ7eNdw
jALbJFs5WY21rAivR8ycDRt/Lo44k55PmegoSzkRVwczEAJFCXM+sxRjktM4ser9/+Dztm3rhi79
RgxrxXH5ahk1RUO/KPM3+sUDTCj0DivCea4/7f2bYnaRgI/cg1TZWkfRq8CGn7daru6ssYtrKMpt
bqtVCMmgfU7As22cVWgQWglidgaFXDX6+jdB/sg1NqeK7ch+Aq6mEdTdBuHVBnnR814q0epmfEBW
Eiv9TVArhM+CV/OZlrCNcTPa1viv0yvrlwAQFFVwnpYh9Po30xU1MeAUWeQloZLOLIFfgIgtMMu+
h77hyaW4qD7LsCxXAqdEqZLgj2XzJU4H4Q3zt7kTh8AqCzCbbPewjy4RkjM4KqcLlY9suQNJgTx5
LysByg0TP/WEP1oWRr/2WfgYQjhq85R/b8O3LXoyhTPYc9jX9URjSz/2E1vy4QS37XOT41LdUXR8
n1I3qgdQkSIAaON/amNgqxV1zPmukjEGHj0wX9nxmA1el2rpeNCjsm6NxWUIvvSsPZxc+0itDBfA
5riBqiTjRSICImJixwKvPVd+knKLsfE7vhWeCLDakOLMFYGMNTsMpXZY8q/yZ/8S5T+aWFOHVPHu
4hVHGe22vuLVW1E5+4+K+L4ryjxFiwXcw/FhdeAwGsJS4C7nDBBzVTCF2u0TeoLq9pH1r+QkuPyB
tM9y7MGCeJpuyKFbPlcDNZHHPkR3VLhzhORKqQ0O9A2A6qdmkY1fmqd/RMIfK/6yIXqN2Q3w4YRg
HkOg2UEKm6wbdDz6MPFjR5JCGo/O9r/VemHiJXCPmqr5VwxsXmAbJlNFXM+WYG/ypgdx/uE6c5pu
pYSb27qU680eZl5fSngSK4SnIGHTJA6ETdfBXsK2oUPsogFZM+qXvwRX7x45db9+nPW5sZM7q+kh
InfLQjvklcHkZGTVwpqSJT+HwHUT6DOQl5Y+PH40Cmik0W04yJfEKyFWWPzxghqSYCbvbNUneXzM
wpo2jfnq/RKLFbNUdOFkQeulgHzwQ6aWJHlVHqeYNYLMPhYwcIRgjZCJDhf8gN/2LHNj8kWoPidf
vrRkPTC58qff4X7ZSKTlTttqtrvq5Vu1cXgD9F+M+q3tiBIRCPoZq1hsUxDpyoJJBknrVFma6k5o
BpnxlYMonMYd0dWJnJxYObXMYhHsSr7yL5B2eq7q9vyjNrpgfk5LZor30y6tr2qwa+8KoNy7PWNP
TbbIe1rlefFA+gdzA2DRDiYExVXR4cahag8SfeAQHU1lSxeBa/ypobZnGSStS488BAMPTebLVR8b
0WZw35C9phwY5HM1FZVS1WzDdE/ADbUKQxJuxjOnthCeGochnezyL28+frXyETRmqqTPZzUucG8n
fg6QQ6dBxdZmG315zkXJ4z7QVeZUiis256eGobzAs+DZFtsqTA8E0RisVvQs6BoarAGkz382/ZHT
xMNUBXi+5Asm2NdO6nRs0r937hlJpt6wol6SW1HZilKL8anKsrIIeivOapCveqlQ1xUNrQqfaaFY
XGltgYQjaUewXcdWl7/Mte03cKOlC8NR86H6/mYIH62CB71uGGY7U789qiTNbxRzR0K4aV6OMgtA
yTzOowE/teeia4mhn8sey7BRtu2tiqb+iaUfhkFrGb+Bwe6va6xavHgBSOjjMpGeAodfRGOiCRNZ
03XH+XKP1aCR64R0Ua89wetQeAHTDzd27eMS533Ku23LGBkj/z4cNsOeAWJrf+LB8DnMgd/cI/x3
iHtm56o5m3wR7681zTvgtyIpKONA+eQG+giKN4GzTetT7iCT1R4b9DSoyq0m4IiJbhM4dSrXBsO+
UclmvLy9ANA/WboYmJnxxoNzVJVembI5F44K8E4zL44zzCClwub9kif8J/Qw/Y27KnBd6QHkAMO8
wKflSPuI1msV5luLKGVaWZHlv+KhQRc0Ek7wcucTO/QpWeAYAIlAzNnvomKg+1HKsI1t07ccIRT0
0tGjfWvVUioflMKuQyN8tvG+yUSZhLP2MUz14jKhxUKsub0QD+QsSyU7XBybiYGyqh9swqiGkywW
LVdCnvz76wwHmFfPevDXNLMFc+iLCaqAk3lFASXX/9bbT3rVmzXuIXu4jE+68+K5eys3Y1b9Kif5
P29uHZOY45Ic5rWJNqnRXvk+4OqXMMxNzYjYNbQMZcdwAba9CVuqqDjoAOgfk6Uyn9hkeypxxVBH
z0ra4pTZBEmjBHtcHr0no4EyllReSeqvqyWDPsJiDbrjwtKWBuZf2w2dALJtKJ7xAT1LBQ1grAnE
DJ7fdcdws6X2kxidxzqcF3Zxeuc7x90OYy2RlAmAqtoW+pu88mnHfYK+OJUWFQoGX9bV8dRzSOoi
8cx26i4yl8QVuMPgAtf1A+ikQi+RYGc+sLCH/fKfSXvrS2OBRESkoZYauVge5fdF8clDcrgZJJ/W
iAMHd6IdF2cgYE3UsJxD2jdzJSTAXX+UNH8Jjh5XIb29QqDt0ts6jtcvXC0kM95KFB3RlbQQ+3so
TikdU6EIpqY7R4W4UI+9sGDSSFm+kdStf/CPaxXM7zIFat31kwFveZsK51vfVFHJhTIJx+0pdFq+
+BfH5VFVRkxGrd/CE5cURVQx7DIf8qhstX7icPXWFmsLej8Jt0pu9Q02ohOt9bXFRpUa+GsTEBnF
V+FaFUOVeKLBHuAOZL0ZP4fin6QiyGCFSgW+WtIZpVCjdsP/lyyXD3Y66EMb8vPUYABwoe29Dsmr
zjq258HqcnlZ/54ZzQS6gb99OgM6jXbsZidejjlqawOt/iCpc9iJhOcNfzDbc/jRs6nq7HSreMGz
6WOLZLtZuQWFSJFY6aD9IRKD/uHfJVqrak+VILVqlfpQAZhZ5ZyUNa+/4G/MqONsdY2Socq0kSNm
vITFoOClZqLTlNuDDfqYUfxOqImK3rNyruU11lrr7B5gMvD569XO0K+KfaprfqtjRW+tKkFfssT7
BUk/Y+7sXjOqufjjSVMivyyS1CcsCNbV9cqTx82QkT0SFlAcot/z+bgAyrGgFhBpj1ajpk/UhOls
C37ki+jsvnVpIAE63NQxlRWXErav3LWIckgrjw8pO6XV4gSuWkkMX+aX0HGwjxFqez9k+0okb+Of
XkmTf4p9TZMSqRSw4tor2WCUt/t+fSHWdnYscA5vOqEBw1ug7S+WgjrwjscT4EvfqZWYHngX/TTC
vZ6OZ5Cz+c2PAFNDoBKEUt1t4G5IhjIdrNkkmiXvfn9YD/cNHpDQAvYNKMLBYqUYWhJWV0R6zQXO
VOwAqd2AEwhKzQPMi/iC7/hPpirI38vL2U990n+leLHVGQi/Tar4dhBVnrOOjaYqogyIIcsVS4Em
8zIEdwQN7vre6PEBAQxWzBDsOVbXkFjnKLqS3CxgYs3BFdDoKlgMicxSGdFUsI2+I/CLhy9osK8X
Ax4KeECwCZwDPG7pFPCUdbkyQPtsRzeJGsYULdaBBTNg0BbC4CEtSV4QyE0+iKcitIk4LfpEYkD1
f0trQr5HtjzDvQTx4oa0O2I8tjAQxwYLCO81ZBfLuV7pywmQ0DihJOCUqMoV4CZ1BuNoM2Zsl4wP
61AAuTGCw2LX0DrZB1I1CZsrxj2I+l/UkL/P4SDsB8UkS3Pag5y3Ff2TbV5nDrT6E3L5gebvDCgO
UC9cYVHVM02B4tWYt6MSRiYUaautGhTmG0t4XyNw63bJ3JdtuKFLURopUD7qJqlyxR7jzE2Kl9VU
nDNTE6k9y7jt1nxAhbgXUv05JITVwtiLNdqersk57D+hWkNhAojqCoMPGhRhFb105hzvLK+Ck8YD
iUaL3+Rlh6AN6JWuROYtlemyNKbE4uPvAUaa8u/j0nOfHUKKHu6i4dKAg4hf3Ur9QklH2vHVXmOe
CK9AE6er3M64Za9kfnxZ+gIxW2tUFmxB2e5nJkGnR++gKJ5rFP4Deo+mPjJIfFNaN7UdOrz6+YM0
SI0AGNCJNOL+6puJiGHiIniiS062S+JwKs+UOTt+eHU62rABp8sE4CksV9lpM/g9PAXSPOkATLoc
rzGZMExXXbvTVR5VQZ/OWIQKcss31AVSbKBSth1G6nlFY2earol3JcKp2VgJRnAVXvLUm7qPZvUl
aKtEQZvHskfYtqQdGjOo4c3Vfb6NeXT2dA0EjZR6vHDZyNzeDt3BUJP2ZVc/T+xN7sIsXyAThoGp
kKfFslmrhxnt9NQQDmlqhL6Az1QIkIUtd/NbzyvzOUmE7vyvbFklyH4RYm5RZUy3s0852rXGEFoc
gO5SKjEHCtKcwMdwlCpmJRFXka8ePYSEN6V8hOK6dRRBK9VVs5/tbgyvZ2qVn39RqG1AnScGvtu2
SnFXwRWHWQnfv4TKrBPuQwaLeTR6UqV+4PDscq4KRaJxwRYJVl+9pYhPEHaCozV9X3K7mFTbOb1U
97viu60Wb8fAiBs849JAZVgUwm/pL917SiPBzA3l0cUe3ym0dvaN7j+85+trFOrhb63f/xuJ6CrL
/1ktxNtl4AyfWHmwr4qUYjJ9vHOWQDEqGoq/Wt7cq3eF7UWsAY7Wir2MhaTS1iztsJqMlA3fzukF
eTOtZiuJ8hFvUrXjyIt6f4/tXQBXo8EoER7MuPPjCmAqo6zYLhsP2dFAAd+rSNGYAkm+Wa7mmy6G
CjfR3SwpKI8g9tE7Iv+HWLSpAjO561NWB8hdQfQ/JHJrh+RP9kXYMg2feY9Wj61pTzj5/GgYJOqD
UTOUoG1Ads3vPfluppJwps8xPeJpDI9kqfnmWnN0mk4IKTQe95HZUI7tDBNF2c3QWTK1qxA6S7uX
QnrSciFFniJvqKPhFbnxqCt6o/VQnnXH9YZ8e3EtgKvLUNEiNlfcvPq/PGncsBEplT3rHy9zzesa
CJuvuT7tEm1AYoh5Xo4ZaxCILA3fMUEXu/LgpNass2T7CKWnJ05wAL8bFgMuJ4yP1HJXIonwLoQ6
hlB6pWUWJjCaISQ6f53PzSrGd0t/DVRR5qeJR3bTMQvvli0BNvxKPzYitJSG6eId3M8NK0GxtL++
9eoBh9gmuf4jezla7Uapc/0iF5278R5jfYOyj1NvqBmrwFpUgY2tIouUrZh9BDhxAFf3dECuU1Zp
7FuO3RIFVMfQ2rWfbnDPBdUaVdkMllBjbZrV4GrbPnrBzJG4MYAcSFpYL3Zabh24/uJrmBNmqnQe
WOTSxcPxgiA3UVkJYkgTB5B9YTCKEmgzsSickR0SMbIyAM6cXLwZwVzZgb5f4Lv+4Ui44DmR6TS/
XD0LLLDNpfyjK0chDlexbPr4+zReK0+pIBoa9LkqJZzMkz6c3xb/S89uT3/UNworQoGzz2b6Jh+I
xILd+kzo41a/CjzAvB3eQPRnDhrxnjov7DkF4fgmw8GA0JAiRuH+n8JW1yz/HfKc+KF0BSlBwL4S
jFRrAXxwSaQnxXRVtfwvR7sPCDJOmoc+PjBNEl45jZb2MW97pjojg0DJzEMaGHDb6LdsrFXOAdw3
EelRBNvplAVWLhXav2sziDeexDiJ1EHUPoohrQ+pEpGJPNfR66qgw0zn3YPkHbopgV8SvEOtd5PR
SOXeLW/WvtbHAJaEQMa4zkO0gaSQGTy30gLUZE0Z4MH3e/XCDalLpMVni8GwRFM6sWQ1vzDy9BKh
rHkIBY6F8lAJ6dd86iKbWqyw9TeCFJSMD+qViyASZ9F2UzGa9PPbHnADWqBCqe9ie4DkBejDweHe
kY0Kimx9ljM5v4fdjyeDgcJUMQPv4uSIFPrXw5vh42vSauPX1+ChJdoXSMETQyxJzVL+4WvwkuiT
th3fbnTKpwwnKJ58kQowBdUavepxF43LPr+CYCmMzk2DvV+XhgRhyCUlmvKKe+ANYHziGfIeCn02
JjoDGajaEo1+d+61KUa3R6B6VbxY/ncLpMORtF8uIoF+30s5F3d7HBKayaeBsHpUGPnRMIl/PA33
vmrXcV9pqDLbMi5EXl6jgxgrgXDOTHvRyDdxZl4Ed7QP6JMlYRmabdn6LCn5yG8QoFznLvy3LHZ2
of8ibV5ikHwFJ0B2Kw3os+n8zljs36GGjDtSw7FeTY7tnM0807Gd5III1OdxlW5C86tyjfAcVIOC
Rz28g2U7dcuvZN+k57xYt6gQ317o3hwg691/Qd2HGMZzyKH9kS8QX4i9K3EKgFPnWOBUmNvWCZas
4/XoUrvZjkqb28xCoo8hfLx9nPyEzWYC0jrzxpb/HIYMadkulWyhSmSUMhYy71zhUcFIIqzom+Sq
LI5oByKJNTOvDyAsh8civjeMgtNJkmYqC0y5btTrdE8JvDGpIYEhzZ3wHrYt4glpbZDPmVuHopIE
4yFl44T+ofhczESNrVDzZd2foG2ncbqzgzS3HtK2bDhSVaCLtAVp00XNdU34Q6KxKIb5YcY/dMyB
+r3J0TffolAH7WZogONLMZ78tjxmIIQ9g3Jl8eJcZO59kynUHUMLX0xGeagPug65pinkQ3Sky9PR
07J0bbCeSH6WxVq0e7HzaOQEQij/i+D8BZzb6KMB68LVuXDEbJ2VjQ4ug9uhA1hWPYFjC/07SMn7
6zG2c576Jnliqb1+eEIN62oeiWsCXogJelnD0LMPGCf/gbsKi1KAVUT1UkEWWhkeJnYqFqZeYY9D
mleE9mEttTYtbkYrgdSCQ/0MJjVySJL2kJOkhk8TXvSNRAG9o1PnsDqGvB9xAkAzv80lqF9MRxcF
yhy0Ex9sksSlyQXrtwsVIu2gChuDQBB3OkACTqJk+7pVPtifPcTlbmnIlNndxLHabz+5peFjSIqY
e+YpAO9etXANO0A6F35aaV405RdPgGInPVtLRMlmWNaZ7yR+XEOkVJTk1rTaE6azrXb3yCOKElT2
m83JDorZfXOGjmkMwqbHj5qtCxJz9JvbbmdD/5Gor/W8sFnuElbDYWL1tcVEQM5S/kv7e6rw2FrX
hiNIjv8Z+WhsIv+FdHVSbrp8mrMjFoSSDA1//xdWcN3Pjo4IiI3mljBhQoXmfJa7JbaNx+27Epc1
+hk4ALs27KXeqlvsnyDglDnBvbeq7VL8HAwHkgXJ6J2otjy7lZDIPpQOz2dEXsxUbYuY24QU3W78
itT0NYeEGo8bcASakvUv21w12L0t9ey5Xo9f59GdGKIfTBxhi+UV9WWASo2D9M6v/7SvlbMZb9rq
8ft/P2LxFOZF7YjnEruEiWgxxyIYBKriinXYKgf397wIrvvY9J8lZtAKTX0ADzD0CW1WTzltnSdD
rW6sgsbw5u99JI5UaAJENlFTPDAlb9bcr2lEKepcjTp3gPY1HQVNuXIq5715D5hxTQAIu7eTUUAC
BPVEf8u4bvi0NtCBVzjT4nsnIfs7lvXbLcoPTce6Xbunr7/1m8OCIV3yfn53FgtD8AoOZCSQey7e
zytzzhAiCLGLvoRQaIeYM3RlRdblT5lj/IfJ/357F5CtkPdl2hJJrO935gLGp1ZM9PRtfTZC9K7z
D8K+Q4bWYNdDD8wrGsW9vwCc/rf7HbgL5a2LCGoEc5V8wurY/9asoXAwLC62piCyYwUeHMZR+Ntf
Isc6lOT4rg+0klKpTKDe1FBi3CfIOKaym3kv36tFEiAbkpHNH++pSxRWbaFN6sWTUJI9Z0o9vNni
7FDh5L5miWcHaAKSEuZQtftv+8O7hLKKSAkv76R8o01Fz9tIJ7Aw8anxzOYL4s4ZvL400pY7zwab
MDSWWdOdJbW7fIdJJA6BHfQplNUm0c90beDdkYJwcufqhIdZO6jj/KfVc1s20X4ouoXNl5+md2bC
xN2Aagd2LvP4BpiqoudvCEYjN2MVsmMDlMSbfVqQdo0RPhWIMQEmjyd6rLZHJM/em6QHOOImT201
Glr6X0BNWnA0ynJYGnvHtbglFCpRu/sSkNmK0gcTiOE8vqt8jJgtmSbB3vtz/ccP9j/Ikx5b5hE5
Y1KEmaIywIm43bKOBJuhCrZXIJg08wc4KE8qzpTQUUS0Mwkv/xPR5+E944Ff+eAG/nZG6amlA7k8
41DdLmWaAf1oRu4JlSeOWB2V6+lsfBunEjbVeFN1nMxg8i2fG6ST4e7NdUL1OTcbQtOH7I1CHEsX
cpo2+0QPLXBllRVuvoyYmTXuT+Pc3/gp8JSuJnmY+Q7qSAo1I+idEuVY7AgpaA/O0OPAiXxSYf9F
L7i4+U9ORAcrtSeJXheKVlYX7WlnEePnFA9VYu/k0jSEZWeDQxNjII09fKolHl6luIr5sgKKvo89
mvuEw1VAve5oqKYekl5zp6dcrNfwi27rTsASX6wzx/ldfqwvQJYSIovv1f2Wn6gy8Flm6UUvZHcy
AmGNzvKY197zTyZsSxMjW9hbO1lAYNMCEuiURtwvwIXktrhVTEQW4inbJJGeteyrKgRlHyJk3Y4C
ObuqzEv7xCt97fkgBkEC1B1iBJt+oAxa/wLX3G173hKZ3zcssqEYptn5F5BcIg/qx0g4ba7qvfVX
XCwx/SjmXeve5cdVBPdMxe303Jn79IndIu+icASGvzbq8qLxvW4dpWvWj/Quc9OmbNtIhr1xG3FW
WPoLEjdd5LYKR3OKzVoAA+6Qz7dFuy5vdrxoBOnfvfQ2MI+NBywOepf/CisRmgMi24QUbhCEzGgN
oaEjxZoCc4Vxb5Xfx4ULSBtzh3CFhwu5z5mzoTQ9qKQ0UG5Gr/WPBTdg63QJpaJrEiZ3qfsmMkF/
mtzQcvGTMN1Axi7V/MI+Vew2T4kW4CEWk83hupyRE28Gl77YIUvSOH1SOs3dYKSwkqPFsnGLjqQ0
eh8h5yXy3h6VKK+pWffXIUirnGOalB9IMWXqDKdl4ZKi7muMYxrDEFf5MEYtch0+r5jFMOIdulcK
sWnn+HHBEm101h4qiLYvxAfK4+9IhTzDKotuyg8lUkvuVxB69u8dh3XNhv9BOIOyh5VuOd9MOfb4
c2QsqripGm9mF8qvW45C7QtdqFMxepSBbw9QRCwtFuMFGCr5ottDwpC42ns+Ee2j8/5i0ZAgyQRV
b32sxAffwjw2fGMqH0A13h0PeJr+4tvEI42YWmHLUrCYJqgcyfOgTLbAIZxf6RRMeE2x5wiKGjpU
02mySm97aTcROPumCF8aWwRgFcqDADfQHkUp9MuEkuOQDoi6YjxAHKrM73srvHfLZSWMHRxZBp1z
GJiF9+V7W/bsp8CT77JHv3RGC2Ig6MWQyzF4GEyHccPUDquZQp83mpkZgD1MiloDC0aj8ZakXZEz
ZDIT8+27Vl7vmQySSTtJ2A3XaV9STurfwkC1S6BETwC35kn8JTMlLR+qCucqWYJiStjP/A1bcETJ
DpVIVEMbHQ8Z7FqoWZPIyLD/BRD5JNBTERfLeAB/C1yjx+ZZE0oWFF76ONNx7znId/C7beP3B28h
fYBbv9xN/7qO6y5Zs+gRIjJSo2N0w0Zl5PXtbjvL3PlfvBl1z7sxyT5lwL+6TZb4eOeWuLJHBBTB
XMP6XNO58xmYwQ2VSyRirxRzB5e+Xu5M1D98kdObjWaq0/Lcgyn4wiX2fkKtTq6l8M9Hc8wYGN/g
e2xjguIljYKwCQnIXRf6Qg4IStuqnqL0y/boS1X6Kta759jdTgcqWLquzubalqwY4e0eCWoYEiDP
ddvoJiTGykERgJ/OfxpaRMEDved+RyEK0LKdlHpksc1ZplKnKx4vIXdw32hpVbkUVPmLLQUIr64R
W8ncaGVhGeO2R+F2NhDJsxsnHfNQ9YMbOYfb7pprfSZhPY+5TyCKl7J5je2NZUpSkSi01qO7rPGU
WSJVxLPK7CE7zLvLpwncTnzDqdjmhjMYFgwf1eBNXnotpMd0dEYnnHn3ERyDUEH6Jh8IhJ8eum5V
CSVjVhuwGIYTyM3L0qKeJuF8HCFl0kPGTnOHI3IzJvHQYsXcowZkypw0pxBH/QEyongfVicLZaRI
z7zKdgYa3xO5GjyCjMrV4Lmstmk3dpn0xjaFcFK1jpQxsn5xEG7pjm1oifIExT/nKev2vGgk93rS
tOXRYzUDZ0HkaqUeTzDhSOQ1QQYFMYzTNC0WN0kqNeoqwo8CMN0UZqp6Vw+dwYyeCIvHpItv8wWy
m5uvX4Cudb5ldetymWcGvLLPnHaPwt9uyfXNFSkUZ8aA0MD1NLvaWn8mTVJRQga9iE6MMRQSlttU
ZJFvMBzRQw40lNpWgZEYKPkQ7umVrEbSynON0DJloT8cyK4ay65cD3HF88YiuSWbzhMGcR8Y0c/M
TKFu2T/+y7jajhPj1KQDA1Licx1BSDn24YUx70niA8GIDcO3t5RVW8qTzLX9ZKxRbcMs2GMI6Ree
lifOOgj9XsFx8v7UX7KRtg+oMfhPjyJbBU1H9J2HAUl9MgMb6ZPZygAZZh4mRRf8jTUHhPG2DQLZ
WWeWMK1DOw391DuQAeygzQcbTZUePu2l42xm16WtOZddGbCETu1nz2vbi0suZkVcfglNkjShSvSA
eagiemKLwbnU7lh833mQg4px0hX/LtlUg5ibnMIwsCZVu/yYJ8JjtfX/EzLf3vfrPfw/NQsiEc/5
tcEzr+tu3LxLRkrD52HJG3nNe/gqRcZfS6C/5+yLvxVxwu11C+ATTfQeVG7Bd58QGvTY/WtLMSuz
qYpZ77WSmN9cI7TO60EAq+ECrscLoIeRKMLieR84sX2UFdcuHfjBIhPXYGfArMoGoQ65BjB71wXY
mF0YX2UVxubCaE3KwP3lLGyMjepcrPHqLkKzYykFqe1t6x0nGFmK5Td1qxrptZo+SrHQjfYszWIf
uetipXauTdvcgimswgeD8H3Mi/Tr9UyIPy+tWe3qmE3BQ2uuKtbNPDOCPmvukf8CgP+RwT4p6tb9
ZWEqdMJgE9qZ19/eeBPDkclhyHjeyMy3ABt6fqplpJkE/t1FNDhw0IT/WEFVj9ka8Z5TRY06XQkr
2euLrV298JUvx7iy/VWFHDqVuj7VS74IUXEjg0sdcSNY65gv2CfL4C58tjpfzjYYGgvPYzD/EO3X
DDHW1HjN3zzhF7bqBNyFivzRmRaRWi4PzTB+47csCO2Dtdw1W+YgTXf2yGecXGB+na6UXHnJ5Ud0
NcDH+mDR4BQ2/zGdZxM1z0uhr/CNkYpBi1/aKPMwm1UHsey5qfngDpeQLy15HQz4aCv/Py/F8M5p
lG72Rg+5IsnG8D6JOfXtJ4aQIJ5kwX3355l/rAOJlGt5vVoLL1RsBdSr7QJJpJNVb60HENjvnzPr
NrQ0SaKbSQ8ePG9pW/VL8pfhJ0RVMwyOwcroqLkC4VEpcY8oZcoCXUSQ3oi4LoGsHeExKqvH7lLw
W+p4Ht3L/8SthNYFs1EylgEHt1zqaOAvQ83FYN28nDOu1XcHdgBQKzwnLoWIk51zU+ObNlWJMytp
sr3Knzbl+brSh9VnGB4MZFQ+hEKua7Jp4xS0BEWIcHX/wzbXk5xRP3YcuvryTwAicpe7umH9uPKU
RoVDnJJ7phSkdx5ELKVzGh2qsRLoe6wO/0n0L0SFV1wLFLG5WG1AsDIK6d7TlaqA47QFDxW3WTjW
FjnGmPqcN7RePn/bLzBImrmz0RQ3BhF5oYKuotuDjjQa5g+NZtR3mnyWUoi6GHkYr67SwQYYYm7F
Oe5DQonCoh42Dud7mwS2X6q6YQKhV2wX7I6sP4i/FSKmWZ6MkVZg43Lf7XU1gRyGSo2+mw6u9voR
QuZKZEmem6iXc9rTQi/nLF9PGRu/+loer2STpWevPKPAcUOlymXTSK/mPuiWsaHW1s5qRSb1+Z4P
0dTpINgxWC6749I0Q7FVs1HxPSLvY87QttY9+3VgBRJHBRF4Xu7dZ4+qPFgSBYEi2B42tpF/SSOz
Qf4w6YuQBYNscx2wJjEXYEfr9A/HWjhV1VtzlpEDiyn4ajyuWsV+V3xFeIAcekUlsZZFAEnUbNiI
11cjlGRV+IgHl4pLNDrI3gDBBEx0M498etTtcz7y9yCelF4mJlNJ/MDvyUBX2kF2w5eTcwsv7f92
GvoUZ6iCW7iD/EdJCo4v2Y4DfZRBLETyN45bphe7AjDyh2w+ZHzoBpGN/gLeilRwljkHjZgyrLQT
VU7D73lsMlbX5QbFgdHtm17oqagxzSfyWN8XUJE5Xb1sSFlmXObeI2hGbb8rAdDI2rynLnx1icy8
12LtRmRwhflbETg+36Heyea4FtZ15RKYssCHEF0arNp0tJAcjt06CftUJDMPBo6S8E2tpDcdjgA0
6tx/dofBFHpCBFnp5ZgQXZ1kh+x4EprorvmOjBeXk0dfE/9d4E4Ws/bJHc6qcOQrWZ8rK91O+tm6
D+QWtcBsxawASRJpNvjecWMWXHWyqbjHal1Y6iZSNGjFtD8hOSuAjNVMBQuV2HBfkxt/Yc5aXFo9
xRB2hidJVPTwel1MsS++7SU63JYkd7eyC6kM00KjzcJH29/A+xCF4AdKwGMMBZS9B1Dp5IGdfcDT
hcXTfsmVAalvBZDjSeeeJNBGSr15KvvhSKCbHBXYFVh6BqStDxtGBi50Lukpt2gFB+Kf0qH+48h2
rfroi35kl7pRkzXUFbUirtsE8WCpoVAnChJ+hgFkJ4iwTQvbu4Mm/zudE53ZuP8jJ0EBdfBZyv4h
grCWZMvdBHjc4YDen6/d54+kKYUmEpljmr3xi8INl4tdOP68Zgx/vkLCTkS6IaZKwraa80VkyQru
MgafwPhEBz4+mjKVK13Jg9CRtYI4SQajMiVIibIa6vcH7eDp/x/JR+rQTpRl1jhVZ6qX/i5N8rK2
cBLTO8vW35BmlhLsDX1oeEaKNT3wgY5euiVAR8PPbMBERCzPJFJYtPwuHxoePseUKfr7D8qcVr6W
TlsxQ0UjQAglNKZmrsZLwbQh5xq3oEilLInNGwvthYNodEUwBeutomb4mkNzRTv0mPI0dv4dpkZm
9m7vmVDQVccBju8+zJkCQw0XwQXdIuat0aOT4uO3y6uwocKJ5bn0fIuY09H39jJ1hX8WuI7kREY3
/qAvb8lxb0KMEmPSiy76IJmSFcbxcaSnTewv1o0iubpMHCrDsyc7AmMQ/01Nece72qNz+EvckZfj
BnFcwUwvaaLKj1wiUGiwxmRvC1IyG21RztVF36Qz4GhfEzEyntZZLQ1EDjK0K4+vxgqQUdDTX1BR
+GS+KX0V5Zs00RdupHA+t0Ul4OItHxOpoLS2+OAeCSh6yR2w0GnmX5SkiQgzLT0+b+PCn5EVjzQI
9DfPyxtA7qLJRj8WkFIhDzBhMPa8m14qrNd/Wnw0Hzhj8vC9HR/siGl7hDBNlsCoj5ntAwelvUcM
PgbSWbuhLT46HmKDWmnDgF8+6amhczwmgDYlSQk64RY+vsZ8fgXgK+XvfXjX6XD2nTCRfAzwZ2nI
TM2RUZeATfhJU5Y7vCTiApEyichXR8m4mrU1E2MldpezOq7uoJ2lyCeU3B754n4FKFADbEv2w+cs
h3ddHD3Xe+wW+zov3bh0p/cqKwW0IlA1GX6tzRYlwi8WLipr0h2JX2dSoEBEe90s1ypnMZaTzIPX
7XRB/pvoGyQTlEKBfUtoFdonvx0VOZvmjsIH4lOODDVxhBffQ1f/OYHt4rWvP9RQx5PS3m51tDCa
AAQV5dtvnv4JfSoLf26iQxIuLytVaC8+VhDtPb/CYVDdAaAB+x6itxL7CYdJ2IjAIS2m4lBjs2/K
QUiYybdsNHtKAzSGAIZZq1sgK8ROcYI7mmcX94tnHT5TSAm5SULfBIA5q3gfjBPlpgJQrq8zdRMf
rIgoSlrjPLDp1hWUex8piwRs4RQE0dB58VSOFG9pMmtqip86jS8sTx0PkMsR44GBYiItRBBghpBq
K7xHgQbBAHSi91ut3dQ6VLVFquMEXlT4FL2iXBPPrN2892ysjv1iAAM5hjo7NtxLN8g6Mn9KNlrc
v1E9JuaXr+aFAfOc1nVAwqS0362MnG1bh7Mmt7G4Hklw8TO8U8Ou5KKhO25r8BJuiAMH3i9yXU3P
KJSWLZiXSJ1W8tFS8Sz1dZc3SJmrnQExvt/PLhxWou33SZadZVl4RPHi6vUCCN60kFMKHoppK80H
rXdoQs1qOPX/zHMRG5gAEoJheBPmVYwGEvnybN9qRO6joxBvvzzA79Hyeq/E9PW4umJK5ZMKZVWm
oBZrpmpwpKuriYWSpU/NDmeIK3p0YDsvBiAEYJg+7ldP6uieaKRkwGSqSk0FwkWUqoMoPH4/SyHp
ha+fu4acQUV1OAyo2l2QD/8UMjurYMFTJefKxYm1quKdBQqkzdV57vZxiprDS9Tdt1CWNZLQGba9
WHLjQHNJD/klnuY3DyfDpmA+0FOKuwq0sMQli10cIuuIcJg9jMR/al+UK4udQZDxzDOkP6edxCQK
gBmR1ToPZs8tqU09GxtEizKheJ8XqvpXeFDceI7KEF25bbNYgw+uOKp8P7bSl3G6KRuhW+2W+YoD
IFlhH4h5BmhVZ0rekwIPUSq27MmWmiYLgsRh8bfcsQ9w5VLnx0OnbkC1tlToXsIy+C1wC9NdljHU
rqXkE1bHs2SHGb90z/B9iFXQmaqRsWwfH8Y4G5OQEDLjXhtRTka8ZK8jmPOciIzZjLle8dEltlvn
Z5FPfIS2IAPP4prQ6UqmCm+BKdPh605NdvaxzXQlIueZ4a9zxGhSlK4IIBuQz3uPMGmnpVbol67P
BSi2/Q/Hu5pyd7TLzPQXy3dE2EZr4ODEqyu2uxEZkjx7MsfJ7kVK5j1C0roocpHG4iSeRCkKPF9o
NPZDQNyGu3KvoVrNyCaZUYpLOX1ZH08nz/ByNS5Cmxbg5qfNeG6qy3a/RcbIoT0gamOChFg/ZOfh
chcvO60HofsU71iihziTfjDcy87cLepJzLYysYsiLWn2Fj+U4azBHZ1LztHVw7B8AlnJu1UnPJd+
3KymZ1xlDl7P+sVm9+wK5MDBlgvO5YXE8soOOfeTMKwOpbVaW3RAIkptJ4Gw+yjQ/vsfUqV/03Ur
Smw/e/jtFdWV8Hlt0/5JKxk9iQvtDdhqOI/B9CBaSpy03bLSW4j8HwZOXxPsHzaLMrxRevU1193W
hs700npX6xCDIfwIiItQn9qHoV4v8qPyJdPuk+Ez1x16Cty3EJjNV0qCyJyHA/8iwYiOF1Xvb2it
5CwkGsuj/iqaN/ci7vNhmoOiMjQupMN4pI/X/nhg1ze63rSstd0c1I6xC6q/VvSS4z76A/MZ9Xz1
ykbMTSkya7zUGg5vM1CtSGGNjMKr+vOH7VMj8dFn6MKchlUKEmpaStcRD1RcdFjZ3+jbJeRQCOJf
/JzmHIyoEl+33tQ07J9tSO+NNvJnOAYizD2e6pP7887a1CQI3E3PkU8Z+UKjvP6evxdu8JqGcNYL
EevWBJx56iP5XdP3sNq7MGdM5uB+Xex2IU5ir2fg2ZWJhH9ugbwbM8oZngQMHFoMabfDm/5wqubB
LMzaSCQKqksipxysigumYOi7vgIsnxeyvdrht0eJ78JxMjmrr//c/Z6MFa9BYit+xgg12yPj4r4H
9dvsQTGybLNbXRvA4NFp0kGxvNiq4gobtY5y1yOfKcAaK6EBQV3k+zUdnyw6x0g1T8C+qDYdyhss
Xiiv6CzJUVhE5k3Vk21QgUjN6/l+0lm1FThO8zS5gda85V4b5LsQkWyoCmfkIdEQpOOsX/Nv3qwg
TzZs7luei6xU9TbUZQyZuHYUXuTwXicdK7DRYxsJOmP1TERJywVjJIA7PSJ3cE1JNeKMA0SK2OP8
Fiv1wDapi0hTntE/a6MwG/z39LpBSs/P6esMUE09/kgIuBsS5C/ImjFi0k0qdbzIr0mTDisv3NqK
5EgdXceJHvJZi+CSHStw38nKlMxv80JLUtuNzgeTIdo/PIdib1FRTwUHHoMU6gfJGYlE1EFXRLzB
bIijcEsjgW2Ps9sIf0+nmaSQ99QdVvim2nByGjdsQfrw77xEGZahid9CK3jyiJgLC0FsTl5Du8tw
oXe25DlUvElqXSPThpiqATHdmSuVJCb16i4qM6JeaMoeyxlpM4t5L2Ts8rLupJZq4T7WSlXCG+1Y
P0Nb0Jfa0b9VfBpOGKBPfmQZ3HX6HH5giAck50SuNZ2NOn4h+F+tHAvA/VZDMtBE2JIkHmhVol0d
T39BiGR8gUK0X2f9anzo7ckG4DO4IKCNueFKUBz0xR5sbO72y0OT50FgxbxV2VTrZWdJa5lIvdIv
YZpcKsMt4blVYtp12hBZjK/VqjimGgS6m3Cy+//cgdANjmFsQdvv+6nfX/NNYZ2F90PPp6C+amC3
uB8Byb84Iu/d6qVbDXUu5gpzdq5Iz3J2bL7FyRPdDPg9/P/ZIMHk1eH9GyxJBqzsaUnRavXLyBtQ
hjvIpIvdBZ8b0LerPM8HiS7P6LKAeyHvOy9X102kRx/nXhJYX5Myu6/G6hXtQSieivmcLpQ0nHnV
E4W3RlpUM+x3cUiu90BPkxWnoPcMqrQmxOH3ZdP5G1EwUGiIeC0L3L+o0cEBbGqv33KVTdKweZwP
kxMkqT8DiwIPjLXanxCkf0u0oaB3oMDUFYGxUtdikIgfVQENBS4wIcZ7TqAhoEOBE9zsr2Fhbux1
RCYNc4cytZ+qAM4hTRAihzVziGvXvjTjd/RaN2WXRxjCBv/WkfLMByqMgu6DD+3dM3fecaomtLFO
d0unLJImtiJ4GYlE4paTnvMUXw/pcLSNQhxAsbx7JNJROmbheviubckCZsQ/ERxpxvGi5b1BAmop
txDUVvJBOfDzEUeFpL5MHGXgLGqvH/8RIGtrNZKvxVnPcA+foW3lm9MHwxMnBQPkcoAwz3S3NSUF
qq445KIIjfxCViIRz0GlceaSo7pVoRgot1JxhrzFjmhEGaF0xsJcObzVBff53Z46eN/st8ix8mAG
gdkfgzHEPOn/MELzOraInMIIBEkFFSKCXwWYX1c6641h9WGY/3CCQ0w/D18daPRj8wQ2RrW7fVZr
jY1ppl0i5rQLwNL+g8qDUTy0PgRwQ6BcoOuQV4HcqTHLKGLUhMFpAR4kdi75Ez9PaJ2dAwQ0bHHs
dnPOU8F3+P4scccvDM+dYp2rg8OeErTPij1+msBdz4eK/cpUw61qhWG38cvZ6EUn7jKNuUc/3c1n
IeSgXGFZnhgtHcSy6B4udgiKeeYz0mz+hEXPw+T1J5GI4h0ZRe6p7+W2WkkpauAknoVP5IyZDUvy
ga54/iyyFQVPG/zkhisL3GVA9CqOgMshLx9YC3c8lMEXmMy78gH4HUfC9/I/NLxkGelhS3sJ/CvE
Fw1JreV25xEOywa7i379g6ZCwMa3XVHZGEWNjbwCSexqCDEqSFyDArki9j9zZnukKZ08L+Dz7qx4
RABvQgiuEbxkxe+fVM9JEEJlsrpIPuwZHK1lyjAWquXJCINoKjU9sEr+JobAe3GkiZFi3vwi11DV
N9shBt709xk3eZqAWGt7SC6YFIrvRKpfKbGrzxZkpfp1UERydmUYjypDPly4+eKSZ1J3mJ7Zas+i
egGUaR1x+Kk129LWffqXwHNny0ancoNBzxRZd9brObbKQDXmROpJbDnEzl+MPVFjaezurKFn7mYJ
PMYnHLPcietBz2KYpywney8Xq/YGFgCjT4vEKL+n98L9+ehNjtn7vaGy3sIMzTKbrnao6P7b5g2F
iOvrpVxOySY5P+TbmWWuoMX/ll1RGj7bMvq18SmmSq1V8Fxurb+66HjGgRPI+P6FiWEqwn7jNrPw
DKKtT2me7M4EWgK8okekUd/ryXh8chHKz/t/+ZDg2/5sBx+/799nfOaZJ0V5VpIrU+ZnHeQ7sDke
XhMpetdyGZnr8ZwScWJQJcL5RL7KmM0heTQ37e0zrpmReEUbzme9CGtloi2s87bzMCXcLjP1M3qA
NIP4FMBUwDSkuN7Z3ioNlPNmQvbby0GZMQFYGoZC9N8xJOFhUFHUy6NzwhlZo7VAXQrzkcoV7Vvz
SAnjzqKH6GsTfw/6NTYIwvDEgP/XWyCL+aOfs4KrUKVVwDA9GWYafQ6tlt5GxjBtcCGxanocB6kr
IfS6kaQ9r/AjfRztnUX9JJh9nLTVjQV+5oK8pz87pLkNhBXg3De5wzzrcaL3pb38tHDSCizbN6UK
HKzuVv0m/rhMvTWBz2IsYXBbf21BgraJwGKppt/I3iMBYhfztxp3EjshQMdUsAvGUnlMuphw8UWx
PwwxWz+kT5H4hdxDY55Q8b18PSr/hvb6eU4QaxhhGqLl83sTXZTUJf2+m+Pjv3wK7CNtYsPKHdcY
FvSp68eN3bIGDjavG4BUdkJSmF05YHAiohhCR5qbT9VLg2NdFIS78u/z0By77b8nBLwKjmV1FsBx
hQ4q1Ysv3R29H3pATabIfmPdWVvW241gp3UZFGnZSOU16DKly0Z3wYRi/4CL0XFoUqw4tfsVLXDy
Gk9MHBe+7ebc8ewzZHiHCHq1Iggbw0NTkSA0gxQjbueATvOKDc0EDonPxpuvUFjE5mgcJDNX8VOR
+BodJmbBeiCsiMks3pyp4xTUPYQsMWAq3/V9rgju7qErP/LFmkGzQ5XbiRM/Y+YCjlGc4tHL55jX
LF4YNkbOABQDB+BLxmbuLTa9oL94nu95vLPExIXMXVR1TljVAJTbhMOZsIVIMCkG8q2CAwcTjMZV
DC752xWpRB6wdU4R6Za3Lb03QczsfBZZBYAS0bKZV1j/u+ZpFTc0KYl9HoY1bW0xiCOAa+TjrNnf
OzoOebJelr7aRoeDHcXKeyvjVdAcPWut2LG0nIAi7d3PQE3esxh9h3P5HgxaAvP9oIaUwCVDxR4O
l7KvNZjvbWyDy+D7ZilmD1jjmisSKvQ221e3/LIfbIrdYNrUkys2wsK83mkyi43+DLYLWVCvPhjL
VuQxwi8nUAkkUCM4JV40F7RscqBshQqdrwYMc6UMKKS0TvKtWyR+4oKAjE9ThcTMIDX71aZfur7o
J1JqPL6Tjyw2eNz5LCx2wtO8CZEY7sSlka7FaA7gxD5uqAyVLs1/zVetIIbkcUdvMEjwkEVz2v+f
HxN/thLOjVxilpZVqvIOYJJXh7ZbNPldT5UFQxeQFqceZUU5B3HcCnCsFEIl5BflgvLZZNnzL9Do
X3Ge8j575X4JEvE2ydShbd9VPfp6wwjcGiiIoG2YDBbqQ5cNquIAxbSYZ7cSRm+M8a8wVig9F9rY
EXM/KKaL0CzNZaN6RPieF7KM8WTlhktEnrE/yg7Qyd8+m6pvhofJT5S0B0S7/ZDCilwoJt9A17NK
4oiPQTklgDM4pYNZTVCNDL4SBeiF01XocyxY9vAKjp8nXOAIpLup68jV/2WAc+ENuu43alHVCgLw
eDaGfnugbx1DGqBT9tvhOgDQbHpIHaGLM2I98qeILbwhG/hkMLJd6q4J8l97aIxZWdw82oEYw07N
L3olvKn33tYb7uCCmUclAqTt7nkNBWzLAwR0kSyy5b12xigzNhDJ9kFeJDlqAhq1cVf3GYNUTCn7
LBOq9tsKUfOg0Kc2pQA3d8d1pumFdVgWSTD8ioKazMYD5sxCRDrZmbMoHVwhJpsv292SssrXR97o
2PCVZIGe4BrEqFXE93D8NvEKVgul08FPsEHcBQzFn1vEnw6/49SjHYGdHGCWjYEem+UA34NGj1/k
XbqgbHEVdeGUt2m4sRzYk6Zto4IrcVF0SvcfrXHkNfBLu3oxRRYJ9rYBgiLnRllr2ML01HxMvo1e
Rh1CjyPuryBnsqB82+rmRUsaqqvgESxz+LmWdl7mpSYyuNHgRaNefOW37VjEJbfHyjLdIauYMeyz
+YcUYfDhqwyJMn/A2yw3sGGQA3BvhuRTgV9/N02kuUM3Sy1ihG2eq9TyMzXVY5LsMdqCzM932DZs
vWMACBSyPN0aHJHYS+Mp/aLO+VJKg4hTswx6Tint9Km+AW3PnjIA6CWUG7JKcI+FVFCq/uSmy6Sm
EHVL2/AGyux2Q8qIryn+c6R6WgmJqd+4SkEjUcd1Jy74nemP8exA5srwnyTnNrSpUAl/+VbidcN1
8YI6lwokZM5Ztmm9H34n3QR6Oswee82M5zLOwQPzDKICoWT2h8mWshypXwbU2aWyCsPoJ2/FHk9B
H34etDRVAlycJ92y4yQJbrgpduAnEHQIA5OpBlv5t6mVjgGEGVk+YrxiuKBOqLEjI/YoxXH3Mrgz
lJxpQ9psaq36DYt0vMSie5IVYIjJfyNzDLRlKQ1JAdW3v8g95uFj9WI8ZCWUQ2B533e1uV+Szgj9
LZxPcNwqsWCTOEtu1wLhdEI8Xx8oy04GmhdnMVXtnMiDsGithk499l5I4cWExTGFG0UZ9wiOe03+
XY/+xOxbNTkyfeZg5i0gz16zj/ttLjIO6B6hULiiAWzMHcmvAbaEgw1p//ZaP7qIlnQjXxTHmLZQ
b6I0sqE4blyJ/lUZNh1ysYERAyIiNDRJ9vXoyB4YHsgYF6aIYIWuzXFwC4Sw6zAYaMLaM0UMiKpP
Bo7aWQaBisYd0cpofds1+wnN7yAZt8Evzqw66Sk0gLYl/xT6F6CeRBwxvW4iV8xcSIAa/w6Lgxk+
WjjKkpdsZPIzdqRFzAjmkuhaIDyADRwIqTPwAci9yRqHMatwgKj+gYfcUVnjZuhIrvuwzb94jhSZ
Iw9toY4Vk3C9dRkIM4AVASO68/SpHCQ60B82qqQVoegmAUyjiiLJNogffl+Mr5hbuu3hn9TyALmc
TiHOmOTjYoakrI3DSgB71PYywEwsMofNv7C8n4dlzS3AC0OVotfHHId9h7vJuyioma+PSbNmgofD
jeWcjVgcQUu21SkRCqv8qn4z5RZcj6wZMKgwiYAFV7gy6le7wMWn4Nc0sHngisziYY3+M+KbI9Sx
9dhVdsw3W2pqKVAryScAskl4V9NISWCH56ZQlNWckShzrTLMQLJlo2AtBQSm3Nkt2Q9Uz3zHwyLF
OVcG0EPTv2DSfajaB/pR4yZOrffFltANQm6bTDKM+EsOz7oDkVksrCUIg2lC4AFgUZx9lKSWjyuD
Vw/C8bJCnmIbn1F7Izh8hsUxUccUcWdQOuV26HiMKX56x9JXfsXHNp/keJJOY/ZfZhYjLV3s+Znn
U0goJJJrXMmpTWc9M59zgNbO+xLrbEPCilv9SiitE/rOZrlYl9vpce9ELi3Tvi016F0hieSk8JZm
c0/nkTrC4/pujzNAKEolytaXBo+uUXfKWr48T23y5tAXX8CVzngOFNbSIIwkPbalRIAGsiQ9g7/C
l57n6RCM1Eawq1/7FsuXv71kBrkzrWvYl2iYE3m9D+rgRJQfKoRqLN5oP2ioL7zhgfZSLhJYApCA
AdIaTNW4JfNHWPR/qzEkYPBMaDyM5EpzAQtxsXpiXXShM05U5CR5+qGkFNskT3rwUOEeF1DTrks8
zWwVvomQdvn5yrg0/g3lC0qqaEN+nnnQ2yhnJIu+QJV4nNmQAiGk7VdI0JlrKMVgMMTgBEu/HgWM
myyOV+8LiU5feal8f/++UHeJS/jECgmuHy3JOlnjnDeElwvOeI7qLULZ0XQvdJZDdoHAfMWl0MME
AQPNCdj/G4O5Ht3BleruN0cYQc/JFcL7pWsZW2lcCDM79hjuOJrAp7X8kTyJ57LFs5Fp34ZGPGMn
pkCPmgnQYVuw5gW/9A08vQsKhergn/hyEuJIbHhifiUZZ3xrYr49lODV7BLFt1k/+LkVhuifBE+G
T34mXAFrPShBxJd13WNkjYI+9XckVW36mq+xvDUPxrXI0P8HBKKscCQ7PakLtCnQOhs7RaE3O3VT
zXQc1F7Vj7uUULTUkwsShbjmj4zXK6m0H8Vpbu8fIzTRbOFmvJTk7n0aOxALHemIhl8tHpZVxAVZ
ta8qukLDhsQRedJnk67cdyby3Jx8Nv62fHC3YZTM2QHO1QHB7tK+VNbTwom0RAWfaqeczGn9JbZQ
wMbfu2/zxCDHiUGDUV4pIt7q37aKkL//8XFJJBu/iratZQtv2YBCR92A+KS4FbgJ7VVTaUJfd0T4
iFDjMohl0tXnltS7XDTI/TEHNvOJs7IflLkGBX/0H8gHtKebbbTGnzkvtRwW87oOi+eFhue4/dIE
YtDqhxxhgDpLMFWn9FA/KMPOLXej/NDdXbzvPOXSMwFOde6fe8p+BDVvJwsp60Ah5WWyyQamhtev
VuQLR0suRBhUyK/262iewtWveVhnnZ0evmodxWiel/4d0ZN6fph3O+BMK20AE0azwgfYfqYmFPXX
uXUl82+fzbbmBimeiEeSkZsLEwo/Bj0+chb5EXjxAcUQf8J/OUQaOMkZaDQE61B0PJkkzM+9h5aF
78TB7onvxfdxLgXp7j6BUcq+fnxeU59M9pKUPeiFPrc+9QqFlvvBL6pKHL5T6yQqaXvPtTgEiVMz
CD0KJK1cszf0Vwy2ahm35VxPH0Y9VH5PyN+67gsxft/7VgHl3I0KLf1UpLw6s3QLx4hM8qGRi6FE
EqWL/MrF6ncBEaVcNO9WM6qJ8AoWMUZxaHGxf2Xu7mXYVe8gicy2Ps3WSnAmshj4uEtdKGMa3iAJ
Mo5zKYd5+R83PPtaUPRR3P9oruLVog81I+juLyvBNy3yt3u/CyXqYRj7tVfBmy5M6vxAgaUouLli
c84DdUHyO3y2pmtLpkIb6Zm4VchYOqoFU3D7GbriGa9Gs1rOEsbwOgLC5hNMKGpGSav3n9RVR60m
MFpeBkSVhyo0TLsBsNcFBTi2i0D9Y8AZmLXqegYvyEHdPx+sVcmFyTEjYmKLltB30LOzRhia1b2a
+9NAo9GmbRYJTyTZMB8RRtBmsbl+VK4PrpZTYto/bVv+HBvAGBBsl2cTCNRg0lIyqcXUiqruuibX
gA3WbCMImRZd9bJAv6D1ULZ48WF4C9UIfUPRY/kySv+5C4ygOijxf6OO5d7SAiCARSjuTma7Y3TX
k6cGAnZ/mT3S5xIoF/rMSEBlXCzeSY9Ddc6VgTveem2mCZWU1DaQLK6s18Wkx41zn2hLWvr1Vf/h
zGgbutucnI3Z48IfusSYaAPPpNtsXTnWIY0lgMHv7uaKd4kHBKdDZoBIcqmYCTUpi067g3TKTh5h
72wSqiNo7P1aEUGLBQCM4vEEyoxbuJeFvoRNF2l73ZyL3g3WD6FhDTRnsE5n8SdAyJBWpT0woohv
4VYfLIOVCbBK/ovUiMWAh4mZ7X2+9wPMSC4LGUrvxNRaa5CnVsgo5r8kR+XEvb7R4JTJldvlsG6V
j0iCfEXFBuRbn2N1T2AXW//ZDlayIbDOk0JyTFME1O9Q8NWNLGPN/oYwa6a+IUWdLjSvSu2nPrBM
I/M0ZxwBEnwPTG6Blk4gQ5grJnyJivxHIftHfXojzaQu50DJGGR+RU2pOs3cxSqN7TfmjEP/i118
gUZj6gEpyP72tEkPYmG8w7wVWda7iP6D52noD1biZhqrINbXnJbK0gXKQxYM99EQZdTUBdWJ2Hd7
s1klh5HglyE4vobEgr3PHQjBjGS/icHc6y2mRsspibIOGxTvxPdxe+UB0YZzfmQAEoolSMmtceDh
AhuPRjN+D4EDXJm8NyyH3hls1kP1jpf2+KoJcNM6qwJRB75hANuqd4A9MOZiezbzmZidsEmADaPc
HbxAqrmtsNaXBS+F4+Z9pAF8eede6PPgRoEEKuruvjsNOwKdIbqas6o/OVPYsn5gotWbMwvhooXv
4U+0YeCYkG2mZhyl5JPDYfUZ9S3eM5UtA5Hj2yDWhGyuUJDteYzFq1oVRBqkAYqlahPdTQOP1AYK
BGDVygAHiK65WQhDBRW8266fwXtuNJhYwoH/Bxq82aY/NJGVlmdLDR3Mkkt+lG58h2HWrzi1c+jb
OheetzeArdW1ELxwKfSFf8+rXXzUQhepd8y3A28fXpkipaA2ZoFUGIeRYS2Izq70JpFBDx9NzhlH
5DrWqbmJ3bBAaYj6syXIz8Z+ca7eC7c5Kd5t/tf2HtX+jxwKJcDMmI5tn+dK8BY6SjWlchWEG7AC
2hUwmDDfOkLgnq5Ch1XaRdmEwnCYPIOdGg3CUiMQHjRcp/mQon5FmQItJtvq97TCsjXlyx77WG8A
cn2JJSIUmO/UGW0WhFN3n7KxrX43JST9Tqttr6tBeHYuF2MVH26Iv+nhqQRJ3q+cR5Ok3isP1vxt
Rp9dTqSCV2dJ6NohxiVBOGbuLHRUEbme9XRTSVb7MfJsEI/Uc+322g+YIz++5+n6O9meUFNrLvE/
6Z+bMoVEMt3TZ/QxGA9ZkRWmk3hwj0RxxveXza7yDJAHsxl4+QYdvLaHRTlCtKnUjD3WzKh7MGyM
yxRWCOfaj5wMs+DGqolRRWaEBs4kMIpJspjWCSDbzu4gWoGMiT8YZTzzcfzO+k2NPRNjHVMaek0m
4hGMqvAqMU1+x5EVAzUBkcIQdapuV7xDKE9UvtFw/kRXK1f4GNCrVw6shnHgzCK/H2LpS3ibi9yc
hRL6xTbyG5DkkMuNfJ08P6OHAcvuC63EHNzMshsDEnw+0V0zAYUOJ4+iM6WhcPbFCGr51jVd7k+y
60yYGV/hFbKjNexjarI8aZYIPpJEOhyRYVDMFm6FsD4X8tbRIw14JKvJVD+42u/s+6leKSs2O9Ub
WLLHRYryHzGv4SsxfApC1dIEf3Mt8hZ0APSY5ArhE/upRyvcui4HCMTN75TuvD9knFgSP46Ai468
WkJnl8S0m1baUcWwNd+j9Bfa1fPGZKiQpUAhe4DTmtL6QnIOaJmCwE4kxaSTx7BP/IM84Dw83AoS
Es4miuaIGN7fiWVj/1n8wPyD7B5rpWLQqZHQH6Vmf4z1/nLMxKzMbG4YVqwWlj6L9QGh/7Xfon31
aL3Ro4wDiFbA0WPsjBcqG/ALBqnhxPVEpJ8wYegoc6fpPMSiz5aX9iG8R2yDhhbQeJ8KvuQi9y5S
mKPMPKc2vPaTq8A1MzKzjrLzpsVc+MIiZalJbaUWPLRGucVWbgU3D0n9l2XyiBaf4yrVYBC1bTG4
A2RHxZaf2NXqO7cUaMJ87q9XUmG10MW+uogXuu3q5luIy7e6JUvctHXJEqqsYtNaDcJdxaASb/iq
nayCs0k75Rb1b6bl2wuhm2EiQAl9jZk/9DHGYwHX3KrdNnDaZIYsqjm4DeNzRUZSDxBxiskHrSOC
poXQ3rXmigp5Oh2z8kuccsFzqyAFES96QQ4WcyetEsimo9Ydz3bc/WwWW+k4dnJElbHVtPk+8Lru
7390Bv+jA36Fo3Lo9J2wz2Dazr5t6kxQj7+gUMG5env+sOrLAnusyPhfukfPNxniTzJIRsUVZoDC
Hawzdyij1A4mFVx0w/jlt5hRiBkEK5LjBCplzGvy8hKsFE+T/CLJKy/mOnr3pLp1B++XsUIUZxdM
V5cYA/VzJKJ22ZhL5NQAwzhSkolWgsEBm3TgNkY+DGk3rMQ9n7DKVewYHUBtF8v6lbP3Fk/ZV+gt
dnqQRI47DXDROrsTjY8Bmf0DnFYnbQTpoM5IrY4hKGwpunzI7WmG/eX2jd2YqlBPZYbhGdBhwtgY
CVxmDasTKz53fREXmVLrXI9N8SNagF1VDc/ur1Mw2s0+h73c4l7z7WBet16AYvMg//ksCwBnGtNJ
tuZHz2Vms2xw/H7TIz4rBIfn3xS32tZZnRRG7m38tpkfdosLnWBsL84CU3YmBt99L+pXSA+nfscf
sMWH3WdHkzeITFmrgyHUJWlaJEdojM/tugMm73u5eJLlmXkWSxH2ABSJdRnSSyjCvA7YjtV+VaCf
2WYSN/svSf0CcXFsxOruD+XX9PaX81adTcIZcY3cxQzH5TzwqIrgDJyi2sQ+GlAKz4AaejZk324l
YjHraA46Kwb9w3Fhnoi19LFB4hAWqq3rCGHIU7/oHm2A+kxxqVPHVVxsWkTddWXClbDaoUnQs2lA
2zBJEOCbgFADEmYf5iAinhfEa1VkXesWjG6Ep+xw1xkAOkdXpb8bvxtggHF0b+iva3ghx0ojfl/3
mqPS1FTL39X2GbrvvAh3PcDll15hoZLI2caf/lrvSWrIFU0vdROEbdTlt1rj8hHAWHQVwNUyunT9
OG2BWcFO8b//vCmQ6SMeZjSVsft4u1KEqaz91sfBAO+UM5We9Kt+XauDjUDW+eV8vwI6LOTI3mAA
eEGWn5elNcGiQh4cagwAdm2Ejk+EAmnPVUE6/V5C3mybfgf6I/W10c5oJPh8fj1J5afIMMyfwTMn
snIowV8CzvEARoiz/uyC/y6xXKzHRUHWdYuBALwTrL0h2744lh1tfywgLe1MqwLUAZDoLrxtLsVD
u5Ed0VN/E0DFA1pNjN1W5nEwo9lgdb29PaF4I/OlEHZQkEBT+yewyun7b0Txn6ZkMDz2PsSCeHWZ
ZwoQWZ4QbyfwzO2WG8umm5BGR4fPnebJBEjEgg5/ThzxOaTddSXHsYH2ePZUAbBllkvsPXlUHlgi
W0RNEm4gFn1X5pVBJCTC+upqbfbgYoC+8BSOLzW4HQDrMItWEOqtanbQA0c9LzB/OI0Hra0xXcsJ
qwkn19npx6R5DExUOc5OweDomQs4CshGtAQr9cnVNRo2Ynm/GuPdEVbx4CFi5qF7cBIKQlCLT78i
s57l/qVz+AiP40dBGYNrWoUHuLgppsKml2S/XzDbaFdi+od/NrGqwRmKEJMbM53Vtrc7RF7Dn5UM
Ml2gOfFel9KR5qePQfyND+2Dg+I7BDAuzW0lneivflo8kIJNtUCWnPBpOgfByqbnGpLaUllTEmQf
9TSwk7PlFYaQeMPRTP+tb8HbygLz/KTCDpNhl4NdUpPBQHiTy09AMDFcSTTcQmJVsLEui5OzZHQF
35HDE0TVhU7NZrXb4mfha9ow1ZR4f8cyhzdGDroP39rcpqhZGlCSsY+kyQGZ72ew9RZhFqWttKpo
SbtGZ3ssPcEO9nBBjEoQsn3MrsEE12wjANXrqQDcTYdjUFGHNpZJnJBw+LsHiYPm4rn59OTOVIq7
GDfI2AW0e0DHPzprc0liIgg5VYv9GsU1UqRKs9jzKXzlo38Eoc8sBIGCpFd0jk/2rhU/spP4uzqk
cqd8Q2mDG8kd4sWfFH2Pw6XfGFufvw4zOMR4UT4p9irHSH8X5r86D2OLkY+gHKXQbtWp3DvAFjNX
B3maDieJASnLfx0FwNYarMHVbo+twPLZvUob/TcQTND3wHTcA2mhhwI2RZl48xsoz+if2w1Ji0H4
/wAJLPcDDaKOCZQZNMtd5L/ASJ2bjAppDN8GmjGbcRfl3qIEuXY4icQOgwNe4vJkKftGPZmsx0pV
4erOZEvklOHBKlDvwIuQEybWAEU2EHTBXUdFRniLYXsOgHvTWetoytRX52MgopwU/VE8zoeuFLuR
+ybq3Ytup38XovrQwFnDcW2qUIUoO5JwqtQDHyokUWEB0uIU58wxhO7NkfcYfAfDS6PcBtotH6fn
lM5IkMbnR55ogz6uhSFkckLXm0CIVP4mHKnUjrGFK2ZO95a6z5BPx8XbaQJrwg5fxThmTHjjfASU
JD4Yh8mUjYpKjePyDb1Kxpp8jOGzifJMEhMxz2RDP/Pg84Wm78UNYO3FzULzzcQWlBKxqQvf0NiI
ATkVm8B+jEU1392gqf/lVcvJLVT7Es0d4B1GTGPI+MXfdouGuSDnjKBQtdTGBONLl8p6JZyoPXKB
1uDxny6ecvJoaQuCjU2GfFrynjNQEqJkYfThp7kSlKU4YixRnwina2KDose+ejt0Rghp8jRyMqvr
ffUOhtD9RlShSN+RdZnoZeadvPJ5AWK2yolemStF5WHW9BdSaGsFSLgXEfGK9YMgwXonx/ESVfUP
+/kiwy+44txm3R5z3lezxYzi9Yz+UmSXgUAFFzbbfSN1kOG20WtRRu5jnqzMF8cwlM9CP7p8soYJ
NvdbKLgcPaY8qM6z5vim3P8qiHu3+YzyGyEx4/LVSTCk267CfSGjC8hiF64/NbcNxJw2/Up9KyKJ
CrfNn1s2DhNo0wHqaBfD/luHE8hcPuC3EtfgGx+v/pGWhRPoLykcxCxLWmmtDrBExguxHIayvBrv
3LjVofAZwV8AHXas7/VqPfAmcTeahS7c+D2YfiC0zLStGpuzz5KxorWNYyvNepYbPHtxXLsVa1F+
78vFvkka2TuxLooqWpzJ6860LdW8jjSwf9/dOTvC+6PZqRKFCNLd5SEOPRgCZc+NcNW1jQ0jdw26
QPGgCgD5qVaUZOOMEMcBs388S2V9R78G3ExhuEA+WNS4UMWmnXUEQNOHyXmlSQf9xqdqapWDp6sx
rfh0TnDdraENf8uFoMZUE9gK69QQ64/Y2sdmcUKfCysv25eRTmURErdBx2T9iaIhsMSdOvTf9JDa
Cy4eZpynE0tLi5Bh3QSiTO6CIBGmowJs9TxEnCYZbK8IW+/W9vDJDhzeK1Lpe6Lu6UynF+AkwDhA
USdANRyy87hKNcXYownEiWQ0dmWSnRrG3y0D23b/7J/f3lMkfreV4HAxHv6Arvc55rpPjbcBcsBN
+JtNM+O38k3jYzwCv5AtRVzgW4/+S48cuxV91ecSDNCmIghxZkpzm3+Zl5WwegejPMURYsW11XgN
o6eWss74RYoyeUMwOmfsSJYil+kMtZW4i4AOxzjOxGu2ja7v6OcAFSST0QdDZL8/t/DDE4NoY24y
E256oGH8SxRxO3tTr8egF0b+Dz4fgZdziOea2i/aalZrgQNAlSqifJcLIWyvrQ764r5YWKCY3ZPY
1P4CJEw4GTniQr4ZAAycN1RZbBsh1rpQW8o6ROkR39GegXfpDcughqh+jv0cpmOmFdylH+Ka8mSR
ewhXFskTPXzk1lxrQJh+/wLzT9HFVpVh2idN+pUpk2NdhzMCQkCUgor8ryQ3Dd+4CEZhJSd4r517
32T8ndnasD4geA5UAbRWRuzVKRduCoPRy5vchwPOLyw3FUxHTu5q101FS7c0dmhsK183SmwKXoCA
PMZF1SlhOcJxWi7Fs4ujdDgkJ1kExCeMZZEUhjtmZlFxz/iu2gik0/oPhdv0yplnbBgCbA5wlj9S
6M69ZheumoahaNBBNDIqmoLl5XHYWhBnDBwM0lMpjTjIi7iGzfVVQqhyyjRoMLW8kwtdOKN+xGU6
TQS61yknGJ9Mu14EO+S3jDhdyUQXzvoAa7Z2ltPWkHkrfkEFjLEX3uOl8j38g+LhXWXGtG9Em2i6
wyvyDVKG1s0/5VStP98qqF8DHIUVVcs1MncFWouE14jLw7GOpn8IBarSe38ryItr/lZlcrOMEE51
zDjHG3cxWwBQ8BxgftuzFjhCbqJzDYxBzqZoOn2SXLoxAOje3hbdMFaEQNQ9d64ryQsD0K7y+sgn
2L37Tt/pvl1Euol/z983iKcRmBTiYKizRoon7UqgYcYbE6kloidhEkU+vtcMCGZ6fAnoKvntVrMf
jGI9me5yx7AC6qxKZCC7Kvq4XoIxsXY747+3MiWydkpSihsx5cC+NMZartDmPR/pkColp+li+LAX
uAUA1x33wH9w5vLpBl2YTrFDwIGODvLef/+aV6L4viwxiVwE3li+RAIa64Etu9X2nHCL4ogyxnSz
hMFsXVOwa8JYW3fo8EvkF2Vq9KI5laLoQObT+hODPn3JviLgp9xx1SDP6ufmnvQCUfV8GL/akWmB
5t8iqwVlk+wFHRMW0zO7co4RdlG0bf7DG1dAUmBWNZF8ZUHbr8Ua7S4SrUGXMU0MOUzziAwX91F3
kZ0Kh+cLhnb+csS0rSq00uTeD6PWTbI+32ZnpGro4Jeo+wWTtwJGAeH6EDuFgtmvVpjkuCX2rdPc
r21FsBTm0LzdGbyg3wECR2aW+8FIXg9hu6qoZ15OgHsp9APgJANKIcDQjW1WWXyzJYP/3wRV8KpX
q7k7bQCWCvzi6UTgSln7xUlIHETCovQkiQtqb8TJfL8gSsbQLkbeXNgltCKC9RuQ0gfRZTwpvzYQ
lkz882IW12zEeDn29ICZhs0SVvNM7/ExCUR7+vTGN4SJ10ynavasSUFDat0+3dkyKUXyigEk7H/+
mACAsTdALFd9o/VkDG3IW99/TA5Oep0DycrVlwKhbLSenKRGKrhbe9KsEUuIWVnl7Q5vB4/PY0+0
PlxfvwlIlE/zH1Tjf0jMapfOY+OK/1oVVolPc2oGJawQAe8Nc1XFBJ7dJQ51E6jiqnBG0UMakoU6
X1gpp4sas8QXLC4NqUyVSbcMG8OzTH0oM1Oa3mpbjqYnFrHTfuo+zTAv/f6DM/+VZOQmeT6Bm8Zb
qcBVcyFJ6R862tQa3sLJOOUPPr3KThX8sB3EVEJMZta3pMh6sG9FVhdqTPtR7uf38JHsP0R9msxl
xbyHP2yqF5v9GhuKnSqaoHw7K6LnOIdLrDGZ3zJByLeo7bDbjgAyhXMS0rXGqhGBjIt5LamvPtrU
WfyxJmcfhLtIxllGX8pGVae7N7Z2dsQ0A3Sd0xm3W5ATTIIgOSN+2Cs8LS6r85G/mVmvwpL6SOd+
Il7Zw6vWnACdxWGw6w+eokbyD0o77tq23G71380nfoL7H5IaRvknd6hXJlQjJfs2rB0A/jppUsDW
w99V8x8EI1IToyAa7+ZFbiUjx7VeZWL9fX+hNHB7SisAcD9aCseUwbfPbJBbG9rj/x+fpfCR1oPE
+LLrJqNseoTpK7719t3MCJczlcddTfQIQxUlKBBitHdvUgJSe0lQBlryMULeL5mA9Jwf2IbT7TjF
2c96qkHDQU+KKn7eDOHaR48haAZ/s/cU0gZS8BCdnvMs2TjQlocMQsQZMlglagiqSZtVlIzE6sOj
TqU5YNPjZPKEkcojQzCvcGvo7IqJyl2M261Buu1Cja1tZ372sZBZvwCPS2IkSHn5HVB4oZn+9eR0
vMWLV4JTaMabxFeGXPKUNyUDeIZPqwqg8Xm17tINC/rosRHeLyVc2yGtvO5O6QRDJ2TTOsP40X9t
rwVeZbEMwwmPli2JiUxa79XLHXrwegQ8xFGwn5KfLc6G69mLzZxbnI9YHPIrvI8n41QdsWxcJdEh
ugKrV0aHJ3oVZG1IPgx5iLVnjFIXo0K2HpgJoEEft0oneYaCWl6SuVQTYfyxFFQ186x4wPxQpwOM
rb7KH106supsBGWc0ow090LZnhoYm9Huyuf5sR2EJxL5/gtUMluFNMQewTc9ypIlxhp0SC8RkDcX
jTDjnCLeh978ACLdWs9S8GUf86ZiD2hC1kXelqCii+BmBmbhmktldcvOnd0CBOecei2UzMD3vH8M
hoowHF683Fo6fixHL9Exx522v6ruuyLn+XrAsf8bOzb7lBR99ETcpb5/RM69QIMKr6d6zG9odk5W
RlADU1VHwIBf+NSoJzaEliBLz+6LFFzV6Pyk46uFxJyAmq/EgpnLDCHGy2oiWqT5//pW26ZeiP2I
25cnosvOGPYCJcU3fOgZCe+xF8dLQPmSScWxnHJp2ELkOwB14A9nWU9knqviFeazlFuR6vS58dob
NYouzhb5TnH5bRLFNlsI5bjLxjP6gloaBSbPkIGczrhQEd+p0HeeJQPbKlRjtvE4T5c4Od7BU1gk
xOjekb1APzSEn93IJyQsZCa2PSbwuboXjGdWEpPzoAYxe26AwLKhaEYPOYZ0BFGvYiIMooqZ1Bxv
vyEyqjYvrSXBy989iX6uz14XADCwWnbgjKf68Q8zMA2zMc4njqJdIgP8pOgMkdMGLdshKHG7SxKB
4wuG3SqnzHjovNS999UiC/91V1n+e2X0pmdZ3qcfoDFdTVXJNhuuCGYLnscSNygefY8s+x0PjQSX
HxkDnIFQpByXvkIat5wMlIT/Thp1vKqJ2MPdJzhXGUNI9Y/1NjLzjUB46kasF+rWyyMnxcNx3Ax2
sjv7IB1AfWhPLpiPMg+Ohkdj9E20myUTULRHxcekvwssBE6jQlLMySWYd8gBudd43sC7/m2ECekt
Jg++DNn36dDbpUMw7d+RTtoJ/3+Xy7qg1bqwCEvEGk1oqV206o4nfTE98KgjhXmcOU98YNkj5VQr
MOpvUXmZlFokiEuHE3KlNaT+iEqN9LqL2GpTu6vVCH4Mdo/gMuf9/rZDh4AWpkNFm54G0MgVT5G+
C41Dnpl4yCCoJ7MqRdGUDIgg9Gc4pA7+joJf376RWJnoDvPAtzhlpmQHCZ4OzxbKV+uzS6k4Mryo
h4d6j8WRTmc6N6WzgnkXwTCG5biAYjuoT/Uh/NKCY/yhOhS3oSNjb9DYn3ETrYNgQSG7yzhcp4qf
Kf89TJx3z2p4fBjPIJGV2iP1wi88LhifDE+H/kdza8VfW0bX/vvCAdyoBRbUPa2ozqtBGYGWp1qO
5bV/bQ0+3ZR9P0zCHxBQN3MBId/2YlXD7RyzweDVJd+1qG28ujMZn3q1e/iSxo68T4X6yRsMMlTa
Ck5kROpuR2Ajy+gHbCwdgEFJk4mUCxnk8DovwDz7eyLVaowA2PzS2AM2JEu+4OUtWKSbTUBs1Xog
7nhUOadKoXYNcVnFnMVyj3m3ZJhtLPn1ciJNo/sRYnNTVb+LGe+QCYCcBFcjbOs6/rzxdmek86j/
Duv/Lk9FfxNhWdbIIF5ofruVligTZ4vaIpDPRkA1cVT+lt3ZILaQGmi/fJ8cvkoPUp90v9mcA3k/
ZO1Ym5NSC27Gdf5xG91Fr9078d+k6uTtGaPUZ2x9lYVZzVwh9wz3DEgz/AjjiEer3cOsi5zCHycm
wsfvt8nKlekBwG7J+I/2z7QRMHNWTdtUUTilRRjzr7t26BH8a+YJ+agItDnNgHeouytVeY29Jj+s
AJbE00NWSzhbS2U9qENSw3AHDglijNFUwbnM+ZMGUVnAvqZ96kr64Isq+aelz5Dr4meea/PHDD0W
p4LWGvJqJNQJn4wVPNQo0WS6t32puLQuBIH8mI+VBVv7F5JZW69rA/4iSvbIeAieISItS9ZDTBTg
HIcufRr+aTex3o5/9h34BXBFEW02AkmBmCUGUcrk+x10402vAhOlUVGOKg8RjqYMVgkMpdJxNzpy
JoC6vVPRyOzDWW3Q3a6HJ/2WD1swtF7In93Yao7wRxGx036fey2xgsgWxooTZoaycPHUHoV/G1En
+YKhyKIH04Cxxoi1sINJ8RmcKqf7ixrnMd1Jep/8jrfOsTxbvg7lLxYlFDCLFLDj3m686K+OpVFZ
S5jcwgKfUtaf2iW4ouPLFf9uEfP9kWGHLoj35XKiSicGXFbvhsN3FP/vLTe9ftZkgempmms/eDv7
iDR2k32UBvv435HyL5Q5QZPBZd+apnsQjcE67cB+IVuaA2TwK7YY07d/VPRGpiOdQo2ve+quv2WS
1I2RK9n747QvKNHpQMpJV0DLcvXM5bDdn2JsPBEyoG+9PB6RocSt1AC3Y5pCN2ik8Wglnwk61Zbn
MpF6gIAJRJqs/xq/M93lgICYbb5C1DpwXQ96HgK1k/H3y2cDRJ/VlkS/YbSi7elHLiJkvV67PFO8
qGsW/+fycLTtoyhbwp3IXSAY1MSWfMJYpybb35Z/BWaE4ZiWb56b0pTw1cV1y3CMcpGGv1mtk+Av
v0p9ekyz+HfOvkFz1QQJpDHYoeUu9QFoapq0EC4Upj+MQvefNqr7rhqDamSYoHn+BaCAv5XFuv1Q
NotarfCn5nNGIZrsPpoXVxXrNKUVqmRGXkvPEyRkeiFJHs2Zh4J5lYZ8Ww2WR5KZ6SiqX1EsgeZ4
Uei7wNbqB4TNor5FQACKrscYDIh9yDg+z4q30fmW0G3U2SX3X/azfALiFxcuQA5tn6KBdjxKl6nd
8C3fXwpz5D4ISS0jJnHhig3fqJhC9+nJJUnojZgzQW4qY5MpQqgqlXUrbmfk6cGXjRWw2neHFx7H
Ibb4nXzDt7+Z0ACi9+DtPIyZLwuRmaE6iKJ+0Z7hwbBYUgiopDhccF0zBylCJBwkmJaFg4YCovx2
3QmDW3jTyCFcceXOJhNh6Q7Un9CGYJ37f6PHIKwkNeu6ILcHwg4fY2hm+t13CI8SZbKLLLgX/7Fd
i6JVYFBM5Lk6+2D1rTMXeOPvGH54KOQKp53bV+lkyW7uj4b7MxKCNqZw4E16RK/ILbYA+k8B+yY0
mdDE6ntQDSixybQ0c3EVlr1KMd6Yfc6LPPf+DXA8Mzvh+mGD4RkDfkNV+30smFItzrFsAYAVJvbu
H2rdilMm9IVC3T61AzwVTobE18ImRts5fdRoxrUF5z4MYqU8mc5Is70NSpMpwwgt1UGzMwB7URqB
TxrDOrUDSUjpewAFZeRd3ukAnnolu4P/aA9tJlqNneb9PwW6AX+Tke7aEoP2Txw9aoVrBl+y7DkQ
cNG8jmQ7BmRvLDs5sJaWuMYKxEHOOBZ42WJdbIqcZGASkwHkXgohh/vKE073n730lRjwlSmzR5ek
l0qsI8hgbRIbzqNVnTyVFDnhxz6WdVnKPs1ceMsmTVmCKLPv0j/cjXXdAnkbw6vSckeg9ZRZEShg
3vaMF0GAAcgdkiIwVeO+ObuczvJl4FOjFefhDGsK871Z4M9G9CDZYSfIuoEr4xaD0pmN015R64Qa
GWBUsHBn4NYBQMCV7ezqy0JCXRPdYLmBpJOgGYkERPhQhFUgDSczwW+lxhhFvpCCWLovilo3CwVw
XofQbYYIiP5d3YE3Dv1Kq5AWZ+Uwsi5x9VGVq/Wv6GACyowNbKwvMD+evSqAXZE4Ob2Z+QWuAdPi
9UK3YnuJ4HwRn/UwjTkKhTcpP+AQ+58JU6mkMK8lFEVBrvUiqk+cTHgmNY87JR7dQbydUSGHtqAy
zhHMIc+4LBOgPxv0BKgGO9FMYVrZGrRusb9lC26IwwsqXBSHU0EmZMKjUXT/q5ps0woXA5sVRC80
SVjqPl+SWaHzSeNYNqzERs+vM7ax2g4j96oif970EybxhN/u17pNTqhU75iwfXjE+1P0rc5UkCzp
B3+QYLwjr0QADHuoEp/yV29PLrWGEWnTIlgKJUfwl6l87L34WoaRv8tPjiMS641sM2GyK34q6JgU
20+T0kNZnTfPtspuWtcVDA5xLsRqo6UaHBXTZ+yiBwBljviyz5FxszBM8HCCfaIIt0EgwQ27jJap
2VOLsRI7ufRC5W135U8tFHoWYO9j9ObNe9qu/kNAe8n8HPJwz8kPe4Uw9jlJ0GHGk8Wzbi3DUbA1
5dcLEeVVdr3MhKnHYJ7rJUyBYNb4d+v+oU23wK9+1JR1CcAPf6+r/TEtiL+VcCIBJZd2ZLa8UEVE
2Hu4sSPHBro/fxusYQDakwRtLCEtjemSUyirHBZh7F8mY1U4Z7XQOnwNQrz0HKA8oljLk6EDDdqV
ZV9y3s6fawWHbPQrKwNA3L35mKsrHj0OeVobUwN8JKPIR6fuOWHy53FrqavCeUwU/aaJMz2+T1jN
/mxj6/VNq4TPxk1kKNvYrGd2qjm5h1u+FIDwZSqE8f9Gdj/DLwE1+ycCpQ3L2r+S2Lhwx5sPtCwv
jRcpwJruaVn371YzMyxbvuYlRiNRFUWEabWi/mtAAy9OCFS4DsV/kdycp9c3yDfS2ZPl79JCj1BM
LUv6w8Gi0TS50wDLbLEMpM+dcVUcqkbAV98cG/gVSnPkusuSGHteFXqg8hiE5KZMP/JStH9FhQzj
3ei1Y/icx23W9IgtBFRZpx4hB7r7YqE/jNqCcUa2yVxyLxx855TVF8ZLbGorrTe8eKFW2Q9VUn1P
yFTKCgaozZ2gPD/UQ1l+CIlWi4QPNDLQs3BjEFebdwAkXeQLFSa/RvvI4DrZ+6qq+kp7QPP/zFCX
HIXMJ+M79Hh4+PGrqIe5PTxCPSR5T+Xr8yesUPdwC8/TY01RZOs1AL4oXeejPmp5msXjbC2ba+kT
LDL9jpQktjQ/nNIIKiQ33lu6k6yk5uIlJ49ISznhiCq8K0wikBCUvKhcD6iEMqOsnMRrKIOaPz6B
Ww2ic6zZMsYcbhQM6b3poB2ys2JdvNwRgK9VmtCpmAVZxFxHt014nvu9uiI1LGMrhqcGJXribyS8
VMT7bzjaOWzwgRkSKbiapCKXlKcl3B16EGl9xvPMXwwDSlfsMvKEjJ9gg0HTOamBaOMWc//GoSbN
CDbu/PXOe3knqXcsIVEIWzydZi012H5Q+ZR7mnQlBMlmahgzEqHcJ84KVu/ooIMSadwK1v39PuLk
/A63x+l5d0dg6TFJGBGallx6/BPcSRwlAMG6OuDDdb3sLpDiWolNi2vM3fUaWZw7lZX6R+qxBnkV
oa4/DKQirkKXnS2EtjNQPYs/n0fI1G+zxU+WLhSec4gu407+H3ybPx53jq3OiQZDr+XmOVnex2u+
6LB7gZBdHLeyt6TN0HNlGumCJ/G5yt82zmvctpH80C8aC5abJBk41wWHQPVKFEjWJE+0g3YVm6c8
zSE/Yp3PapyGjzWRwDZWTsPp23RR6oaJEIHdV/fH8FAtnN04AIgVvcmPS+NsEU0EEgvnipWkxwcV
jNePMhalkLR6fcnAuPAX2Pi+0T0pzpgp1TttGmvLU1Hi5/dcfKg70yliZFZzNnXC1CWXU4Mu4W/j
ZnQ3yYKwiTIPdDAPrEu/lm1c4KKAPgN+Ho7U5+PjvamNzl/zfDe5UTaXwHaGETzkOrAPNwcP5cPt
k5dpwOu8tiqxMAAYvLDs1mRc7aivrsBdbFDEfrzqSLBC0fr3+O9uQ2MpGVkK6M5eG7CVolaZSd5d
t4hj0MctVsMLkxXkDbNykZgu+i8KXFfJlR3pO0/DdcLid4M22LJ6rpSlW/F7MsDl4ZmFMwWQbrtQ
SI5cMUbJXktMjqObJadvY75zva3MuI85FQYImYJFbsDPhiLRXsTqiOdywhiEeR8CVdihAnFcd84y
UaS6VxZVc23Z4nFoZkj/95w4ScFzxJtAAOQBgIAOgCs30J82SqfZ18uWht8H148O+hM3liEsAhHm
AauvFJ8fQcEGMryOW0swgBW6Kec6TwquqMdH69F/jI4JX/ck2rZ38b+yNtGRp8jRrgTH2n6ST/7+
Qv2YmuCiQsxsdzwtRu3n4ozQMlj8Ngjo9y/OMfpubrad78roHh8GgQnLGh8us2Mg0HPiXVOF+6vt
ni8eAzpe7NTHms1pggUDrFRkvK8fqNwtOY1Vxfs5cf8Owusc6fWGqHgWurb3nqqfuKA3F1GMrVcU
8+cWp0tac06TCbLTlmeGGOLstDdvZm+3fmWH9RdNq12TABhkwsAVSR4Bn2EnLkqqMVjqFSuSE/W/
anuxy4vFW3iz1hv1FxeQPct1E0wrt8mM8TjVEl/kjPeuxxHEcVBRU1dvH/zXSxngLnQ6/ZOqu9X1
35cscHJaAZd8XXx6d2lzmy9Ul8jKDyRqFpS3AQbZ5WY9XOA2Arc+d0iKLeiHrx3BcXKNiYy6P5VP
8ZLoqYg4lJNWj+N24YaSerDBeuhZ+e1fxDJbHh6O6aOzf0dQZYEuycRkYE8YkOXB8sh87A9DBR4U
6tmDqJHay5aCZgXWMMK/6dOt4buZY9X9wv1+fshNOq9glIhwgFxSvstZ7BOMhK5dv3b0ojIosfT1
5RTT/rLknq9nhEP02/CpZPWUb637jNubbIueE3QEclMjYJeX8x1QKnPqsTDmpB3PlonY0hrPfNvs
t3beHEKvSEjz7xhjb4fbNuLqWFp2QmNpIAyb95Ohhl+JDRnBTzNdi214cOONnWiAtGpUJQb3LzSz
S18PcckOydA23Xu9mXM0wfyBzxIXvyPMVvvTJ11lR0V8oSm63/O3gPSj4Zt5QcF4/4sH5Lel0iSp
QrDXezuk28qOzgzCwaGRjm3yQSBfN3OS4X0lt0DcU3G6WjXyyEiVdNlSu0QLca953XOAFS2wsrbn
J5Q2ccE7vjPpEcHLPMLBg0tH5jMlCcfTh0bXm1u7aNS/lRC5T5xG1CqeVKIBV2KLWg8+IhaJTk0f
80wy+3+boPkb7zd7CW9pWUzR0Wryk5cg3D0UBbyVjM5KvuH4Ojb3ys7EybFdjuk13SFb4SEnIoQ2
yj0RN+unQZC1q9CddErfhFiUFf1L8CIgeHqKzwEiX1jw8f4W/2euFcOlwEXyqfolBt3uxLQ/fu+R
sFCdiWIcp9vqh3BAfyXVKNoUKP5XGYEg+RX2z0+my8G3k1IxbOREMJlfOpCOTqrDlOb6ac3MiEYe
wt4zP0Kws5keBTcrMDOeGcO5zU6G1gG1KrH+NgFFhy6CHbpGumOXMf5z/tosxlPAeVXslKeJJ8XS
ZktdFjPqAyRiIx6hicvdGYWo7IGzEsGoKgfoI/P6M7REItlBnufXqVYnf/K9a/ENXxlsFSoCnCxO
WS6Q+bmTJ6GS7hIqJxMqV0/JT1tU7RATmrcIOdTJK24QIUOzGFTefpS1o1JHPbGTXz5qfNFzo+Rx
fEf587LmaIgCGOvRxM+tSEJPBGpXHRaaRQq5SaZBWGvLm9Tmze5rBaJIa86oFFror8KLKGqBYPSv
rlVPt0ha5ag3a5iUIx274xPjo2ee9/lhOftoHrbSHsYNjXDnJ5Xm0zVrgP7rgR7Fv6NJO6yJK5/v
S7UMhHUi1q76/w7PPUKEfzw69+LFEA5wgzyQV1XGuI/MlaiOMYzO/1fSnQYIL1yVF93WZb+AQoro
Vi6s9K7oaB5qRJVkxd2QM0b+WX8lFUNVqZqpdANILgrSqKs4Yt1oS0KIO7cGgaiOQNRsSP0WR1e4
BIOy3TyQubfoQf8dbtD215fJflyO3l38SKB8LCdnP4rWMkw8ZRoNW/Sodag/MF3Bymg70CmlpOSE
gdkreZEVIEAIqPKwDBi8OW8hoRC0jY+3tIMVkZU3PrFnrgZd8bk6nHghKKMdzW++XCl+3NVX/uZ5
NgAHTfVkIuA5rfFIcEsXpXfRnbEhA8dzrR7UFha/qQfJTmmUkGWgwVmrGU66nS4TwPIMYH1omiTA
rWJes5P3YZ7pm+NnrW6jLoUVtjgRoAJTB47OrYIAHfBhPCC4Jml3ZcTFGpWHDrcWNpLy9geS+8XE
rEk1YRE+cK5oORacMsr1WIdvyjYOvH1lL4w6FQ4aUwIFPAYEyXgG8u+Gpdjxi0efMXUoa6J7eO/N
TPChX9bNI4YVkSuxrAMmrL2RTXGgV2hfLxNYaM8Z0RusXLvGSpAS00tVUxOzW2X0DSM9MJQRq/jB
f5t6QjSKE/KnyKN7Jeefi/qcQU310JkWKFryyU9suKa44O2+SJHjvC/I9Ic2seU4544cIw0FFs5D
iiHtcJq18wHFF7a08XR4hNQJp08QefmOL4QdtuF9prJENx7MTBTUqxLxZFQkIRGri7vjWRQFljAJ
KtDAPiMFDQwzCMK9GGyCFawUVHsQ35bEsjnfmsdZzHobWttSFYYqw2vOfC8jSgJryr9Zie+NQi2R
sXllWK7pxzcAJJHEe56UeWZAqYEw9K94OwoAhn4PZe6QIm8ZYpAsTWLeRCuvZ5dea1ZHK87uN7BK
ugrbpwY7CHLLP/pd29VHlsgoRocNuSA6CuuT4b6NT2eh2Z3QUAL1dtaK69G4VXKpgLSTD/K20LWX
KZCDjaHgso6in/GfdEBsoPoLP9V0QYLmYYTM8+9cfmLNN1XrGk8ytWdBAlZNTZaf3exG6dzBYFXw
0m1aocWjuV+iq5UK6WSMq0vQPCVg7t6CexPmUcMMrZAYzOmtYnL/MIltoQcBf+kr8iwqzSvzPzIY
7Pkw3d7IooTgjkIC4lYnHtEvkGZo8wY62+VaJiGnslRvIK8Cdg5DSqDtH8CEGT5ZrOiM3xoRFHDs
nEgwd4zfbMqMZb6SjufCQkipGZ4pQTWMUWFnh3AcOkbEDOmWEeyVpDVVGMsHglaoQ14bklCfBRw+
qqIywJxd9joMqshB7lArYUKLWZKeI8qamnFY268X6qnIHc+sMq/Lh9p/8olageYkA3M+3eTDY9vW
yqsKb0ITi3pNBNIuT3rYjAYYBbpLSsPCU+FPAW/OY0dhNMvQfhOrGRWGKeC/JmURxd/DiI9D9tjF
IAVJCDBjRE32Jl041Tz1q7uoAgM3qqJKWwjVLr7KoC581xZUJN4fVrsx8pUkLjHR6XzTgXEBOoZz
5ZOmXD+j4p8338ku/d4ohqS2ocuBk7pW3kz4N1aS93XEbBuhtMV3H3Zm0KARXqkJQPpfrRU58AQV
0lXoTl+6OGNlyR2mnlr7FOlsegxgf40ymyehFPwwbnDlFgQTBZbPKj1XMw+aGhkWXsnAOqi2sTHZ
KQePfs2zy7XZJ9vV6lk4MMhmfo7ecFlJcnF+9yFMjW6zn0r44zh1FmF+zw1wHE0ayWvMMm5oP6rE
rzirhZBbe2+mShCjQ47Yf65qmjk5tayKpvDJE1vr0d5XiHFjkl/00vU34wGtQiZ0AYdpS/RUvUuF
y9ZGDFCDnetatCw4OKFSOuTvATarHDgxdyJ0dICQB55zWb4kTBtUMA/Vt72q94RTITcSxpIjCucK
z7PMaLhzqsy/Fc9DJK/nt6D0fdld8w/Fb2PekVvWSseQCM21YVZ4C/iAHQ/OXVUvvN/6kcXufeRq
8CEZvrEVMgJQYATy5h/ZbHRZXKD9cNcAY+1kYYH0gAS/uBoCfMY25a1UKf+MQ9nciVX9yg9YyAVK
T/AUpSjwTjicMjP7fLd4K94VQK0f1y6yWC9xp9R4WQBp3j9PiEOr/tzwLKqV9KFXTRgA+8OM3YV1
KDd+li71/JKRDXE7WxMF6zYbl3UOJFapzYgN2oGK2HHfWi/iPju473hEUPQCFmhwxRegrvSeMKQA
eFE3h8Oy8oo9AJ3DZdFmIXtmJEtNTdKwr55z53s8+N69dIx+Ymkt12A3vp/05CE8RAqXR1qNpL+X
9KondD9/ok2QSJZ3GsPp28oLKEszQQ96J2PHw+m1VpTU2nnTFlT2vW6OxnF3asWB0kMDs8WJT3KY
KIzNn2H+4G/R6UvFCBd31MmUyleULQrpUADt0Ppmr5uH9Pa9BVul9FTfSoCz7SieLQc3OZ9jxgUa
j7xoANihF6xWBRDDnO7E0kOJQrkfSnd1d/73R6kEJTgCTPfv1g0cqdDSIEvoX1RBzxIoQ9ok1lod
C+016l6G5F+NXWT/EiQD4Bku9XzJ8EMkf6XVbWROPRQmc0enIVkgFPGV2X9qiaZvZDKVMgShcOJ1
OkLfilsI+CPBcD7XoR5QRiTuC1vvRsgbFL5fc4sez2SnvkOtM9rsEQtt5cPy3jAszq3mUBlCd6mz
7dJ7CtMT150plrHNLeaDIYhiaj4Jz+t5eU0DInsZ/Wa4sfz7Qjqzdw5gcKp6LIn0YFPqm6fLfuRd
fCu4bhkgDU4QOPOOFWrSZukXPWu+mETod9J1hAIDZIFo4T6Bz2YR0DYyOgBZcbuuUdb85iGP/iF8
XulgVO604BiIbtqzdjhwHlglbF1yp4G/mtCslAMKO6ibsmRYXBZUlEGvqem4H2Lx6HnzvqdB+tkB
d7Do2pOtdQljHfDKBBI3UYlfIxyv6PTCvLnndu0rSS7DsZXUZFSpXFZ3fmBhE9F2k829yQCUpGLd
7dcGsBFQ0zZUY6N87+FCkTVU2GI4Clc5d2k/smWbQVu2sR7dztdzvPdTu7cqsF/6yhhhhBMWVK4H
PJ88+DCvEiFsYl2UnRZuIKhQ7bXGWbvfr3Adoen2NFMqTPaHIKb8Pb7pR2vSSCz+k8VianlDXROr
vJUt/kudIgfwJaJ7tnuqHexELakmkEByVEnQVMKiTYS3Rf1yYlm7xPXTIoulxVrQGqn7YFSnHTNU
oTciBm+qhbIZMiMSCPaIfrC1nwrHXDpbNEZcTxfCuDrRiEybjwJ9u4Fv+7128E14YzArGB1GpFok
bdNaR5AV+DtAOR9VLwqB8LiPcxagoa6mh21bSg+LtL1ZeXYphCO6mL/Trv0zCoURa8pk3yHavYJK
f2dhQoEuJ7KVhjv4w2uImLiDfiWfCja2IqCj2xSXDQVHrhl7f7yU60PgBbhiw9b33pN0XUngYzmb
kPCWK8ZiRrbpyETLQo3Z4ih/GKlS3KCW8ORps1Y72w7nMZfhtX4Lj/R/+WeTTXtM5+GAJEqhYGjG
V1VfUmBWsgf5BS51Pn9ipoB+PQqopa1oL5OjNHK0w7hiibG8AaKZera3Qm7AT4i3kHGgqeZs5Ueq
CIfI32lNNq4MCX2BVn9e4j3sfq+xi5rbgTn1E2+U317gy99GcNlbh0aBWAp+e0Z02L2abjY6RMTN
/2G+gta/yfPM0ufXIWbCenPojDGV47LgyrFgjxVtUQJz+9hYCz/rJixXSkfqL+4I7MXIv/xfEMrn
b3s0Qt84gkASgFXgvEmpCyX/H/bNbYk7Jn8N55VCQ8iP9DX3DufLW9w+cEHZnVXR5+VZES1XKDN2
leZqmBc3fBn309PvCyqioF09y4WzEBMe5pSKuTobH9DXh7UWS8FgwTyRZ4leXSs8GWQoHyEckwrD
usUpQFo50Aae7eAeUdcM4DozAiynmSM3Bm+7oeQaO4oIbnBCRoZPcMbLYkiitWcsfU7RREXr75yQ
9cbTtRhYPlI5RsxFsQFFq34l8R8LVRVPNVWt5SceRBARnS338bydenivZRpJoBB6iLfLahUn7Kyk
Y/fAPbKp7vhDzoeFZ6mklKhH2rBXjRsxCsjXP80NEA5y6dmS3KyteYapvBh0YPgcXh3fBmARSruR
lAoTmywiMYdaiThILF9pd21TJq7EANCwBGooO9dE0dy+YUxp9Tstvhw7fCvJure/JEOCuIKr74d8
ZkFbYnbcyNBIcaWnKhMyCFkjDRVyQ2m2oiuz5WX062c3V3ASI5grhA7eZFDdSuAAuMt66BWLWYZ0
rlYZqYhstvvb8Ojwf8OBeJpQDNDiWogIAlL3ntEekKRjFg1bYOc/sLJhh+gHSFVg1OhLY3juye1I
huTjWxWnpa6UG6w2h8C0YmL97IapkxLQfSmHkzIhlSg+63V51xAJmbzeSOBx4Tro7Mdi7wyfh4Bp
zZFYeOyAZMihNaYdaVdOjn11CdA8t7Js47xQpKK3/gQdwuZi1OvMrWizCdxBoQarNrQ/RvUnHk7A
jiB28d1idWciMZLGv6xfG95NlKbz4+mrfWMi4Vw4bo09eBt9g38fdhWqQBenFuhHuHf2WQVIkpqz
cAMXT7NnuDCBuHWhUL+vdUj3/fOKX1NrwbQ/B0a84V/FmhIx0nFBQgcaeVMiMUNhXoKoj13yRZHR
zEIKfPQsZvJepwr3tjVwhAu8i5xoWXrK4E5h+qiaVDI2QIini35XPb86iU9QUG7x2ObfmlNjsy8I
I2VMhT8x8VpqvVgbyrJq59Ly5woLP++VJp6i9QX8dp0cNUU8aW+3mx2P65dITUxUa6d3kqVQairG
pOktSHaYKd6oJpvi5U4/axgxofuE8OO6FjYR3VjQMJ7nethubxt9Rf6v5sl7jpdA73d8rBx7Pymt
jsmUwm3SZqzNKO2hIG8xt/xAGViiXNZjePskye4obIXpSCsLnJ+9HOu2YobkTQX5ubgswDO9Q4Sj
Bc4R3hQITSGYxNVVJo9Ld1/1vVvb7xTXcWUcwqgEh5LWkl7BxEUBu75AJLIX0uI+x7SPLNze8H8h
O30oeSV2fGJX9k3vwG3ahL/0e8NNrIKmQ0Gx5KatuFm6XUwMI2PSOiCGqS/oXhFlHQoJLqp5Wn4t
vA2SmwGI7sDDTSqeqC0B8dR4GLFT8rITlVGxW+JR5LhxpUFXFuVzaRCkFs32z/CdOfjjFfOjYpbB
UoWnGWT5c2o/kew49LR0SLu9Csv3oUkpR/panfKlOHYFFnN+1HHORftPL/DaqeWFGYCTUf77LFah
DV8P3HRjATlE2aRAm29t/eKNZC2sgYCsdyxV1/sesJqrnyDpgwxQ5wQY++MyYZeEjq8Qpp1L6S+z
KoeQxhGaoRfTTQ0abwcmU26BdLVy8IzPpZ86ZbSBTmmwMmGedeVo3hvfatglFgah5vSLVrHIA3ec
7apy/x3LNBgSg0OOdObJSNUHOOVtc/Jhb5rUfH8gaVr5Gv6UtUFrHlLOnqc4Gh2X8hMTNyWzlFGR
X7idU33cxnV8idq0XTo8KP817m9b7VBluNILuo9eF3PWr0v1VJsEY8aSnLkaYgwWqCUiY47y1bi/
tWeBvcZTBL6ATWu40BCwaM/7mok8CYLmi0zaLjnKdiFMUi9FZRGT8Q+nUNNyIk8vUDkB4EoP0zOL
2WweP3l8WlmQjCfvopjwD2JStPEu/APSiLe6lMr/1Um7o3iihSKHcMAeRKRc7MgTNAMGbNJ3TxV+
QKKsYhDDHWdcQZUrRQ+tmMYZOuhROj9o9aGbDlJ69Nv9TCtktBck8BxbKVGT6YbNgYD551S1v+4m
RZ1y2X/g9AqqBGFJF2cV2aYyNwsKKq6Nh194gzTDBAqHJDUM+/fJeESSdtYCXWauZy8IxiryLcFl
O3HXQq/cq7s7mIjGgscovYJngEDZ7uYSM+qxP14YVB3aOzPvjhMtG8JluVGJwRvK/AodFuhZPghX
rv307OLx78mXcYcTYZQ+hT+618UsT1Raal9j/O08Z0r9WowPkA8lbMg/TrZgFMk4614GEEWhY7d+
KEg/jDVO0qt61w+TSXrlpCWfgPIh6urs3oUZ5DR619pFmWL+zl1pN/duXdlB/fbeAIoZCTqi/67j
zSJs4OKKKx9ZowJpEa9LlK4pUxr3LQ56Juy7TG3FHgZ+ssFXl6K0My2fLFCEEsfik+mx2UYZSLxx
uLkeC9dbEkHrX3RKZ1Zjenmy58KO0F/XgHblVRgQXs0cmpZ8ER45oYi4Poa4Wzr9LXFJA4EEj14s
Qu1JOYuL2Pu42bi0bo5kY4Zg5/uCN3cP7unjeaogUb/Bk1+LY0NN8SNT8Ci5a2Zk2VQjbLuaSWI8
SL7Ns/kH56rNKwC+fo2sD0/2nvqIFCBKsky0FGvKJ7EGNnoFoVHOyzsBUUWsoUlNQUKr4tpsETDd
PjoQlFg4FA5myw3F91PXqh7N4qDPk2Cp+M8QNdmYeY99oICh7vHHstwl4aMpG+NZXX68NtWSEk5F
n0ZjAWvAXqWUtShXIAVMR4Eb6704x9g67JZ4UiLcUdpRNj5ZlQgh+YZJZG+l4jIESF/DtpV6/pvW
WRmNHi3DaBxck5v9xo8cpLjj1m9HX2+yNtgKICwasc+xEf0pXHePThG5gc5wAPbmHE4d4J0/gq/C
z7XaIndAoieQPLh1Ab/PJ7uighfZnpdEtl1OOXTtD9oAWkDBK3XUU4P3B8RAWGE0pT6iU29ZihuY
FhnXtbtFSTZB5iX5d7mc8PZ4JN2x+6Ag1yL994hsowNfziyMTielqOnFWqgoDnzC7ccXJ73n3Xev
ihzflI5RjIx6kqMAocUya6wMbrx458VIJi1F86Ycp6RQPBnFCU646i/uV/yyVipIdIXPOaoRuDJX
UMZvfZnou1MaQaWRozF0gR8GahlSYAoOvSLzJSo9efhpdf76+s8s0Fi4vIQJ1lAiJpDbJ3viyFvq
yBDKSdTFGvLDpjLnnZbiTdnuYvpFGJ2WO9o6YcwA5Ia149N9zMXbi5Vl53dbkx/WzafmmKH4GWO6
wBQ34NPU9P/wjGNaC8fgt/yhdlWpgFqo3uyVzlZYlb8EE+IRoFLPbAGrq0O873EFaDRygJ+BcHjb
q5fmdMGFfFof8nAYcwSzxqitvIauh7fXKkMtdTAnxZkA6oODQivLEWcC/f9/xSfi111FGy1E+xhd
Kj94tLX1RsYllsjMBKn9r/5OLE8SU6NQtjz/B9VpxljhR3bJzHxtycpT4NU1c3LK0iwjYG/NdSIK
bT+XqHMSfQtv5PUp6BjwkCfpnP+17BNRyc4nshXePdZ1SeQXwyEMuFyLwxSoU1p49R3NWYWyM3FI
GUeZQ7VRVJotobr9SH/7utQcAAj/bEaBnIjM00cDgL8ZRk4K1YBUuPkcSzJIPiPVRfGXenKtpNIZ
hhSO4SE4RYU3khddjDUEQKbKjbDkT33VqayYMAdPMiYPNcUxLqWpjAQyqphnAOHghf4Juu2gsDpy
fOuHSRqHA8T9UcZu1Cnio/cmIOCtdib75LI6IcTQeKa27fWuBQ6DAtWKK6+Me8EmcUflXRrLMuxl
SjPS3Dp+sVLp0s1z+h2KhT193tH+oXC/yFSeIfonfw2vyswXr1yzwUD9yAoQ0SJdwtgac+a+/M+a
0ST3V5tmQIruYBvffHTM0Pi8s/RAaBpt6PB12Eo9zRCaMhnfg7OLgKm/RSoXZWbFgeHfMvt57nnK
igET2qr1AkJKzfvDoSS6ZGBVw1dlV35Gn4LcFzzJThjIkCBJrBW3iSIRToqkNF69AfvQFFtBceu7
WxfSixEeLXuA6C3LGHYhykbITogsYGG8CUmDio9o7QW6PCFI1QK5Hsh1HF6/JiJ8u6Tw9AfZgsVH
esOIBP3L94oUZDC+g27U9bmzFsP6fK1XNhb/+6w5qNgZVqnst96JRKrKBoRx8hafwamq/mq/dOzn
U5w9Z/gzB9PSaR+bWapPHzXHEGRWAve5qQ859Er18uDyRQnSmyFFzT8KOoUF3+4IDASwGNnwroNi
btR4vhisRMGDnijlTX2Pb3NoYGsIkTK98GjvOnHJsUb5kJU4TiDtDy5pLY7UTyT1CC5ojmyAJYAH
tLMI/rb+RwCPwSjOsJelorNw4H06KYgHp4j8dpFaGKMtMTeYnxOzQ1fIvXD548uYIsnPt2Nw9a5q
qgXzh6/C1xJpQYqzIVKz+VxAN1muC+a4tkvq212LHQEcGojKvfiQe3jnmkvzVD7SavZeduAeYoCG
UDsS4vx0anIunxahv740VqzFv5ye5rLs5kNA4eyDHvHNnskbS3rImRjI4a1YtsOf9SewYfSuP3Su
WYB2oronL2D/P/jekHigcOkqc/CWrFgu0I/nBI6KbrHmL5jWF0/tEv+l67FeLIy0yO1jgWNt2mfN
R2h/Kfgi22zs7NaNdZ8Sl61c6rdmT1NP6ciYzEhHMGU+2oaFt+q/JAZ0+F2amhgxafk20Q1/2YLf
103nwsH56NetGjcvYbx0Mn2jyGdBVhIDyi+IPH/FuSF95EPyPCc9exmPLYcPcWZsXyIgquQcjqqe
J5cj1DPPkyD4ZCzgNO44jc0kOKBZ6Q+h4F0OQBAulPoD5vnHS+NSs0IrPxRA4UzDBjuf02TN96iw
AhmMc2atTNuVjh32GC4exgcw7ey/NG+VC1snCEkrOdV6mxhLhY46RdgMQEXgvYYEZuCFX5WHVHGT
OYJOau3NNSFP/TuhwMhOGffiyH5gNdRvotcmohf3tkYT6LvKeVA7ukvIhAZ/1i+41P7vr9oR83ws
DdsOylu9XP/z3ef1gTCGTV3dcjm/G/0O97nIj5QYl3ya4cgQw2RUOwmIMPaJuhdv89sHBDl2pzHn
4pnU7zULRm4Z6OeEWPuCYzILvrn8MV9hIVbU+/yWX5ujoyJkS1sUzUwwkTuMAaPtA920jZqvN0LJ
YQgoAHwxVjkSjy7QCoF7buYrDi1psJJy0On5PZ0iT+SD4HNxG9SkkhZM0sfy8kEvpuxH3NemGeU+
emudfWWWEtJ9hrtS8ASvFbzNh8+ek7qN/Kv+1PZWlWeUsbUW4payeZwjnkk4I11fWHaOxx/B8Dyx
0uforHL8claqpGVwHSzSP6/d2E8IoMFWdcGqePgx0hMHoE9MANBa7fuT6ASW3f5gfeLgHy4M1qzm
Pqgc8RbtGRhFhBZO8hwE61HrAgHpxB4Tiuy0ehnfeqd+rD3aa4PGRZ3h22i4pzKijoiJtRZxwKxJ
C2DZVv0vMwm7SedD94tQBqs5YIL0G7CoPYzouCd8UmbfEdc4stJ1WSiLAV8ox3MrcJ1x1K4XdrBC
qmjw/i8B49J2Phie6G3WulwjslUDO6WBZcTw1V/yiFU5Es+UU/XbkMioSGvgHmGS+wNPPzVvtgmv
YVFby6UUVOcDk0cOZgkQzyaPl5FYPE+TjTNXD2lUBWbxz8q4NeHPp0lV4Efx/xXlo7rYvTDsd5wE
WHbDqc+L89UVimrb6XYg4LGlJr70rhc2DLgGVEg3QIi7cWK8Lb7P6WgtTE75Z7Wutc4bwX5Mbyl1
zkWPmcgnIjMiHSt42HMr7bwivZiSKJOKcQ7/4EfoqECDXGn/0XPCkfmPU43NH57lsuuwQVdOeZyd
GDXL2WGKSAaA+zqNFFH+vX90tn2YDanvLit0IlZ2wEOPMqhNyorkyGkJljozV96JKNFqcOFXImhF
CNkpvGR52axFlQ9VP+7W0yIiiwlXBPe/0BdUBgT2bfmM5CzvMFtYvE0RhFgNJOWZJBC7iN6Rj4Z5
lKbOCOK27pxmTya7KMqTrnBgF3Hk27MWw8je5W8Ox9QDPXrcjlO4QZLHrPL7uuUeoSx1YAZ161XK
EdqB5nEZdLXtPxhPZX70yqkYzcNS3wfcnrnl6KWan7Jqu5du2ddrNs6m1pb28FqF4HFtz6D9lZ2/
vHbzc6qYRPA5OKD6jMBx41rU6BmVUaE9vlH39o0TMvfwmWiL+N9kK0iErIp3wZyat0qquCqL3nzq
DlF7n5ZfYVJ4OBXaNpGkO0gXDimlPItf+AtwWXA5zuinJB9cB4+tTYVQvUNPlSE9nCN21x1k4wMn
gh9tfsWYGZqFfbOvpGVXdEqHQV0gjqr7+xTaNmCg509rOktrCHP837QfIfdW0xprEONg7H4QqS95
aZw9tU1unbokFIIhKWghkAdS863hcqX+mHPGJ6oUX0faYo8vbdbDSCY6opH3x6DnCZb7P4oycmkx
4rv80OyYSEZpHaIyAXXhl2JV3AIsP+zNB9BgSLYdI6gnNgeE2UYmsPJNRDX5DNoY7errAPHT3dkf
8S1DMiVFuihSyUvFI/bqyzeTq1Ar5jmbgnvGlqtk13obGbokdUCYm1QtTKxAK3+jkO65ZP8w2Mw+
KlN8pljNym5KtuFQFpXvEhYrbDcWfRIQrvhG4qqJYkiIIqGSR+NRs0FNPCcG95JBVU61Bh1pJci1
75jnL2P9MbxBhYWXOg6+RaXMu+j0FMlJ5Db1LAoeem0CNjboGPob0P2mAE1nwh9kQq/M84AHBR1T
PvtRi/up5t1yk/rBVGMYLZjpSFurO1aSsk+np0r6zPl/8D/m5O2DqImLX1BXCFYicnaKiGYQOBZt
XOWq0IX/YviJnDFGB/45BGnWCL8KtT8HaFMf6yO6Nx7do/jY4QfzQkKeaMXPl0+zVNqGaSRB4E+V
j7cC16gRSuV4R6EtU1v9p+3iuf/yOBzMcgEvzhyghItMaT0SBCXqG3AlE/VXWAzOqvQsqt0jJzQN
9hHt5m2z3aHZ7/68QwmQLGL2FmqI69Yss6J6eh30Lcg1qYoLY90OzP0PnxRQz3qkTgEabkY2+bTm
cECIKjUUeGW6pJ70a4zE9R9rq01nsMaEctv0Ddetibf8koWHRcDV32YlokkzCzlih78IN7+pUt0/
hIK3Ot34BRi1L416LcmW+VoSn8HFXcCkYuBabfCXlsB0qNCE8Yj7w2rYG9Bjsw14TdAmHbZldaW5
ySecckVY7HCDohrToIDdaYduFP3hPdXFcnzjz05eeZcR5KHDvcKKFWrTuhJpq9sXI3EYv166XQBf
mOqCaYWWOSzUPA1Za695SRMgEN8MpyL7UHziN76JDerDdfVhn0+G2EL/7R1y6KTi5SOBch3V2LaD
X6uoG3PoeNvb6hLIfo5xYlIPnzp5/ffJ6uu/MWpBY9jCFTEZrMsefJs8ca4RTkM3u8HtNaThQ1Hw
9lwCltqrv92B/cuVNTpfbSMdyEdDCU5jVRBzHTz3yGjWjZ4hxOxJ75D29hPpVO+duFmCsTTSGScD
GyHZqt8XrZ1N8M7Z6ftuEGS50XOb7KprVaQy4LazNOcl/io3Vgwp6wGCohZ4u6y+odLZfQC5p9uy
TSzmnKB9Ap6oPS22UWcc2HnF0tNxEJyHKKEXKiLX1v7OTUjSm6EcG5iJ/v+5/gkIxTqyl/HXuzt+
QFC5cZm7FFKS9PzYatmfGsdejKLicV2IzEwjqlAZxDbqnPmwL+Rd/IgagovV4i8OJ+/rJ6acvzwR
01/0/cd9b8UZQcDD0OJkimVw8cqT9wov07o8A8b6V2sDqjWBfjBLWd83iClAxoclt2Fn3BtDyM7e
LwsskOiZdtW+pZBDJx/askgtwbHN95gEOmi/b0LSRGcVv2heRBw91BCJgUr9RrmgR5MwPehYital
o/PUV7ckp+lyrt8Se/dv+b4Qht8GMwFMDtUaBW1OOKehnwsJCZT8hjI/AWTYwVYKxEGkoZcZ0sPx
kqBDVtJhH8xEBUOysR1nO9Av3sOWTt4/zfUUoAeAjPQw48006NNm59KC4n9P2k5MvTHtIo3n32fh
m7nGiKgXL/KdrY+xluiqvwCN5Ux6i+cvEpVj75OcQoQrRrAD9drZHr/0VlhFdXPiUAX9GJF3f6k3
wAJPAEtSuIxssd/ZuSlQXUqtqRjM+gsdHjLeTYIwsEZ5WKV4wASuN8ZXTEkGFzSpTrhP05NszcM1
Zxik52G8/JH7FtD41jyXHt1TesFs4lNcKaoFLGZNRb92SYzoP3w2o9Z9fEQ02M2+x9PazR4PTF5a
s98qTyidQqQ97/n8QfTNgdnr4Wy/zJZiW7NNCC+0kBvIFtvJQT5yDr9xZvWXPo4X5fr4+MSWEY/8
UvFBtlK/uvBULJXvKdo5fLPMbtonrACXqYSQkOsf9/V5n8yY9AKw/xodba1THUoDUvNzeWpvp7L6
TktqbsBdFXCNCykmJ07WiFftc4a/YyS8bb0xHUv0FqVLvmfRThJKkNEYfNzd6jy8bkk0S9HFA2Ds
LI6hRPUQPBwKNrSVUTnhT1+uppmeSbh1GmIZvApUhrMBLoRC+Ak6bBUcDNxp104DotfSLBrfPDhy
jTecXXfqqhaHs02yaofXrXNaInggwj0+LqS++8h6Ga0BtQ1qnY0amMlCvKeuuw6JKJqF48ejiA85
qSue2yRRw1UbbKqAu08TfdpmGxOHlYLXMKwtI24YGD3kPPP2+iiOBa+STM4r5Z7v60uA9kbdfn83
umJjwbNUABf/6qXkx2uKO3aHrRIcH7/LdJX5usmkBIw/Wz3cXaLXGvHV07kP8uPcd0LH5GR9EJik
Txuxg7VGF9GzY0sw3R/XZNKp53mcpxJk3v+6T4IQlh7rmF86wU8pBy3G6xX8UoJCC4Fjr3kRY5cW
SfG8/go46Tkdj4dvrCPjkcLGpR0Q6jDVFw7v1erEulyLAEl0LChlEtA5cnYI+FsWeIKmEb3tIbMN
VyYdWMeTNacBtWvcxLv8WIc59kBcpj9+gHxGzlUb55mrx0N6Flhcet7TGxFUKuaeKiyp6/n7830g
4Vsa+vWgJ8xC0qNk8jaff4hSsTd9SAJdCP8m7zFTq0HGbmSnTIL/go4mJz/z2bQ42lTE6drS1440
M2t3yziMiiTv5aMuYtalrhvN+cnIH4x10gtE11lNn1/fU7EKu9eOPPhddwAhibduQvcv7h4P9IYR
F8X3Gw1E7pwQk/wT809zjUqvf7/1I8Gy7IzE/q59Ras46Wiy5D4+zD7+FWmMfX7hn8EL5Q92wQpr
4RmbHJA7kyGiyx7khetfpdYVq3ZPoEQcoue6avgo16N3st62qDEcT3Y8p3+DaEzK1Z76A2jtNmRp
wiNXAtig47hchZ2ZvJhPzuR6/niB3MOWvY4DcD9h+xCLYk1Ur9TQXXGGyyKcaoudJ1N9RDYdrH4a
MTyRpjag3zMOCaZlBa9TI+T4Ca3WDBmKsp6nJJRRvaDhzWCdnIvnHjo20m+5OFBUJ+cxj1F3/3jt
2QbJ10mVZHVGP6U89730i58fTUhs5Mgk+HwOnG9scun5n6h9oq6GGM9lTOTKPbeCR3f63NfW0CZw
TqVRmyatFhnCgSlMq0AZJ9vQLabQFaw/9Q7nRoaVYdiG+1K0U/OHReuEsuTI97m8Zq7grlc0JjSQ
19Yycnm54SqOz1mkigmyG1Ne3aBfWgGyJKkfpUsyg1ieHqbmEHbGzp/O+y0w6TWSufMDFPMGZhPj
GIifel3KXR1/PIeQEjR9LfDxsBUxxKER4wLEwcZEMbp5+vvVeMq7BhmvT4IUVXF9baq43J3KyMlf
+TjcwIT+TRU3VYb5zRJRYvg9NKERlHjSSnsojPOvXZxrmlZ17FI8Mtg6UuyR3i5a2/THnyYPw5gb
UkTH8SS7jWHYES0g6P7glhprHXZd7xBZ5aYZrR9RZ7f+5Uka4mx3Mc6TGdMMV1sZOdojJr81t8pE
HwaNkxE9IWbz/d6yzMoluYxI6QGSK5449lvgcL42l/qDLWCNLuE7C/22DMHPd/0tFuTbcxdn+g+k
EDZDGgV8WqXhSWxDGvDPpUp1j7rSs9CHQO3WrbcPenEAfy9MioW8/iFW28zShz7UI0tquUpzcjcc
SzatpKcjxh10VpnCo6aDWuAJMf8MihDPdZtvxx0yAia/LPgJluez/QEmOl8kvHXiPWmsRKuHJgCu
bAHoQy2yBJNVuti1iMBHK9+/autJxgoHCCjunrgQHAPEEESPvWf5cRKQv5p0K7AEhwsZKG/mS1gz
Npx9V8ovlnsLrPHisZ5MrJa6dHJf/IpwbdHAnlCFvBLlUNpm90jBhZ7Z3Cq3vwFfalIswzIQfnw3
D15ByAzCYbCMbn3za/mVcSKRdP45GFMNw4k6PKfXgYpufljx36vkdl1qVp7gUj3UH1hiaFk1KI8U
kZtIFLkAp1WKRngRHGN07s2wera4WFIbSM1YUhu1dNYEHft2j7iFphCLnTWFu4yqcqguOWpGr0WK
N8k2SGFqxTKSe1wVd6QB1Jy88X4PsjULH0va+Q6sSjIKSq4LzJ6ad4vPCOkE1364IxL70UvGhco0
bwHFI31hgL6w6YdW43+US8xALgi8FwxtqsclM1EpqQTUF38zXZUQSAkekUpy0JFr4eBejyw8EIFG
iv58RUQ4MriZkmkq3Sn+47s+jDdRxssN93zyb9rsCp5md8cYgm5crGqj690s5U87uNH11KH5Xypk
dlcuX1lppMux+IcPsZvBSz00VrRgH/zOOWWVJZW2Dcju3bDP4QFI7A+e70y1C9+ExjVP6C/8inJ1
YYmSfBXliNE5gQagUqOSb3SoBVqIPPT3IfrZC/QZG85nH7iLVZC6ycBlhp/uz5IytW33PVUu6Cfa
Nlz1QC2k7p74xbUxp9Zc5wnFaSP2ofBKYKYoQr2kNZP+ErLMZDD8OiiaZ5gbSJJJUcZ36616kMIX
mEj2rf6I1fsfTRkQwLi5lLxGGptVNwYosfWo9A777u91CJVaZlL2BHCAhWWD7n6QhJl1f6IXKFr2
qZdujyN/dCZeXpdz9evCOEyv2g3kXKohZIstiCe/RG57TLfvKXpjQGt0jY9rrAnKuDU7f4uYxyqL
G8XjJ0pVNytPg0IEFhJphg0tJ74H8AJB2L+ItVQN6GFJjTLzmFxRYUcjv7tvfiFtA0d4pWZL14Ot
KdmNORWSrs4qkX7sRUulxqgW7MdbbVAbvKXF6WPKRLsHJg0QmzTbRKXdi6W1E6bAxBErGTRoxXgA
XwHZ7do3y77rmHO5kJ6W1e5RHoJC6Daz1ck74KHtb8jHu4uSMW7vDq5lOLInGLnuFBYaVo9CAymD
2xBBVNxQUuABRk2BOcnBM53iQnOgf8vaIgPSejRtdJB+O3g1iCyoYAR7iw7I40ucWLhzOdGu8yvI
6Lh+A66OEOIuR6HIYPJtdVvU7MrZQYqyPNu5S2f5JAPTU4hqkwHVBAc7ilN66LgbTGMAiwwpo5ja
7e2SSfF5bajolept/E4RKiBsiSO4/vj5b2Gn2SYAnocsp/Bu3fQouHN/AVaL76f/pzW+arKtwd6f
FiK4g9fmohBGMFE6n4dbX/GFJ8MVVftVcw1JuAanKCGGT1HhJkoKZt8cQrkTmrYtXR8/48wem8zh
yCWLRmAU/SPWqzEvWk3FT7VXm7OAuxkpmTRhNW7CkEOL7z/TsV1CHN1+yGuBD2CmVdfrcmg0oksm
WgakWVeo5//tMtilmNKGzg0uGydVUtBJabiw7MOoEAygRk9fOKtidG8Xtx1JlZQzifyT4Ssoerdq
5iOvZJQep8wXy30kmqz24uk5GluqkuEwZRYneOPjIghmT+/KCyg3j5JbulOUQ15B7TMZN9Tz3uGg
7dI5x1aMCabwcLI6lS4a8cyz3cUiom8F92Pglz3I75yti2VDiP15jwcdCPhaPV+5J7aE7gBMCll/
FTd2CWh+e3IljoJwRTPK2kolazkhPMuNuvu4YiN+e8ekqR0XhXFoJtVz/kHT6cvsY7QPYX4ke2FW
zOExiKyLuiSnKu/KaIpo+48Sctg13YpfHO6OL35Y7kvkGTdUKkQE6HY6ny3aeLBhMnoVlLM1r7+t
dj3dtqU3lCUPa8rB8zcDZsqCgAHiQJrl3pms43kpFqrYfGr94iOplycj+XykJPqixl6QNUjYM84H
4vNjH1HjOTwzHZh61EEZwDQ/QwZ+PvGEq+iRFz4BwKwSyH2j+ev6bDq9gtVu9+KxM18nSn6fE9Sk
LDhg5JCDfLE4oO/IrqkJE4gpDb32HzvO1gV6Oo4iU1iKM/V6C4ygPNdYb8qMFQfzR27PjJJfmUnz
EiFxPW33g2XPCtQQYWCu3BB6esNLc6Z8RCTkkXyiDOD7pq14oBm7NFu5GzIjL/n6X8/NuEb8a6Ht
0AO0LzhRbiOy7aFPdQLGetAsI/MwgZR7McHiUC9Fgob6+qXSUsPdDQYqj925Sfyp7yYTe0v3EPvH
b491rcM16BgMqUSUpkyTaYEbzzSLlOc5LtaDj+k3f61B5zAetxZqMNlUtEkCGmHfj0qsw+APEZze
oqHwWDUoYp/Se0Ef0JzIq9Ef7RGRz4cHO10PHqpGbyrDvZQ4MSmuYIGzsmSIDHfzWc/vAsNczyiW
T7krEAZQjMS+W4SeUgb3jxMqwTVizInC2O0EVWRCeYeYqoJxkhRykVuNyw5K4YKMt6xw0Vm7krE6
kSwT+2NkFGrXo4rJ60H6wZB5uvis8Y10etI0ptSknP9EmnJ0Dm3TM0BqUYk3jGh5yjrXuDtVBXxA
VYWuXrDA2d/C0HCmZqQlXP6C0OEnIlC/zlWFeAu9+vkLbHumXtT1ToHtnmvySF0rrfjQmjvH2v8b
Xw61YqKeE8iNPeWd2VWZkVT6UVsFQnwFVAHzcjfi1GAEhnd6d2S2ji2zWaVQ089391mIzBnYXNzJ
mBBDIDz7JD2l+e+N6Mh3mL4EVZQGo4UDLTSlSprCuQCLf3CE10+Aqv2+K22R5UD8+nu0gnnCrOtC
GPYW7lVY/S5VK8f15QFPpR9QlyauRZt/u1lsbEBSgCUncXWdYpXisEQhrBlT7PIhX0L8a5R+/wua
7SIUPg3717UrTOwMmOUsIkmxjKTR6FoRaK2zgdyTUjtuAD8Cjf4qoM4YxXoVG1mYNalzFO16GVwF
4Mp7UpGhlOMtvkj1fyaBXbNm4h9b33DkP1Ta18Z0AlIQPB0likvK4bGTts2iG1zidBvyVn3xYwqu
63fwpetzml736wUCsOkkGCEwMQQQWGTRvmIH1zAL2ZXImvcYFgTS8GoJ3BnaPsTnLvjhm6CCq6aD
mGR8vqMEOdidHRnHyi0F26rsnBnGTAKbg/bqyRFh7ciA8Lzmux7gqOY/ZFWwBjfGPEJGV8lJYnNe
jNsEJWljixRgswfoTYS51Qikfyug7tdy4/oko3Ech1X5VNn5Vk14/6MNHwqfPvebJrgqNBMq6gVk
7atoWtnWy7s3LmEKXYIoNS8sCIg5fLb7CMpm+DIV8sakTsW7gTU59ow2xp2z/JZlmgnJbSjcXplt
ggW2W4vdIy/mpqL6HQeqM8UqKgrJV1StedMz4F/Vxc1c1m79sPEUbPAO9gYF7xJZTtb2IcyfjfNZ
Z6GetAaIh7i7EoPcsm4MoSTxiNn3EfRwYLcUEmj9xBgt/xUnv486zfTUfNDba3amyCPK2WUSxoXI
CoyhIwqXxloCJlhDOyNb2VrteTgcaKSo8gysuBb2n/YkVu3PNOCq/p/7EuFcqlZkG8rTP4ALuQb/
RuXiMNBTpz+T+jQJVu05TumydFbcuHZe7dSZs/28xn1H0UFmfHWPa4Tcg7TNuQ8oZDGY5J9qsYRm
/mnm4sPewjq2tY8rhF8DqGltf27sbF1ugY21MwIeHuG5HqAKy4o/O0B3+8uoEz4INo2GmZP2zd2z
FDpPX7gX+no9f4rO98WSmlX+IxywVXtfPJISwrTArsJkX8X2K+lkyJUAvrOeF1lc1/r0lxWWpXoB
+KjwbIKWCiZIafy75antS5SzZFwjlxa7KhzeR4eYSp5NuzIp2wZtgij9LdQ9rGKqualx5YyHSi2q
xeJc2LbtXsrpaNI8mJr+orWHnyJq+LHXYE3bMGEAGDVxnYR4Fks5nYSeF3brGHnwHFyopwGgGrTW
JLFs9wX4P0yevIfKig6YvLAuweLtTvidt8flndRAbguCKEWkhcxOtgpW+Cd+Ivx2EfdqHHHxKwfI
Hbg99WQL+VO7nPwfdasfyyXcRyQ0nrLUK5KdFD0nNDuxlBMLzioGFq7Auw3hasW0n6cu7tvsv0u0
XyU/46TjP6ab6b3ooPGZaZZ008nQiArxuEG/BEvH8nQGMkTuiEZhpqUnlXSNGSB8SY++TCHPaywa
J6Ffii+7uWyMMUtPoOFROSQuFWZ9U+q6qsE87yJi8TddmKD5Zde8tDxy1jcbFsej/OkRBYwuHKrS
4SEbXfcP2licBznC7qjE2Q3SGhxDNudnDguQn0lkukIc0xgQHniMH/LSdryvxP/TNyHfqdx5I3uX
kNnamKTxh3CNO7qhIuHG66wHxgpqJdt7pYyq7lVgKHazVtfzwvuBxBQi+7IkD+ewCBRWbzVJ3D/A
wuRJ+98QT2aVIKLcOPJ9pvqE0DmzHsjvBtcY4A1VPYhFGoTo9dgA14k16PefXsxSTvQ29yP9PM8e
nfoX3xxmMhuw1+3Hof0/JG5HbtpLpc8uBrf/feRGb7Pv3Uwr1YrQTuIb90kjdYwy8WemrJMfdyyk
A0Adbd7ynXOw8WDHqfO7f+yJOs8Wul8CWlSTDrO0L/QiWX80YwzXqk1VBgxDo/T/9ul6D4uJSMtF
E8yW/Aj25m4HcXq6c2d09lDDLQNtYrXnz8nAxFxD6Hx/WpUkmn93nRXIzSGgOnr9xHg6RBahztdf
gYH633glqpAmy0jKNC3lM9MwD2ZhHbjHaZn50zSR2ACdnY2dqsl+cdGtDXVrqRnYLDrTDdHMuMg6
H/JSg5gHna0yJoHJBR1Tm2+ScODdSimNBybQ4HqQ4GAAVEsEVlERdVECAmdFao2sNxmF5ESOX9G6
4sushtPCQL4e7Y9m8O1b5AdVgVc5T5tGmkj6ZCvq9zFbCniNgMVAQlW/WF+xZRpqZwt9P9RF5apg
TjWOAEpfFNeFRrmmSelUBLauPh334r0Fp0jvYnkWcGt+VIPlmMEiRDOxmC8Jcw45tR7UfkWDUwrm
5WIDgX2Aw2MOxMAPMdK4RPng0ZepeXpKD1E9l9cIed34MVt6bpcTAeUt69XyLOUa1MaWKbKmh5cj
EvDs0vkraY/RU3gEXGMiyITqfla7V3FwViviR4/BctKTDrR44cua8KLx/yf1R1o80gyWwvppWpE2
qq+AaB8j0BB6e2Mz16qwwwiJxSbG9pL9Iw7OWCfZjFR1+0ZobMWMVh8MQr+BgfaVDyThAB8BDGs0
ES8IVuK1ABnBC9rBk1MQioeGCq0q0qP1sr22UFbWFOPsa3VOTo6xxOuDsR9cMa4DiTV265JeLaRV
HITolDh7PWJO9dyzHni6qLeUlhEzxZF44wjJ1Sv8vVsQbdJz017/iZrHH67zDoHqBKKTRzuUsEuw
GwZBRZSlYYLbcjpG7mPPp4v8Xh9Lu/dbiygeoVSPDtRtF0rVqI6KwqQdSQSy4HwoV5YWErEJc1vs
830p0jkybFj2kfx9lXOj4JupxXypbPLRuxX+ns9AE0zCmzO8T2ByYrsMMXrxDMgoV37c1DVttHLA
xM2fnjG73WLwy2G/MFtr6Cxsc9dLe6UtOBOX9PdzhRBt5F4wWoEMAQoWXVT1v1pVfUgWmYdQdFKp
2Q59XpxDCBg5zh4CBP/u9kpk3V4VOUZJxW7RF0BVHpaCYmVBQqPt8KEECAop8ZCAZdzZBwnh6Qdi
aSmffbDqegZhHr0R8RM+gASzRVqAI3f6XHUsDoJyEs/l0AAmXTgXYaD3shJqc0C1YyZQU1IQdkLo
KeOsJmlbMO4ZrsWoTfaITU0SH+gMumiy5dsTiH4RGOru6cxMq866OVzEu0tSEUKTabNDmBYa7KGX
q45QE1tMdTJ6cQ8HlSGbBpficbH76b9qisPS53aEd38n+FBRRp+XAxTa4O4KP2EKaJnV5P83vbE3
8EDEQviaAigIQ9ToOru1hLRBt4ar9Ueo0WLvMGDlTI/zZe86gUDMSno4NylKD34CARNXW902X6Nx
zws4q3b4kLxIm8JaaCu7jEbVn+Ln6tdDSw7y+J/Jbm2HVMHI5QenxxNXDgvpIBHFLii0h8vW+Gz+
68u4OI/tUW5Gz7jnD6IsfjLVNqMIt5IgIb63fGigXT+KbkgQcTVMOvfvlaBfjGkjBGM65PKQT0/P
PrNFM2L4RuunQv23tYBYCGIzV0UFaGGcJ4RtI9/UadCSODy6O7/8m1hLsbjdJxWYWRRJQ+LG/+Q5
LdzOpM0xSaMAMfR7z2w+QngaAiRNJhUSinJU5PXPdNNQLtWszN8IenDa8FgCrORMiVD4gcdJgAF4
GVbP3A+pEmiycwJmk/AtkfCYTCQfmJFAKll0AOKGr5UmxIR+qeRZr9gLrz1FCLQEweKu52v7KPmD
iNUY/XJXLmnkA6ocnZc3MnkOk4nmZOWrUvA1R3N8HNFcG8mK/SAR+V6gYnaX/GZI4nMpAV/Kcudx
78Ggndx8eXY1TLW96fB3/Yva2VHGa8CuAACRxpQBB5ZbxI/5UcyIHwgEk6RlTwjtErrNNgkPpMRM
7O6ohlrwZdyBR6xSSGXyHNZvRcwfdbIEarFsHV14vh9FkAl102nvJf3wCMitmyLUxUuqYOACQGzv
R6Tn1/ZjppM6rz7ZKov+2C9xi5+ZGVDpsA/GfvZ3BVvLwfHqrALH+i59ad2S4Yf714oueybVg7cz
aj4gRGMMFHcSOerS3rR4/amrGwgLq5KR9RbbhxB90aRdL6NmNKSYDyuu5zlkLQL6ovTpYqv3ghE8
L3b/dGuUS5o0UGl3zBbQJEew1xv4/VHmW6avD4sw1TP4/PQGiqJ1HyXU0+X1UJonnZNNtu5xz+Tn
j5+kePVE/R6ytMOQ+jCBxMCT26diTGP7RyESRLvVATA2vwtrFftWSAsOP968aSelodZqJT60ce/J
uhkF+byTH1wlPrBqsCpXYlYd80RZI+Sn6rLjd3MDSyM++jqjI899tMJAuBYTwcFQu8NxOuJcglEq
m0xiTekGQrzpjRYl614TME6KokO/LpekvAx9bcbQQKvJQ+WocL6A6yhFk0w5XWg2CLJSpeMnm27P
pAu3Yl0E1gOmhC/rxQSGBP3b4xwwszXIfUZAOcSiqIJ45eFj1pfoVqcVR9oQrfVW/12e8NHERYMG
0wOFcB64s9EQoThSa5iSCB2aSMNSBS8p8MJCktctm//KMmh2PebOR347iI9MsnbQ6uFkoelO2KlP
l/Kh+AK/SMr/zGVtTGfFHCINvLXqGfLMQBOrHo0XalGhQeSNAGoQZyLeL2cie0plEiSy08zoREPD
C8SuepZ39WjmhqwukhyBVkdK6Md6xqY8XAMvKzeIBm8ubuUZmPrusP/KA2K7700czpP+PA4jS6Yw
YIistJEXwOnXgS4mC/gS9AMcDZloMMNnPouY87T6W/fP+f/ENOXE1bCjOUvrVnEuZ+OGmxeXCcVc
Omc4fbWDZF84FTzqU2KVUBsh2bZGls1wI4Pjuxi/Os7HfOY7YdWZeGOaPh3fCZvkU9L4L9BBBulu
7DyV2pAj8Lr47SZnlO5tnvP/2+87XAFKsqo72dCHMDaXl2QIU0YRxBKOHxoQ+cmgcqbVke1n+99T
VU0TzEE5ERuh6Fnhta+0PT/eZKQsCmQ9ly2Y7K1IW2lDrszJO6Eu1j1sv8TaxbQOcDFtldZdYSwE
YMlkP+PFeHr2jeid1IbqiTtv9/dKPkITAvBJ3YKbHiTx3Rnmdjl097D2QQeYTOUmI6a+8VVS7/Sd
ONbr8mdJ6nJ4tzjXF24+X+5K9/eEA+KRN55JbKmtM17L2x5PylYw3JiQrZhu05ZOSNzHK6hnhCMv
xOg4ULDPVn/DqHTs1LrJkrgj+cnjXtpzg/Xgp59ilfMXD9W8J8/U680VnM3+KAFI3qK1Oo214xte
mw29HATS8DyLQWVV3Fv31ZBE8v79gSsPlKVt2vuwLIQF7ZyxJ7YtDA5UkfIKXJZYTlv4orxqczWl
8Uq0L89eMv85CHQfaSo5LtRgkPxUU7dfGBegqa29ARACn/6HFjBssXO5zeT8lbLGQNEF3dctdfaf
Obo0O0i4qRFvTByQncJkraQYBd4q65w2piPVyHhfZfoFIaVayg55LJWA05MXw/foRRY4ofu9ZWGx
DMdVL7qZ+It0sIBq5hMWq/caslsnx3/N5eapiCQpNfzb3LYd81OYltNED0crr1lfyayWrzeIZzib
O/e3+F1Y0SNF15DZ9VBg85redqweGiA4fqKkzqEeh0FrCdB6pUDs1Ly38f6GxrDfKpyzFwaK+EkG
fG2TMLnPhLS4JU1FOgRE64IKDCNbE9eAeuC8rr/rGqI+ezpodxaaPSn4sqVKPXQu+Kr6m2HVmr1j
d0y4teQYRzvGx9zPFqxjLpw7+eZsnQfIzpJgtuFUQkHbOXv3xCjHzXWXMWu157Q7BHnqClTx8Wnt
lSbqT8eG4b9F79WBS7Om8h92slsMex9elk+l/BZ2bTo+7dJIF00Lc+KTMF1v7CAidystLwN1ICbq
Jsx07a9VCMm7iYR4n33OAEpbwPL/q8U8Q0ghfLZ2yJcYt4avpGuXxPaqCup5aQ/d2Is5UpzWI3ei
n5B6Ix0blzivkB7eObno1LJ/qmyQZDoJcnSNwtPaqmaKuU0sUsoKx+0rV/lY+zILl6wFVJC+T7CL
OBSVBA2sp65s3L9MrlERedLlJ6QS4TZOGO2FC55vqDU5jWFSqwhdUEaPqw7HpymmobxYFeOg8wCm
DXL5H2Td9E8m9Z0q98fJKExkg2olQwS+8TsxL9X5udBBkc3rFw28heK/+dQ/CulrQIrBaOjDrNfp
LOO2CAaXxy7OKtYrM5+/QfuEx0/fXUbPZ85paNsa1mEHI608pE0cAJTEY759jQ9DkVWxtpY673CO
/ETHR1vYYyx3ycdgE3Sm2vJ7YkMIOeopw+0oI8oh6W04sXtOTdnRlRGRCyiDK8rdP65JkGL1cYPs
WHe/Q++6M1juRomyot7kbxgaV02w+t3nmDhqhHUJRpj8cL9EIns83zCSbQ34ctWd/A5jmvIB0x1u
vNMsOJcXlYd9KrYLqtbXyJrG4/pcH9n0Vd1PqUlJGiPt/Oo8DZi4vPUN+H85cZhcJzH9+mISyd6R
tS0oo52jXz8m2050dSv68tR4Ck13akuyMCjEGhcCJTQPfVZhJgeLou4f8cfF7BV1eT3Ge6kFL2xN
aOxb+sy7gvxKPdpTUt52JALFjGlUY4G2jIyAWepZiBOUUA0oBW0O9KpXMu65o2D7op5YH6jAFIvc
aAwE1/OJS5cxW0fBdG7HlFrqLH7Z4noXRRYy1Zgg+fzpGxec2IbGMzIMLUe//S0gPZpaPvXjTLoS
iCWWHmy2sMNiYCSmRXFU+PvWxDNHEevdxhRYXR+hFPGdvuf7MWw8h9Oa4pzmXnfRWWVsJDmZXdy7
UKTXriYid1LeN5JUXfVD4XhNwvbbXEPjEhCP2S+mOTB0olv06YjgHG9UCiFB5MrnIW4xuJLedPVw
NOEXLAsHEL+rRro8QBXu55uF9vlb0O1g6fWv05UeD1TbuLuOCu8BYnCOdI4Sh6gUgx5e5l+rSTbx
FluZujePLvoYrFURIrKYaN7OQG6gJ1ahnpxXnsJl/HM69j9gxnefEGUVPSmM3UXlzmY1uYjH252y
YnTc2iK3Bc1xdEN4yhoChf2YXMXZQtM5PIv3zoGRkwUzNFR8QIL4CYc+uW1oJPTtg9kDMQ5tXnzu
LzdtPxuIq+rSDk7dfno57S2golobKE7Z8sE1TGq7TIjRZcMZ0OwKReiszV553F8JPp9WCQ13pdPT
GD08dnIvmX+kqlK+CCLjWQUidzqXtT1xsQg8RXc9e5HJX8Nk5tOtIC2caN50AJW5BdL+QNrSNf5b
yND6aLW2nncv4WUodLotJyRlYlDZzeG5vsq9px2VgMPjwYXK902QYj4788weiFDIihEgHVAaMZNG
7oQKPxD6I9UIM7tx7iYovp4pRiiR4QawJt1VOi15axhRHJgeOOIGaQN5AwZwlrrHWRuaXcu/gbdM
4Stt2Hyp1KtJPHFjixNvzv0JYx/54Z6c5nKfCsMfEkGCa3zMnAyOLWP+alDPMFjukBKFBhFmk6kB
9/3FTCWp5u6YXKoxSmEw3GTfJ9viyVDNJfq67zTFx/yevOONyoVuND2ugdVqz7HHkCKM7J9u/xdb
nAEPgt/msLSi5xDBrVSyt6yTbwqs/tKtaLE0JkklWNqpEqwKIjeC1AkOoAI6QtS5pKLNee/wFIVE
PQolEhGXGppudi2e/ScKcMB3roOpJCnabbfTgmFJACwiUxhG1Xeh5xeYDLEhDdHAuU49I/kmYUB/
FIRmMPP/lXugHmb5n/VFD04Ue1JU7Tp5WqlyI/QpKAM2VgPmNW6RDr7DaAfE96zFRiv1r9/Pz/v3
dGJmc81ZMpdXKgiiMp7TnihK3WxEFtoqrBR2t5qYtMem1xk3kH0vTgFJRQbQ+o03ZLc8dFPbh72P
tGoys5NTF07E9yB2yY1FF2U8FuKDQr0yfrnDap9fQLEZAeK/wUe6KuxurTBuQ84FRaFb43pJq43r
rRZIhRqMFuiGDnwh/jhV+XoQVuqqzrs530EILKrtONlD+5zMzzD1n3JV6qzAQSo0Lcb2A6sNDYXf
zmLx51oaiulB7gyVrkifPN7C/JGzjLyVGK+b63Y+4c959bJAxdagt+8ybj7ybnkT08ywHGS7kXWV
UdYi/Se8ShH5Kb9JrYRaVAKVRQgn1dYLSM+r54kEglVTx1wLMNwtjMNjhdYhTWhi/biwBOLWqSjE
4jJDMnMoeZ5JFusshJ5qpVfV5MVXDvN40JFpptkGpzMBbElzwyboIwaJnHk11rVa/yoDjkBRVOET
QvEyy2sFqZVZSlXVIYn0Pd0Eka8rnKk452Or99mAWAqioP0uP3JnvjksR7oT5iabyugA4ufpOY2M
VkTFgjOfUs86O6975j07APC0y8ezRVRNk+awh3c3c93iixhuni2HCzZfh8sPhb/FLiXQXUfpC9lZ
J9ROVUDoGDJTlu6Bk3hXUaGWK/CBvEBO4VCqKT+5Ia/NsJGhHd79rSN/EIpHS8j1rZOZt8glp4Qb
siuYqFesTuRHjL7B6D05t0ilWt1tr8IyJMQYcdwz29RcHkznrfFdcJggrKf7F8onOobu7vxqIoPK
ZPu+eUKmAu+SfMTGmdgEBsAMsoW1UxiY/p9Re5pRFYG+0LKdDBcT6/HS4081/qov+ux/roHrlWvB
tycxEFuRtoYGoEoBAnlcu5mAr5tBua/YOuROPCjRPCYurLsA8KuBx2QbW+cXcRFMJ2UNE/d5Ldag
Jz+d2lLvUYzJJK40M+88wxXp1u0x4rpZtdvbZx7mkHafDOKRpTVPpPlUjgLZ2/x/xO9NIpT7c+py
v146XWrkOnJvmPXpg3UdlBGLv9KCXQ8Bnfulo3TEdpxn9kT0tLNeg/SQuBDzk1dzOe6cDVdrSCM7
LF0VjrPRqaQlDuraXdZjIop3ZDse9XXfbCXVAbWTLfOJuPiwTthUJKahnnlj9xu/hjlyAvW2YSNM
NLF8Y9ysRZAYZupSZOLuyV0w0sncWMbxrhuDU2e0VJwa6bfzXA9LQBHkflhFgLK9+1/TB3XTrM3E
2OrKtlmXCCITDs4N0Y5szfploGGsabu+ggz2kG4UsGBhXneEQPWOM+58djjYASqGrOZJNsGkj70w
M+vOQUYgQ9GAWPtkXyRomF7VFDjd28F1r/o3EC6vI25jGnXgWXaQMomrsIzyQRJnReqFkcnWjXxW
LwZF7riY9LH8kfoO9n5lTG+dzsekc27y0w73r0xt43xqn8B9IugslIEurI7WAHcjzh2ASxYJv+nr
V00c2I445kgfNbO6id2A0KK+OCSJknX2FFl8zaaIwRRF9bIU4aXMlMZnv7dbVXN/8tlrYNRqNNBv
ki29X/rNRI3f8tAe/Zm0DvovBBxwldwVUJ3313fH404RbRnQ4hlxsZ25PrL6c9CEmUajp8s4WV0K
CowWyk0ctc+RiH011LgpVoDWr9ZHrE0O6AjdWBuub370gAoFX8dB4qaJk4dbZUJWaoCWyzxOXyjb
AVjMUHYtoJkMfYbl59/VDZ26e1qL5dCEC2y/R5naC84B5i7qBmIv2k94mI5YJ9vitxevoXWrGcju
GcOr9pUPsuca4F2dVAXwLdzaBHwxx7+hEVBAsDeJPBDUoEQK3Ah8sTdoNFXzmU4Cm85ye9d0xWkr
xcL8S/2DagjRNgEgXArhyr1hF+bLtSaC4yBrlThSSPrT8PlNfgz+I4490leZRHwGlLxt5VdCswsR
5WAswrWviU6KcRnejg8IgWXPhAW63dXD/MHADKMOxWWgUs18V+z/KMflZ2SJn7TbaZutfgtZ68Bz
lQDCE+Vs67eC+RUJ5zdPgoy4FkRseDINb3W3DgQsBK1/He/K8ivefaFV8FyJgu0BPZ81DMS5j2Oc
SODaCU4nEBUrswS51B4lONrY2IgQQYj8WhOUySury8KDgsR7DbO/4/MJWCvPGTUabZ/d2qAbVhFa
n0zvtq2zbe9PuyfXf6QLXGxZtIJy3i7SB+s4IoIM7NLlVhAfDm4NXR0F1cUyWWR0dcF1g++0SFda
t9PD645ryswKd4ZFkWmc7ZoDhXzfB8Rn8rQGZNxLye72zR17EWSlSujn8JIsiFwjurlbwCN+WSbQ
XpcrsdDSqnWD5ylF0gnn1C1BrJdvo9VEPE2aiNX8y++ztYU3EXjsMWtDLQq4d/WDgzWacGVQWU2N
k9OFLYjUfbfJFoGE/rKAJXnyBJWfgWEbtvQ8hRZAnJbMEH2/kRzI22jp9C9jcE943QJn+1Ki9OQb
SqbXwdZ7Rkjv2KZJfZb1I3a9fjTDiODMhNJiee6tdPpq6fiQTeSQ6t9FVIJkhErZbuGExuknZYKE
kETySoTbr7Qr7aBtvSl+U5Ur31CWLqI3KgbZckTOVf/graqRkTD9v8479UwrwH8frQuICi0flsRz
0qWIRiYSLCKYOhU/6Pc2AaVj6ZmJYBtE+Aowd8TIpNYMk82XZc/HCzMamvpoNM3Kyrz11dXjr+i0
a58ToKK8ryzBEI1mXgaAMV+UD2PX2mt0nr8FsKN3V2FjME/SOyW+9s7BSVwQ5Fh74ARC4syVVX4Z
ECmZmKkX+jFvOfxPgoFiR/xwunprjI3/Zjy+1FNDwXsEucFlA+s4mNVj12G5NwLVnFicc71pGRcH
iHYIKR9LtbZ6SV6s6khmQTEIRJYhlVCRXLP4+ell0PTqrBc4LCLbcX+8v5QEEqpVg8aRLPJXd/yc
bVhabFSmBELF/nneeEvzR7OspsMeSQDTjRgNhmF8a/4zSqzcIx24vNhPp16nyWcAHYGWgnKz41up
fNmGgHaw0lVGHNV2kt5nABWhgEVnUiyapVsOEDu3xevLdn0O1JlluPkSIZK86wMkuThOJQF6+WDb
OY1SLPQ5F5JbFQxRNLZzOkii61U+RkLFg+OYmdV6JhPQeXR9AaZjd3HpAdFs1QkoNWqOc4ocKB1Q
l0hDyHlJ8SjqP4CFfeflOJTO35jmOo59k7WzfxWx7hKdwALvZPgINC2ETb555/g4VA6PLTfwwbP5
iKtwDwpgo/bGzILcxFRhfFQNkYRFkDOQIAnad+Hnen5zmnYGqIgHWWIXGF9zc3z7H09U+iptTlDE
zsNdPa7lQka45j8lGs+NJxijAhn1neCAxzytkOSaA9R0peAt/ylhmQWYHByc5kecP79GcmXmZk3D
28vLc+dROuN0Fhs3g9FdGiPPtYXQjqCea7w8CmiYZsGUIbDnSKcsY1gVB7MtZx9hkbRl6KeSBxNP
RMy7o8KeRJZmU9MCMYH+Ep6gBLoEh2Qjju3/5yXPNtQ4nZM092AvN1H6PNsl3tvjREojAh0o/eEk
RkcJ+ht/HlXNRYhimDkAAGykEvJenI9tvBW0maJELPLjLEL4wvDbASFM4QQNn2AZviGA6+9aNJna
tlliB7nVFvI7Lerx8dU2F+4M1AJoVcFEWLT9m6mptqh7UgzjnP/apIBzTkqm5kzqITl/2WD9c2XI
kLpMDj5hRsBmJ4ivOfXBfII0zFWXl7xLZ2EVslD33le7cuB8+8iBVHZm4q+AsmyWkn6ZQYFv7Qvg
zwE6We+kcnFKGuTKv9Q3czFtUCKGbKfmbBCIRsDrQUENWgGpw6W6FAdxSDDUznqWlD0fp9VGQmw5
YRBs38ympb3ggCFtz0vxRExQ3hH1XBfbBQaJEKBbf/nLcpm/VsIs0aVUwCLwJq89qX8Bl9Xqm5ZB
QfLoAfm/wcIEfXSpry3iU75N073nxTBJAJ1ncdbyj8wWdM73nVGYemPfaclYuin3hOPOvoW64plA
hS2gMRpdCjncC76jTeDIuwAnPqZ+0k3waNp42OWw+mpolU7UDVYUPox2F2ini843t7Fm2UwPm76D
4WEX9VtZDXUJWCd/7Ew0Cb0FU62z1WnEVlji4ynY0TaWX5oXMONNfEQpBuw2KGwQnSAID6jGaWfs
VBO9/gBFw07QkBgG8M51c5Ez6ki9oRtd3v0ih4cWOe4SVeOViCyr6uuYxSFxnYgxJ0wDb+H/N+vf
EzYcdwIT2nTFY1b5QciOVzHFGmgPdZY9fJ8zHYIXY6lwxNiTLpgGBtT66+iaNB6Y91eNyDv8FXyd
sp3Qr5Lw1bvBTWtXwfUCJ3YiNZPaAdIOT9NZoM2lfUSXNHZSIfMfx7HWX3k15vqvRNg8VmRefvpc
niuuHZ4y8AcC0QbjG/aryPTJvp8stk43YqgHpPB0sUmWPtff9Ew3TPviKWk4asSq2jgYT5KC3L2H
qcrNSdW+7RDVvBIAqvuptX1685IBWC9kLgasGq9fpNCGM127nQ1/LqxG35kONb9dWTGq/llRgq0D
RxUw2pSPg9c8wq9zBIdIZGqh7M/6MI2V4lAqBhD1Ujr5SDWqqpBaCPesXy/19xUzo9BQa73m0CA9
0+entkmqvpJhiXwcXZzfzZpRpEglUrCoFEflCHpvN0m0AhsQ8bUuLtEBakAsjNdETlsB6SMfwvKU
yWQUV0G87C0S1T+a8vEebB2CKSXu2xPqr7UKK649YUpy5BMnHrVW/n0cxSXe1oFLdM1KJTAs+/GK
uYj2HBILsLhGZEVuIykoalaXP7L1j1nplnt6CWs4M09IprcjNAbJgNaePirD+XsrBEJFR/p7uHKa
koo1evECnPjD2K+2FUXZmFN9Vvbce3+G0183iZwlabkCzmwSCcgtCc/aGnr93wwwgY8jrTaQoiIw
ApTS7slIorG8R5r2/30hZ3lV6LA6X51xlhxdMcZg//AqiP4oECn7/4OoNgUMDd9qSqUl8T7LO4Lj
rpmppseS+rtWArfCKsKV1J9p0dEaTptTs/IWyxYOGoSd+cCovRtJv//yhfcJBKVMWiKdp5T/pW8c
IhNK8A3gwOw67lcr6VH4aPHhYScS/YseoJPXeBPftJ/6yFrE3HnsIQEpOAxYFTQ6nbzJjALaQzOd
oOieqoOTCPFrhDdw2okgjT9pe0Nu3lo83Fsb1t3Q2of2+TjbwQNSW55rV4tfsObhl0qGSGY+q2LP
3dtEymF9u3U9v8qa587kgtXvN64TZqtYl0vgfKD27asHFAC+sY6ROfcuvWXF95CG4lHJIkEVmsXI
4AGiseH+0Ik0slnDRdu4x2kiMP1bPLVP5P30j7ZZSAHbyqZq6lC6PrN0igfwpQCqJXeQnafI7QFT
HhOZmoSxiKe+v5MuqSHgw4wgu+VWwsxtX4g2srIPlryHg26FyBsRhePKMcd7gtFAbLC31Io3Jpl2
S3818UPpx77ZCA+dBL8X4eNpKxTdTDgm4DvGYWO+a5XCixv7ou7+6xKZJLFFc8cTpuaRmr8r5lQ6
KxHgmLDYWevpK0c5xcKub8yczhh8KpLlMgmIwgBEzqNb23n3XxY9bBAEiehAFi/3lFQzzDN1JqnQ
OZYPsO3Kd1z0MExnjKk3huP8xDVPC235zCyoSPx8ch3ir4exRfdBFB9sO4yZ++ijd2blFR8cCmO5
WAPSa+WKMCcZKoXerK/AORYEMWonjdJPVQZcZ0N6GIriUyAsDNmUw0Otrsbr8mAUmq1GIQ3bl692
4vLzx8IxmIjEhDSJ8NBbkiGK6a7P6VqXQYiv+hK8UmH7sQzpG3pnbiu/7dgEkBt85TZFnogWcrke
d9+glEqQmOnXusXWBrC6jhj5Gwto+yZlwUu5ahUW2Bz4csAR85p/iAwl3u8QqZbXke2ycPT378CT
J1tIkwUhTtLjeXHXfTyrgiraaoQ8lywu0Mz0HNo8Rtkn2CaqNCn0ENz14a4lZmzwa2mRx9i0+KM7
S56q3mFDbgTgjAD+XFBr4dyilOHXdSvhvtXeBb1bznCMX9kwHxhLYeH4Kzu18urh0f/m5UCN6acs
TO1reJ5euNiu6wnl/8DI5CNXaSYLE5PA00G7P4Linh/ucdGo+HdhpbuXFqUPsMqBtnS+XOpR4Eva
QnEi+21DxX7v+Yep+QAgAqdZa5O2fB/aoFWZuYKZRQ2MC9KYG1hDHEMsSVHvGjT3WHLFEUdrSWg3
thHLNZl2v35lMsam0tIl6WrwbwG7v5XxJQ0euU/g02lvg1wmtYFWnUUy/kPK3hI60QbGSAdVVZO8
r7exoBFECZooKZEx6Z8ayzavw8Jwr43luP/Qj26u7y90ekj/d/w8mnr0x1IW0FVp56ss9X7fH3Jo
iUEc5EDgMFxo7iD4mYd1r65Y6y2yi2LvM3tAKdIbfhXhrHgXvHXgWrh6OGV3Sr0Os96XfePI8iLL
HS5BX88PBWvDUqZHjL/JipVJBBcqrky6t3S/S4HT7roNc9L/8klgcTOOAqDXvdnWjzBUYXv+FwdP
x7NtIScpSfp3W1hJ1e+MP00vbXYBxYqeLRzNbSS6LzYHH5B9H+20pYojxg4o2tKqA33kk2xEawY9
diFOlhKxhbAJjhIDh/EmEaBSKeMEiUoQ8AHarFBA/6GT67J15g3sa7UiWL+ymsmkaVkoIEeiIrVZ
iL2AKR6aO24tnp0yNC/h7jP37khNhziER+QJg6K53QCePpSZk5wlhKbynk0mbrrF3c9xTw9KYYiE
WnSc2dTSuJTYgP+VMKjelosc192hdUq6tvBU0oVDJS1w2/HNTQqJnvJSs2tw4s4xtmjPPHA9ir5x
YEovRH76nC5i7of1ZkfpiEXzhYPqS7RbzO3M5Qnk+PlOjIkk/G+8QQBfqR0vOhu7di4jY7H5mt+T
S9oAQ+WvAkqA0driUu1niBgZDqalxCXMfKiHEwDvaQv2CSsExwCPFGOgRVxRXjQlAU4XiMBO2kGF
88PJ3WnG7sH+yYjs2yETUQfLCJxoXc/F/CrcLhXu5R36yCLlFJBZb7dj6ZBjojw9y+Sa5LPUmpM2
HX6AvkyjbeSl8Tsq+lDV5TvdB5XaxUaemtJfUEBieDaJYnbfwZTEjK3n9ZCYBJj12LZNCvK6QPGU
XUqU3lQN3EI0/Zdt2dkNuFprCg60PC6r7LqCt8iRuCdl0QnaNJzk6nEQvtz8Lcf/3DQa1yuKiPwT
8mjWZ+uDyKa6S/kjKqCN99Ju+D+jOuONeK7JsBRJsuGtwiqEHIc2U3glgDlVXbobQ6ECeCryQSbN
9PfV2xMcWNPohoCyElBV0SS8ZpQppyKbzfTXPb6xv4gPhL8GZiCDbhgP1J/Puf35Tw4fnkdEQzcT
yOHE9wTWj6jd15vAJMig3Krd9ApdPtO7FcRgDksU1N9ARTJErERGJiPjPVlXQ8MEDaPkc+WylywY
Q9onDI7KvVDOFAFXkhGHh3BDjMGpK/T2V5jzMsfcOy5oCjpNwEzyV5MROBSZF6J9YcMCUnOJHygW
MzAHYZC5Nc9HEQvsi9/1zXxayz6YCpyHqRnjyI0KXyp9Ff85maPH5ccHkelCdxdK/kbnmwM8etXG
vw1O3xVnBJ+HVpZVWtcwZ/qI6o2kREENDOXPP1RXRmBKOwwpS30N1iEKWFyhX9ZpCiQQCIonmFD+
ZmqsjWGaVIlwAME0mJLGsDdZtSD5xWYDpm7/REuxNclq1kg9tgnweL7FSiFfqYNeKCr8Z34ZhYJ+
AJUyglWMRMMRRW5AmgD2ghuFar7QmvePzhGIKvsT0zx+DnHcZKx94/nnl8B21DryGx1c97GzPy3w
hCLWshA4RRsM9uB2hj4uasLuMPVheC/lhyyZU5Vi8t36fPxbKtGMZXqT6ESW/xcbZjmcWvidW1H7
94hxsjb0FSC7xO33RcqSTMksckVzB7A+FFs+CKXsV5f/aIAebBFjA32A+8Lc2uY7UiPnyVBxtUzp
Dj6uZuxOr25R8UfOifGxMHBGmv5WGrLVtxEkJm9pbTGguGSZDqe+hA2yG7NCX2gXENTzcPVPNYPt
Nwk+AIYlSAtRha+FWOxfYg/6LtOFqIMIjGLg8ClAJG6TlrWPooninYxSZD48eVkY8Pn6T0xXboIv
g5uzo3+yJMnUm8tU/uulSuKjfYpJUnYKNv3l1In4asJ+6k1CUjr/6p03w/uKlG5Jk2ZNOOYtbo//
JWvLhuFwCnyxOqpVM9zP4W17Lipd754lpLlE9yDpHJ0FTHhxDG60N3WC9FkbbtoYWl9UOFPdHnSC
pT+6L5s1s5smOy/lrXooM0g1B2FEkjWMvt4+ERurwUfTvCtVHNtuf/1Br9MWOy6X3tfVEdciWkbC
iUoBSIU6ZeRtuFlulDWp90XyEeP8FKjTbwCTEHHdPpoIBWsesZWxJYXwF3ERmyGkOTEzw7dNXXCD
d2VOEKMP6+KiTM+2LIqg/3idc39+gDZdDbQkSoYKNP1j5wTJbzbzhj4vdCv7tIgJhEvY7sKLZWlL
cZcRHYGY9ZNUsHoMnAk+zHL5DMZfo1TSxrWqcjxJtKuQhMNTnsatFEdzXLoc/tmlm6a2PS/UO3Po
TIyIS5LRfXCGP4hT33AQCcc4yp3yfjHTvn1qyll+JCWfvFhIxQuWVfgU5dwG+++dFPWft0tOm7Is
mvPRiaBq7XBG+cU8S2UNzlFLYn2ijneujqQXuTBfUu4fcEYZPwW/YgMskZF8NIwZ1PUJ+vcw3Mca
QyVOS/YEXOaeagKYkEhNzRsxXHYMJjbec0o+41DnNg+nyjJaKsWvUPF1AtBIXcEQ+7CXWV6TtoBx
eqjHwlfFQsJn6Wgwn9bIZWeUKenJM6IGuNN0bmGOlOfflzeZWiyGO06EmOwUeNbGrCXiUOFwJNaO
B27ZyrWNS8lNu6t/4I2cJhBcVgY+zb3UsBRKqUjskJFFodIppdZC2khQtW5EaH+teuSMSIvnQnzk
63OtNM6donoY5uaA3+xsk1D5CfEplT/EsZHkggWWRoavF2uHSN3oqPKwkvKw9Zc/e4NyQYTU3sfl
/r6kx+rb6O8SjbjiFWXRT/c/c/H+M7QkNU9IGmblZLicM1Y9Na1DsBS3QmUeOUM/eO6Tr06B9LIS
68JNampONdnDgD9kMDhpRXmJQbGPgflMLuD2EBC7jT5ewY+IrKBfH7dUMNkhnDonusIyb54Cy+X9
Znj3QgULXc3XL/Zqf8f5Chp2wlWj51eAOTdJPmx7nW0w+JFQxVtpOVIYHeDyB1IfXz/OA2ojtqP6
GKkaTckyvHB5uhTOiSrf9yKgFJfAfnnxKOGepPZezad7YO04dE/qNo5Cz5MYekED2O0h2bzcdzSi
6wF0lgDu97CkwgDZRR6VaAGwBQ3LnrTp1s2fYVTazS0+DdMeS/9QUjedvK4ToO2OJWY0T4l6sq4l
J8Tgr7o01Rk2R4LkqFt/vST0hfEjLcnn5yN+UZbLdVaQIupDeRpcL3NPbiq1yR3L88HSgLTaAPNL
JK3pZmD3nlqepd1pyHRVvaQQ3ol4+PRT4WeXeOqDE+KdMBJSM4XA50qhmaTmuHt5+peJkEcBS/r5
ilRwIE1oH9kWNXrbeQhBx5DxtEy6X7ZDCX/6O+Ngc8FW2vcxpQEkIAFna38OiQV0UUTR4vEN/WAC
q5w/0xnEXQNLMMi5RQdjLZh3f0BcSsVMNyS1FYMfnrRltnG1cOJHQhgfwUwH4NIEjDkVNjWBQ//i
7ivpqhRKgg+NzDyaqRyhEFErmpsB+sng0T4LDaif+GGE+nOlR8iZQlyjrbqalGSt6cfNufPTd+VQ
YFziN4m8xi2E4ZtG0Bmw9xI0Jj2c3pxnQJ1ydA10/0GlL+Z/W90G07e1JmvBxNlY5qJCs++6LLrl
yDZ2m+JnwBzUNMcgofkVzd+j4icfy4k2AlMg8Abx8VwJoiVbmHq/EXi5EcNwGCbJJ+2UzDqmpA+Y
DIZLfcFPsrhu68DWq+Qa5EklTIX7TszAe97V4Tr5iApqKEgrELgwQljiKEqCsHcRzEmEPoeZIw0O
G0vNEiVrau3QfJCJFuAUimdSDrrk80bsBNjY/rHRHu9nkX/5nJpNq96V27lxhWQm6AdYCOFQKQWb
dAym3wj0LfomVBnBCUjBuDJwBNRDj9l7vOni/Zlo0qJ8ETDKwazJaD7WAfQqYWuPu3RxLThrt6qY
EJpWh4I75ngI0ES68YiV4wc9URfPgNxw9Eqx08Jjia74EUnQnp1KZSxIK5a8rsTdZepCrKEbNy0T
djTfofn2bSRzLmxltFNxP0SE6AGmOlhHzFvdu62HwSWVG2x2JsFoBNaLMf5pqfC5/UM0nqD8AXaU
Lg5yqxSSYCHVoM936qVv83ap4WnqV4ApMaC+CLcuqiSUwYSKEcuXMmiXdEkthW12GQHTaJRmY39Q
PtP930W1fJDfgUj3XFTEqNiYnHgrDfk1kFYtxEe1XqkzsN5jQHS45EdRLklqEPE1+ZokAIjkg/oR
O7I2YvmpM5rJ0HLnIa7kiij+rEvsNL154ogjPN+kDKB8nrsuT+kvrtQs7NupVest/qMuJ1BGGK5Y
jCLSlgpxsfDoOP56p5sZDcUMppkaOM7N4FX8BVtJ7npn7O+jyUr1C9Ulez1qWoEFmwfnJ5PvrFph
FO9imAI8j2iqbtBXkV2KPXECuwKQEGOR5WpTVLKaaMdoA4MGBSqHC0X6PFjJEKjbn1LUCVwYVOqZ
wd0r5svL9HV5X4DvTocBdF8Iet59aY1GhbHfZOMD4wTXX6Ug4i9mTU0J9TMEAY6gjIa1pj7zgI9X
DaRhF9SxaEOJprvxm+q00GXlW7MSxQfS7qvJZv9ybe5Y9mSS0+qzbg4FIPjRi+E/8mWw52l0YTLm
wqX5ge5nL6/oGjpdUUDkTzVmAXCAI2Qy474Kp+pgtAiDAHx7X1S2LtAakgPCdTEmKMdHtgtDM/A4
pn80hWk7QvSACyq87p/8MyCMzfqDFdXDfP+A9basAy2NTgplyW2TdRshs0tx39097YgnEsddb2Ea
vT3KEkno4MqSxOClUCpaBOavxrBTjsHUoox6AVZ2aQ6G/gbIt6um/h0zXzKY3Uf95SzVZhQHA0UB
prHxelUe5rRr47bjCrT6K7ef51CC3O6OdSEfhcGJfw1GYYxVBJCnO6qOQ1pxO9xLgAHEQ32Y0x4o
wstq4rkXTRyXPj5Hi9BSxkx+Ak5XNkmBb9wXNsv/LDj7BJV3KP31EYlzH7hz+XUEe0nXUDxXDWMu
NSTxMqUqgjQsJHwUny6XljdHM9qfjdYiZyLDMcVYAwso5QPfVBzFlBS3DLcHAlyrfSKD95QHmyAn
a6SzI92fD2qpFzs9WRSNRde+tM8/PswMZTZtxVFEo0a35EVn+w/dhnmBvpOR0a5Ohr3vS+Qtfzb8
hBsWwT7PDNCKchxSfTctV2iZlT3v9x1RRPzBXq5h3yEWK7d8FAF53GXhrkZ7kLGUlporbSlmJNhG
HVi4J4Y6LS/3zDRGJ9wVGTSiHkdnpamVJb6o2PhZJvyg86kJY8t4r+ZaX4aDdf+yIKTFtjWzIkDK
YXX0FM82kbVRIXTq4WTufbTAqX2TpoNmNPlaylfApth1+xX4gIa3+XEry2W5+jMlEhq9HsbQPF1j
iUS7gB+GhzNGs0xrQ+kHe7mb+ncak0OxM2QyzGzEPkkFVEd+mbYEx3XxgoDVHDFpYThGS5BdGxNd
zgMssJF75y+S+TKY8GsvtU3ZHoC85cn6UKVXkHVn7XYnvH+krc31UAVBPXRGPW4TdY8bkHslSIpi
kezYb8j08iR9CFVZvypxX8NQiSHA458L+XhYuAhsrqL067fsw/YoUEnjLM9bVwfSOlu1KHuDcSRS
aYjEWyo5zwbESnKgPC6Yow6L33VSflGOm2n7/umRt1BXpnOvWDQk3ooR0DPiCssEEEpRQax7EVLW
cF/I1DIXd4qnHzrw0X2EDx9z/Oq6xE4cfSnyWRVArxvv8vDmxItX47BdgD1aTWau84AwDTJzDOW0
SIS/tvyefxkxdBpPlNWU0juu1R7CFOYEyc44h19GiTPveKdXD/W2NVdOn8Wbbx3H6ZU9Un/txHlL
RdCPpUZWctguseZWvCbRrE+zhoRGgGRWkW4KpDNdYKRsGTq88wsycTIqPeFmswWO+d0bOWy9zelt
Y9sx7WQlveT/6sleA2UAsuY13MagyBvOIf/hlHNVxbKFA+RuhzZgg+SOBcbgu6UYjnbm4iGm1uBO
l6CVjFMeFfNaMUeL0cpvgPfzyh+AuUlrtpjPztJvkWCUMif5bvBt0PGp/6vUd2iAVvzHcehoSI45
1Dj/DRlRaieKC6ycvNV23nqhQFKrBxZasxjp12zZgKdQENHxKz1UQhOR2ywXbOoavBgMGbq/rXO7
Jh1P6w0T0oLwip0t7khB9HZSfX+7vxr8BwAtL4V3Y0+aSQrnUaEF88wuV6tSaZrq1qHXh5dvxjra
R7Cv42hC+6hSHpKXj3DgIUAZrusBzx5/+zyFJoPiV92m1g3cVe4m1oi6dbxv1E4F92Pm8FU4Y1xI
NE8jTnnH5VSp6UmbACHAFHPXufAKJeaSEHQxFanq0musU6UaD3Z/3lipiKcmat9R3vSe14jM258F
EWLbFGKo8yKSaoHhPgYSBudEU7ibJQ32vIPZMQFP5qDHJFl6jPJTlBVdX7eTgm+jiC2qAROkI/wl
4UgY5i6jU2NHsDr2ZGh8xQZvJd+pBb+5Myf3tlK13uoEWAgnYlF2b0q/6pWUpa23gGxBUrJOEadx
8pBQb0tkZQNVP/eLtbtpDRWF+HsdiCbtVpXkVbkV0oP7GWgP6FkPV0tPdswrmmMcvX0TT6SLWlW0
OIO/Z+25G1vWI0zcOjJ3w0IaIKKg7B49DK+s8pTNIfKK26DAjJf+OwNv2t0YIRjA0jdB+kSYsQ8+
ixN9oRzJhiNcuQA2bunP5D19HbJU2t0+ywswojGSA3pxrFpv5zsYbtFAHO5ZynS52VCSx/cnU/H7
qdqBczuIZdzH5UF2yW6qipBu9zT/yGkII9FSi/fJv5/gXRJVmIYWIRmFXE3x5uOj9IPFRCJgYpg4
SoupmhfyEOFPDgQMhKArOLSj+TK9UBU0WM/MamqmMnUcEdBUMzgyBHmEkAQoe0uZz7iyUIkgdfKP
+834QQGMjaDCexKYIhdkat29Yol0CofjgSbl0XuOggmvc/B/Lr2twPx6p7k82LE0DAzPXLw3CnU+
mWBXgfrbw5xXFx3Zjd1qu6n8QVFKPziv7pl2gzrpJWyOSScUwLNaPir3eOtJjoYcW9PtQ8Kbq5j0
ecib26vSkh8fVi2RYmlAiYmNlsLipP8vQ6qihWLSVgZ3GLzSH8Df7oL1fTi/fgEHBdyFHLERcde/
TgBa/SY2d8BGNKxdOaTZqz+3cl6y+seIPTakBBSS/9SEmo0yxm1G2I1T5o9D6t1ZkMs4Oyg5OPcv
TyHL1URjBMywT2qJ8WVvLo49lQxNss8uUplgNlxTtZuJqW5oZCkuUVUpGRYMGSWlFhXAGBULRXkm
GyEpowD1zIsGT5UTsDBsBGAMsYGXNq3A5UeAiOt8CaSRu41o7HVsuo/tCLeimc+5/T1vmRg05iyh
3zLMvGSNsWc66fpy3KvtGak+GIaZUSKq5nveUiU7Tjad1g6ME/unBUkFoasWRD7UK/eqiZ5kR4py
Smd+f9HGOIvklDFjDJXPBQuhWaBGXsQ7oHnS5t4DnbBtFUDhElie3Su5o0llLv6Rtej+N6jWuGih
JPM5qSVC06a+Jhk+pJayo4UC2883tDtmyd6Ce+f3fT21jQKSS0vcGXNV8u+USBgXuUoaukTFCqUY
WxOk32NXRRVWLRGhWm1wsUiQ0VV61X7SpdJuRFWBVlKmIMxHaqx8c2XEUiKNZ87PV+rusqwtRZAq
gxmLXwB63HO5F7Refv2X7hzbRFHLCZo16coDmL6P1LQpe5p+/UWxT/fbtzj2dteRIVDoaZDUh/rd
AHBNjjpc3LDxKW1QUYTq5MzE1sYkxrE4YfQTjcfEDV9FGfTMQvjPdBROuQIEEL5G5PaYTqujFYml
ksCDzJSSPoVEVQkoIyWUGsiFvKBjJm34aIFy12Rm67E2DCkDXCMkWAy7veBY/2g5Ohab6WCUomz1
is1aVLE48ZX+Z8lEhXDpb2TEEjpGQ8ZxLiaKVsMI+ZSrPoUjFdgllrQrMiJqHDPAdnNgnfPsL7dg
NycIxB0QxTi3UXSDOlHtIDv5vWuC/2qxxcECLjUEiLoU7nZhy2DRXn+looLco1ojSACHfb5kijJ5
MyhoHA/d6fJ+3kAIFGjvaE2lcHm0oLGQzL3W5M/9eytKM2XN5OiNjDR6c0dpxM9x8ka0EnY1QpVL
8ssK+M+5+HUyb+CRib/CbYi6Zk4ccQPmSS86DeIHcyTyFXoNfBNaGUeRJpKKUbMHRUuxqXBx/Mut
7XTIe4t5XP8fEdzTjj9Bng354ov/9yP6UPe8YO1uNZmj2XsjNKIIwfeA/svBZsgKqzWPuq4EwqCW
ldUirUYwJfFaVVRqP1fpXlQRYxbWQ8ZMgL+jDRcxCqjKbxgwV3NBQ7oEFpPUEhfpuAIkpEuvN6QE
eRyOT5T10oFT8wAcZKqf3/Y06r7pbui8GXoxuMb/cg3Xyz+P/lS4tu+3rsqrRS15P+cvcXaUk0Q4
OV5lTuoWtr2+V2Zs+/M+MNHzKwX2koyVI6aYhlPxovsq/z1QRW/x70g9nw6e36OKIh8vF7Wynb/h
8p1El5eATmSoBt85LNpXAz/UlwJEJPkrtYv1Wh3Tcom0vYVCERKVGSg/KKsu6XQmSVAcS+vLHs9C
UjsgrdPEuAJVqm3txG3n+sLXZ8BSee+iv8F5UNEwFd7Cg/SqJj2HAE9dgITEDPYHtIlzKcUXzRrQ
y4OJlU/v/GbidCIjQwHKNjNeM908oZXu8ayFl2NumySVZcvZ6IU9yMddxC5pdMiujeg7xBOL/1ut
nDTKxTtDQjV7xiLleoBtRkrrIEqJOLzP1LoU7SklTLlQAVfnjP0j0c8pSq1xp5IMQAEdTBAU91Xj
nKVoSVMnZAJkH/fwUCcZxQFkBZstPPDG8lNndUViAOgoBO1yETjNY5xB57rkehXuLiUHvfSD61xE
X6RW/52IzIgxXhy+FIs4VCoWaXNi4j/gKK5tq9Z+mhXqpo5Vbfji2KkOK97ilkcgrTotimJQy0hM
BEhgDqcvYZzHt0laqHwBBrOY2QtbErnKWFjnCFxbcuT8KiF8MU5sQQYTMi+4Al5p3M7WksctVUdc
4LLodJ5fwpgTgjdOlBnQkJAumpEiV/MQtt2V8XgFIDf+HIfCd8dVSTZOSNZ1ZBeWQoE8CgEyDr2Z
zvq7RpidXtyK1Lv7CCjCx1FZWMyyrnXjIcioGPTQUy6AVtTkoGCLx04gLJkK6fbDndRExrPy4aF0
bwxnQKf/ggltZlz1lnLJGN5wOvsrfRjkUkPLavOH3tOcEDChU/v1T4H2ldIzGi//ZxPb6J9TsS2d
epXv+t9bNLnN9qt0NQ8OHVThadas1hJXlqRSLsoxJMtcyinr2sdMkvvV23QtKBYVFtOQmqa257Mj
OhqpdMUY7RZZRRU1cgeRpbTW/LAdOK44gHEePiuOAaJyO7h4obTr0ereQGAOJG+izn7bJLbNHGpc
uJ5PG4wE8mZ57tlKBhUZYO2nhYEB9T6oQwU5Hy7DdbRss4uzyb1z8X/9UFaYVLKG9sbT7H/tQbJG
x3grteeFWwsBuOW50MbRCfejLC+OFcCHPiNzEeenqT0tB77MJtP2DyMXG6kUBYjeDvh7bGevdq+3
tP1AYLV0DtZTTHcEu5tuS2GZMVEiXKuaIJfPiZ+Llxft800XwCcvg1R57o1pugVyI2wXk5clQptm
x2wICdNkmievF2xf/PSpgDOnQcV8sJU5zNbS1I8rVq/mm096gbqzxka0VDfJIsq7phWzkbY9QWkv
oSl5evLsoPD/JI52wO9rm+QCx7oCCGIVR7cgIoi7JZco3oOEbtWDemNR4kseTiRzV5xN8jrkqp+7
YY5/aQ/JIqMOGv2qR8o7gvzBfWOs/HVoAMlvmr1lMojV74zuFvmpMQnwa3p8Z9bkR1CcaZp7pXl0
o4yX0Zl9loJK6TggEohUKsvorirpJNb8uXAAK+CnKZrRYWNR5aE/cPv/U287+nyqQb/HokTUHoFz
VuOSuz+jbIEzRAcsLSEyzjdE1pDKVgUPyfkxfWJK2x9sOBKLsvkhZ9Em5CL1FUVU7nO4mK2GPpi/
jLbFrV9/sNNc6VcV3EojEkT5r3jHDom9CCQsoSSQ5b68Wo7BYrHiLYC5mRGj0hVSl9i58NGOhBuu
1sEY63wWV1x8hR5eHkv0ZY7Ryjn5QxIlBZQ7y+MdBFAhqNR9/nsoAtwlv3xXZbvNropYWwhXWYJc
/xSyJ8qpxZLddjxbzceHl4c9njX/QnCI+9vH7NeVcb5UMg1cgD1BKcz6vjLhq9vMv996+FVP0Tjk
Maq69ThBrZb1jEvzC5V84weeSX9kSiiBfT472JAtyO1OIEaypoXAal2KsiRBF4VCw4DfRz55vf0X
+iDDu/yGpDQkO3/G6Y68ZFlRTNrD5sBP96KgjHWK/SWtNDo8SNN19RX6AV+Uonw0b3peLSxKgVsc
TKTvZx2OJrmOFMwoSH/gSVjBq7/yTPMNSebEtVbD9g5d1mpS0HR7+BtzSLr/QfPu9Jvvin882deZ
hTBPagp9NuHDYum+jV09mwS4aiGzokAQq2H9447ialNwgzG/3dHdVNPG/NhY0ulnzPxMiDxhXG4d
XxJEeFoU6jjhLP/pzymr1dWJc8H4818FIvdeYsIniiTAWF412acOwsw/V55vJQ39lnMEbSwFhGHV
LYVyGLR99UnwJxRAGHkRGr2PYFAG6KN6JozuVuKIerdi5SSMLCemaNGx06KDD9qLzDtVxqKk+Gmk
5dYoWWf/tx7+mn2jKCpRzTHn7h0VzxCxnUfvIibIWeljsxzmMW2sgb7wI3OFJ3mpexKHt3cxyOCN
jOxD3Vr+AVKYU4QLpIkCqP2muqW68hnVodBS7z7CK3KZ6TdO/00376nDEyc5AM5H5nRJTmltgucV
PBFSnYGIuLGMZ/3o8jEgqvQD5bwogRHjyr0iBofZ6n6U1slD36b3dgT40a8gpl2r3LOcW1Hs1+mS
PUKA6EgIk14MjS7VLDp+2rKxC6tH9qq8xglNfdR6Txc5hA/Rd8aOrQtc03uw1bUkJjAB9+WNU1oi
chZA9YWM8sv0UaFtxs54x/IMd89XU24ItJL3lQmkxk7QEBX1T6kluuqmYSSidVZ5ZCNqhYs33ORm
CHlvP5hyPIoQn3RlTtWHQ7eKx6ggbHhAbbDO+hanoYAwo270PYrAzfyHYcyN1tj591uYTKOx/p5t
Aatw8oV8x+JMWtioXYZNW1BpzzSahy3ADKCAq5MtSQfD/hGP0HddwdzcBQ58AFvW8396TVipL8N2
VLkXtJiE2c7IbV7+hUKnJKtqvQPyXR8c5kOYU1bIO05Bo7aJcZMB1bCgG9m22ZZQdRvV29Hy/yEX
IGx3rN9o9baJ/fr6hHbztSHUo5KI1E7KlgmzLL6jq/r79Szcib+F4MQpiwPnMGWu9kj63Z4BdEVR
O8fG6rtFWasCMJ5a5AhBAuAchKobaSAPVxuY8e28hY38ueU4rr7rIH+dxeF2+0pB7C+jcY+XpFGP
10KokDbJEoMGZy5Hzt7mzgojhMnrv26EePEEtlxJjDlLu7PBtC1pKkBpe6EjOZpf1INytkTiJwda
pUHqkouPBBg9Ib5LGG/aqxPh3w+wwdCF9mQufcupFcqwgLe8TTZCELlddrfIS6vDMDtE1jfQD0VV
C0hJUc8TGITJljPIFKMmulcmXXBi9EFxAFYGUCG2sufwWLpMS7+yvysk7GHAOGGQWMEY4d4UJqj8
KIv2N0zSYgb609ZO3GCjlRYad3GdUaOzap/5n44lBoPJI4eqi14WQ/S0EarhhKfRsluQ0fhm4ZR5
SohnRzHvetpvBmXRZ/5ryr8L+ktFxTQbmXMsvSegMcJCS6pM41LpBOe5fpBWT0mYbntnOJKyczCl
tLGys9+ENi8tKn5uT9e2CyO3GezX1qmU301+RtbHWSy3YBMgUnzZoIJDffR3flYNwYeKYlb3EQaL
cfwEMcf61vjUofIZoZv4ULQDA6JutrVWk4odfvBT5Q9p2wU7MZ59sl0uFmQBxG3WNOtBFoact61v
qknYdTYtTI0FWYYMOkBEwgMAbwL5USvuhoLdFfiS8y1tyaMFHV4YplNxVU5PcbBcFWhoHzeSxa4k
PXI0Zh06rI/ZAnDo05u6i+sd0fFU0tvf7NN+UD6czTfeYToy2lc5eva5B9QnFTfMdvmqkFfxqEZE
H9rlPNWzei8dZBU3TQW6KcDBYDOdWB0WBlb3HIfciiJ5L4U+6If2QnNwPMdv7h9UnHxAQuCQWnFq
RLeeWouYU1j9HnG7R6yAnBrymOQBKDz3UJN/jVp/si/bQ4SFdkXVScgLnkJTBi2s9WfoechLHAPN
IW4EM+b3hSTEx+jSWIiG0OZeBlg6VOv++LXnmlYYtZoyKn3YQSDdKLySRCYgDpXfbQVxoxUjBeQW
dU33WxZmxW92QpcKDx0fKGrHVF+q0OhtRJo9Je2NTEmOTdAMBXlHzBrwemWBVIlBWYfE4LHsOVYi
nCrPf53bTO+I2yixub7n+pjv56Vai32k13J5sIuadghleQ842PjHD3xWEO2OVhKJ2NWH3yGJo8mF
jmHvKNHKCFLSBX9zyiI4ZGl6B+UPwAnhpz09AauwWiqkIxX/cUJ6sNxTnsgWZI4jEE5lFVDUAH+U
akcv1YeajIEc80NcC/I2H/ykX8JL9eqA3jxjM+AAkgh8YLnlW+X/vF7mgJlRVG1EMDVBCXFoPAOm
vKXnw4tmUIrTO/QvX3qrgXjbav1IBhWjQQag3aOlxdqdDFWZpMSWJgyr6ZTmcrIRDPHrKYRLLHdk
pvoxgVDhx3M3uczU97LNgw+4L6KJD2DhtAHZ4JDC+O0gI/75tT1T5/8luVNLtts/Sk631R/n4Y6O
HJW+x8/P088WNP506Lxl8nMSbnBPS3oo0AOEq16IGpuns5Y3i6vIqiKKVCo1GdTnkt+QBF0E7YKx
VEzbnGtcrORjv1MEuQhk5tSbgygTiu0x8CtNuhAYp//9fN8gq0o2kjeKFLx7pf2C/oN23sg0Y3oE
Q0sIaMpZrakjjk5xOLRuG/HlFTnIhON05/acDEHARAB/C/9I6RrvH6HzfD/s6+GxxykL57f1Nw1k
lOgUtxSfSb3xF/dKwUALrF1HUc77cbsiUjClgYlEAkamJYbxYFRuWw+WdwgKhN2URABtcFBczm4m
S6gcZvOZyvHZxltk7DNrPJQvo1AzpbhE5/H3gENHU3X6ETeZDKGCtG1kUEsiPeL6YDDKb9oXh8Pt
sNXTm4yFrzN53KJYGzbHUs/prvwlUiYW9tT6MutZIMH57NLNZAG+3q9ZZWJ4KEmLC34xI71GXMUG
/Kv4TS1b4pmIid8nM1S6XyG/Cb9iZjeFhBpn+pzoBXz7sU/pY124bnQB1VdNC9CxFphwHrYvcjvE
bzVbhutizXv2lLr/5ZzQgh3ZuyZDVDyehI6Md1S1kT9xQXVLPNFUSOiuqHnqO+xMCAepg7D3GeCE
OStLIhbpI1f8gY1O3OT/NDelgkbDaxsmKm0iToLVz6Ebp3NgJW6MdH1cZ9xDlZxpZBr/BxW46god
67RdzmtWSZxWDwj04/M5FIEIx2dcnNZK6w44jG0A8h1eOWkeGksPWGRFRmxxuTfx1b5CykHzO8k6
3YFtwxBsgqGzRgZahu5Ul7MdfD82Ibs6LE62YuHh6BzHwe2UChypvS2TijYy9IBUHLDYt5vWl6ss
dmCh/xqtb0icjG2QnrmGuO6usQ8S+olkk0npWEmoXGv3975JDX24+N92xM/0e3jVhZNbLvu+SOap
uZtrs2G1Nd0K3m9DPou18e1Sn1ch7rv8ZhufMb5ZakHafRIaePiLO+4+9WOdqWHyHZenVx8YjJA+
VgXO/4dSOZpn/c82HGQkNiPaAL77ayUVwhOXQe2kS0XpYWBgrIhLgqnCzmd7T3FJPtDuDGhnkOLJ
h2ZF/KnkjxiHGyIgrfnADd9V11PqfFkhyi76pwijxxS2zPUpsmtEhFwqMGc6eo+O4KWf7wJaU/QI
mbHfCKtBADoDJg6tYRq6WmJD6tBNq5/1cC0wfA+edQugwWW76Nw3IqMOGNQocop0AJ0Br5gwhE5d
1/YbBM5/5irJO+lSQK8I2CdwzZvVN1GbHrH4hDvd5GjtLDV0J+HVG3FHM7+no8A5xW2ZYfigOx6x
tRITrB3KjgnVcpQyCkx/o8zuVqq+xSLnnYPPea3MPCfA0c2zfz4Qe2wIFdWTuEMXKd3IZOq/0/TR
gQzd2UEzWeBZtFLxCvKfoOVEsWMAH+H/PUMUG00sjg+2T2QQ/D3EN/p0SSWFmpWWHRkz1CWWKBjQ
iuhyD4DdB4z+UW57U64p/a8Bddbxp707+wUgr7ctNdbDhpJyMj60qHpAyRjcO3acKcGfSwor5C7D
m3Tnij2Qk5HggXnDoDs0On/NWB98CEpg6U2DEVU3Z7cVelWR84NFScN8Pob2ffHuOxOMj2fG+4Dt
7ou6leQzJWLFPmh+/LPGEeDM7fTibNDY50T/A7jkydejauZ8I9o0cOfch0LtxIT0aga4kPpcMYg8
HpjtF92B7pPIHUOrlMg8ArgmawrIPWy1WtEmbIVdt6+v1SFZNqHHvTZiJiSZ7tAfk7hookDSeveG
jXwtkaL9HNYdgtlgYkN4JFo6QJxCoRP9Uv2iKCn1U0FSmlQkc0yxJ81mdNtZEmJvFJRZIgCUoOw5
FD+9ZzmROArEBF7WNJouiPpyIQS7wOnpMrC64N2bIt7OZzMh/FMDz0T1XjiD4bTBPulHREao94tX
VSeLMru2DK4rD34qmSrJB/wYEq3LWQghm5x9kFnn7X5RyuTseY0Ud5tsLFVopR3fxrMeCtAs2l5V
bbKxAseIrvDkmvTqWY5XNVhnt1RZ9eMCfq64HvhlWyE+gHuNEwXY8b1qrSiF6zO7yFqrvU15TtuR
GmPQ1TWKktWTMgQhYsF7hAIyVyiXJqIrCPkCxd4ke/uMEuJ4Z83jozV0DHJtHGX/OQjtVu8CnQ/A
1seiJqHkwau+IjHBddqP+Jw/4GKBpd+hLQYWQCv4oTR1k3gpXMF/khkFNIbDrOXhrLYoRkfwlaJY
DdN1wHMUu3LsGR2bUHVM5kHAhJlTTrNgLP4ejF5cM/TySWLOd4rnPokF4AE9/lPg3tg5cLR7svOh
Ilxdz3bdJ/MNxJ+FM/MXdI+tAkGu9RrDbZRvGmIGDumN/Y+IWQs4wuCSJm2g7qv6q6FCD2n/G7Nw
qw90EviZ+n/6H+JTg5HW9UOPmJORefPApsHs6CAwJERouIAJoC5stHs5Pxfr/MVwBNJsJOtTXyRK
tmsmn7+iGZyraW/0aH9j/mNT7+HPB7z4882gF11YsyI0mIZX5YPbGYEV/qURVnNwqWQmk0ppKtN4
/OaEz0GUxpTtiKRRSCnE3f+B40NjpDBZJ4r/rPk/YyXwZr+42fIsAHhCnIWrHCm+FFVpp0+mDNa0
+bWNpNEkfvz/6oyx9YIYFKeddQ6lxqpEVJCqXdWqrpYRQhaYrlqASqg3xWpP57oWZPj76m8SzEHJ
BPyztYLR4pWv65oZgRwY2qwKPxTlwUYcglYdqm22h3sMSBXysNTVxKCZjtH/f2Gi8/gczpQN4Fmo
Ta3Gq0j3t7hRipQ+b7py3WjB3/ZrjATSSY+PTVrL/EIC535385HZEN5bprKvGTv1SJHzNhvzWSg9
tgyd6bAMaPtyttbE7zTqG/yNDmtFqLlqXs4GkB1wllizrQbBcXVbcFT/4QIWU+kVDwtsb0qj9UTG
Def+6BBy4P/tb7ju+Yzd11hOHcGlr/4rg1czznp9FSeFKdHopkwwA19/T1jbYkj+8Dl+u4gbKfSi
5T57f+SDVdGQezlq374R01nsyXuz/+zLCJrBltZU9PKqdcYBb8Fw1OVPnCbZHKWaNJQQHdC9nTun
fnhxar834paWJIPX9RXY8MOvevpeI6EW44QKWEVVmmnjND93vMBX3kPc49uWG6iNPIOCzIHCSqYw
ffVpyCdWDQyUyLobwFhiaFdqyXB8atzVTrTgoaF9TxpX3XZlYaHSfCRf6KJ5goPNQZACpXRLFZvy
ZwjNnvo6sKflXKH3tRfAoSiYYyiMfceNR831i4qaXxaE1qWQLHPF8HhB43HNVn2u/uJ6WTurEo31
nyJkV+uSafI/N0Oh6qgBc6msT8o/PhuAaKHrML+ZBwA5MvtsM5Uqe8kkHbnS4x9ZAtKA2N+BYzwB
WDYdKoHtZyMaAbTriwHXI/M8/Po5zSXQuptJTA7RleL+enuzhVdVws70VMBOt/oSkc/4KeGx8FWr
nNWPWiu4C9cdDV3kC7qPxP8FHfQ6K6e8tkG/VhKV3LLla7JF1hZUmaWRTPxvIF7P1v3aUK0O9AUC
h6AH1arb8z2qLYUNC3jzcIPRPy5px3fHS5Q9XGM5P/7374Cw2DkjYcXF3PEjkoumJvWXp1qFlhka
y2nX6wUvNA99lPLg2QGqKliSPYV1AUALEDXcLBN6wpbhxE4fGqxRlkf0hXw+Mj3iCPV9rMTM4Byf
Xs02q51pT5rhdg8SXgXNu9FVADpr140TiGBQaAr7ITIaPbfCGvwKsySmH8bS81QF/sF/LMA+IouN
4VVuNiBrfrwopDn6TdPiGr4DfFOnTdvqLBXHAxA5O2HlcHjR6EhZeitlQ26u/1JTRlhJTx/qP5Rq
xo5V2qLcLLTx2jJhuO8zUvE3B9npQVog24GI26qEYOuPceGoTrBtdqmcLBkP2AceFl4qe8ZDa8ZL
0LjorV1LR5ldrycJNcQqnAjK1xdeIj/kdbAz5cP8A9R8j1HNxEgQ6wlrt3pXo4rTiN80LGJDCbrr
P2d6wVSokAdLPlpN4IJQY7G8Qd/CPL8sFtFpxC1aqCP2ju1t+avO+JLQJ+HbKTbxJgGKHW4VZBZc
XhFYM4B/zUMCIQ50iUZ049rfDEo6qZKNNELvt6xD8jrnXFSgWd7KAGGP67I7NINrb4pKmGPlQMiS
YJLW1AjmW6uxZuTyciFJP4NWgb4VvHKS3eSvCzAL7mzLJ+aqljvbFcOs1JuVFQ4DShKb9J0MT8Ci
PEMaCR4204o66O5IP2pwyNe+H747QUDHxgfR2j+97rBWwCKIYt9SDkLNVlu0wWs+LDHl7aPKCNk5
PSUaINA05Z9LXW7MWQgNpXLw6jl8CNfTEDCluuh4KU0kh+l2yrCGlsxOdTalNZF176HRqx4els2c
Sh3iwLYveqMrB9jDLCZ0/MOmpEMZwnGq34AYYYkCJWaKrtm0oSvcO5JzjFCMaKHxEkuPZQQzCToK
n0cDCch7UUuqRTyiM6crMOSXjv8W00zUXwwr/hmWRuXFUu4IE78BdQalJpLnBk5H3ePA+qyu1u/I
hrQSVA0kQZI+VWhIVHnk81xJD+HLPb/33Gc3NGLp+7nr1E/kRQz7xh6DRk55oEkH2hzBcp0CGmwZ
acaNsDlqCwoICalmJn6JF1NOkYQxoXUoNGdoDpImPHAZEnQGJj6OGmgvCDz3fetaX+a6mvy9cLsb
/w5cQwXYXjYx+HxH5F5YbU1v95+Md/7TNfWCRvjhVA243JidE4L6rv/cu7mteZ2HW1EjKuntqc6T
aGq6DDe3fSiahF27WUU9g8dMkTln5L/RLUMxDeXnjf/HkZdsVhB7P8ELrywu8qSACsJgvMLdPbGr
iWamHfwrwTiln4pYGoswM0v1ab6eGYLSs2lZXsF5ggO3hknoxiId6yXD2SI6dh8xzvgFyYLlW8ML
KjVRGSAJANfYRoP727v12siwWxaZMQL9/tNEDJZVzDvAy8JfNQXPVOUQ49xKuE8MuPNuRYUfhG5A
lGFEOgeJK6Yg1fm7lrsHOsEfeF0su19ygt4JyvxHvtY5IKeYT5YCUm8ioxzSqXDvh5AQ8eU/YLPP
9YwiCG1XG1RjomccEQfliPOAgXPsfljOq57dwaXD3JnNfpdgppToDNHHev2f40d/AVaYqdp7kYJK
7+tEWqK0ppto3e4kCyJf5CTkeg7fnl9ZwKEVHzSP69SvvnJ6ztIaJuV8AjTLniRMxqNULGlwfzJt
9au57OghCjnEi4LgkdcseeXVi2MGK/KNPUODroyi3NnrHCb8iXsujJqGkf7jrHJw4NaG7xfsto5Y
UgBC5n7Ivue5510Xo1/69HVKjUAiy6Q46R408XRnSnSecFMY2mrvoyGB+6chtwDj0F74zPo/d/eo
apYxzHKTKDJwaPRDeK4oaMoc6ZPmwX20COssR5pRnxUPp+0ti0B5LAf4qlP/6m2F1ZkSdfZDD1HA
Gtx8nah9GE7VFhKN1LZeluRXAXuajxnVxxIYbkMr9dyEZ+dHoG0FhUFUcOOyOGVYrN01f/JDQKDS
GVOcFNHnN8xYVZpqV10aBU3EbjTEdwEvriDleLrKc61yuxnuAoPJ2pnhP/nw1Iv6gFclT57Xr176
CMWtKW0kzZy6FnEG83FCFtDcwMyHI+EbNT7EomFMso7z+ctr6GHykqe7WTcVHwR0npw41I5iu8lD
kgUkQPNxTpW51O/UN1wieQcyMtLMYWSjSVzHJrYB2z0xbRqcbK/uoM/XcysPSWfY2F+tHZy4/8ov
02G1Nfk1tVLjBFlSIrvcCaq1RKgdv61w+ur9AXChwth+qwmO/YhC+vXqY4ZT8ex1f+YnbTelkoHi
QE9KdV1zOfMFN0tt/gNUIg03vZrSW9idgkGaBwk/JpuqxwM1+8TfR7wJxdNiODgB0H0Nbn8qn0Y2
RXXtvmmknuJoixFhg2wNXc7/0Bvph4T4Oj5CuJEli3vw1y4svXDQSRNAk9T9agHsqQnhvNmEPd/o
34OjOXBXc3uIZeds40AteRubBAluYbyXSZLZCLNFNDYFrbU7RDu+CzkTaQ1FFdXkn1JziVTQHu+R
LIgZIwV6DDNYnzlCD08fr8nBQsxzNP37U0DT9v8cNzCBVKaW4EfsPa30yaxOfjgtXBg+VlizQYEe
in2/q1NQy6K17evuxwsI5NfrzyMeZHlu8NUJQwhNPwt1IyhaOVOsb+Pv5POkVQYpGTvSkwALdjvW
rw3Cq7wMq8aDAD2l3dE1iHOR9FXHDPVctCQ09qZA7HmyYxlxoWi1fzDcMdUMEuGRLCiAWeyVxY9R
YM0i6pY9/uTIU3YY8h5MpAzv2TvM0q/xESnQ7nvVG2ZRzz3TI2PXzOGf6Mipd4x8fS6tQ5Fq0iDf
gd0IV/Ml2ZOhC9ioPt8x5A5dVgwo5/OnKSoqHONVWSX6gdMcvj0nesTW/s9XKkjdA8u06wTvJBxQ
M2LmYDu9Jh5RmAXw4m/qfROMkLR3CKz5UH3y7Kub1wYp5p01nIcedHbr1Aee1hWaYFqS4nzqQSbk
jvndIUwGPBVjVwZ9c5kqkJws2bkENR7q2wCCcY+woBHPdCeLThFcPf4wIrLe/FvPVgwCnwYD9Uxw
JNi2SngytW5ENrCreBZkEAO7gTGesQdy6b4/CC8QtS5zGbys8Ycl90AwkwF/wtB6lBc/ra2rQMyy
TIranaT618IMjBIT8z0anQIbEWohupIms+Yn6NFqGGEDlFZgVDlDYiGI4seqj+lDPkELITO7GYH1
YzmI1QykyvDcojsTJy54BzPa5eHiYUHXXr0mDi5Z1wt0gZ9Gik7dB1Tx2tq7O9qAjK1m3MX9ocfq
nkGB/ZUVb4UkFUYz2v+w2od7VPzeRlkl0RLxA5zEirjeVBC+WhJrCaBPypVgGnVoDiqT9P4MfAp/
I4s+MLULK8J04i4FdHcyWmz7bIK5Tll27bThoWsbw4N+McO38t+QkP3Rc0dRtp8HqnzSeBcnGTDy
vET0chqQm9InWIePPwissN1xisb8jryvD1PkZi20oceKMu8qh42OSIf11np6qd8SlDercMOIC3rs
OXjjNV+yXqagB0cJSpxkPh/dnphJDPYAQo90mTsdYt48mypyGIVWweVHhIz1LcoLE/3hK8YZYla5
trmBtsSB9JaHhDIT6F/yidxoYJxAoDloeLLesd/K0FbY/i2AmPvblLRWZBCRB+fta0PbY67vGXgM
j5ibk9cxlDauBG3hAvyR0SX/dBLGXbLh0VKkfOf0LATkifMc9CjvDwUy14ADeHQbaQ24v9MraaJw
xHpeF8wlDQq0MeKdjm/oZ58f4W3wvZ8QgiEyLs5IPzbM7i3OJGODswuNam3nOTtBL/YzzCWGKf1i
s7LabOplRM5EgISa3YgPFZzyuoIP/6NXAhPtMHNODxZ1I9HNBCB6oyrbAkKsP6M8JNJsh8QS/gYI
+jVI8u3dLQH16edjQ8KlGzZVwsN6/fvFwXiKg/7vdzQkDbX+WXXvKr+9SxmGio9ZxrS1b/YREbMd
goFDLxkTGwPriI5o41N/wmE4VP+gsTyBPtpVTtNR0gnEozrtNRUrHvvdcOCGaw8NcxgbiRw5St3C
nXVmCf3mTtWmx/kwjA7zLNqVuuxjG44HvR8Ulm5N7qtFp/yHeAgiTLtL81bsx2RAwNdwoOJhJlF2
YZWzDU/CyZjDZf1mYatvr8smOK1R+xzRUvJ4RTXM1rRSQAGYJeSX9h2yGM/DVTRpeCUTK6BoirvZ
qAksle6PpVELSqDUY0Ilvr0lLzgy8/nMeXYV3u771kyzZEt0W5/9mrmKKOd8356QhFjDzMlJVevw
XYha+NCMnj5PvuIBm8q7pyU8pzb6JLM4qjE69M2qST1J25y0A4AQcrh+HMStqUd3aSCKwgtO5lN3
xArLGZDYBa3htNnG75KSGsRVgILFoZj6f8dIOFjEtnlu9bsVx1+7GtCmw+818GfLpil8cYjh6N8N
nwQSRGYwdr59TkbsFG+mQyOQbHmQbcLKmyXKgEvGA/IYXCMxVVYlb3nOqgRUdJh+cJnY3CQpKuD/
lOKUDiE5xJfTqNjEDLljEf/etNAq7f2EE/NNI7p306/Gg+K3Bb/hrvM8bhI7QTPWUJQ4CzzpBq0l
kdw0sTPZWxL/PNOe1vZJY5+5NLrGuwRgwcCkEUczSrLSBNaKgaU/x6OZjzy7Q2RzTxbxXKVKtR+X
L+PWGp9RzAbu/CJuguME+Zo84/E0GjYQlT3QYw8jeaL6f2206WUPVC1eUnG+wW4J0rEMItPMBJgG
v3WlcPbiW3XHygIwpMeJTbF3AwsW0fcbeMGQoOBDE5jnxjIjGiHti5lspLd9OQ10MTlgforTmZ1Q
mO0wI6xshyHwEK7CfG+fIRUswOde20BQri5qGC8TL3EXRNnLrIP/OZbvayTZe52GJWgv60MLbtu4
HGLd3oB8ZE3BGe0QzUTaAfsFFrnsV/byLGbA18ZhkWKsmGmZepfg0mNcFuDJmFOa5Gd2CWVxuODH
1Ty7/IDbt99spvv4GroMgiGcyudo8gWqPhqNet31ronUWjFmBntfIMhxxtANdz5RAR4jvPmoiKk0
0SKc9KFG91y6cXlzj1EGaTOI0n3Qp/1ircGBaNz0zC/51sbMIeVfUNUDXOV0xseSYfgg/mDaBOql
b+i3XpGYR0qz0zUzrWUaKpp+n/McjyOx/CXqAgXlR5vIyU+psVito41LAFGD1DEcF3uiauVZJci6
vd+JkyERjHiyS56WTRO2XDDI/E63vy97sW3euoziDIJUwlVc2ehTUdtZ6BvMofNMnPPO5/dNqhNj
GZAtK1xfH++7CZUmb6IM5ffX42bkPUfx9qlR0YeXoQsUVNcjIa8d3DNcBz5NcHAj87XdlVqRRrT5
NqUnIQl3Xx3EWZb7DFzfIHfMZDjx5aP8aY8QUxs0XAI7dIiwbZ0Nuwecv7INwm0y1WpA7HKKBW0A
t1N0dsYaX6LvDaoa2LYeTKSpc4jqVvdQkPFfnLR4NiwWNbiZFk1wOiY482YXx9LWP1g/Ig4io0OC
OiH1n6r/iJ9Fv0ZSQPbLtd+sj44yOqbqb8YKXWY1hBJd7yUONpAXQ4GQuih0ZsFeu0kGOb6lq5ps
XerYEqHoLaBxW4Ahpy7gf0EYqg+cBHrcWM/AyQTD4vX3dQnzjc7iqjZcevnWd3FPToEW3AFqhCuA
la6Hx6OrhfdLdiecgzCcwwKbjYqBZdRCGELUmFWgdgg4WVUMtVxCxxv+8AafxW2MBdDUzC9CogK5
ebRiR1ALyXEzfRef1CJ8ZCJOGszUfzOX2C+CvfFNb9VIyRcGxw8uFsfvJk66tRjYpg7qrRIWdZJ+
RMnynkJxjcueyf7+V4E74/pceiyfdNjNay0CgBXUn7Pmd71gjqqrvXeyRoDzXn/CF5v9WbmSxcNU
25wdKhD5dyb2KJJb99TqfaxjEf+DAYgRou+zRd5/pl87mjJbiHixYcZhaqNQ1BhMfA2beoaGSPy7
KGopgOy2fVSTkxGSdXg9kKFPO0tRcL+g0fqqKRd8zjtjaz4JbOMVpn8DIQ4JlVUuBMOr37bbh3+5
1kgRmonx16EvHo0bJsDcZlROfQ/Z4aP800oU8zSBc6lz/u/Rg24vJmv91wnD7Fv7zwV7n6JzoGKW
SEHhGvXjvErwk/hyCTXag4ASlFlcf2wQ1UiFwTil8FERVITM2GiX76LkKK7PEDKY4Qs+u0oqrDah
2v3NVn2A10mlGVzfEGQB87cwxDftIWmonoQFAsKEKEdkDmVQKk46elnz8QCZ9lKr/H8gNfeTIOPv
mpGDx1EBerNI+W+Btl9g61YPaw2XKUbYj3IAwmMAmYG+q3tDEqdJA0px3WnVwDr9Z+tL2Iok919m
SQIqFnTcL6CeH45BcUulD1qllPPl2lQ1VLdNN8XBuGGAezdaLhdtkU/uDgzi+XxvLLm7XKgzeNJF
5z3Mgi3upv/4o6IxuSB6Dd+zck3IQ3U6XiuAn1OGmyH3mgDWfsIWJpVrQXmqka7b1jUAKU5zzHWz
GWuLtd7RYRnTUEKfobV1gtHwH7iZdCL1s5qpQX1jbsM3enY/QjetPnUFP5whYIMFKZjx57hrHB+z
7Ijkuo7M4/saiFvZBY8/J0XGCfdzVlhjNGSHskMJJRhQ8h4bZ3gnHYoOfjDaZ7D8SR3qiLEB68sA
zoLAPnIAT3J67pdmD6Y4HFKQO+jd+sW4lodUG+VjeyMKM1RYmOgTVVjj1c+ep1V39uzi3Dffen6N
y72+mdFAF6pNXav4T0NomrxMystV1Rh9jIlI0TEZfD8BFxiFGAj6LPMFYJ8xiCxFq2/QF97WOQaP
PMcXbt03yuMi22f/iK7s/U55BUSV35SZBPd45MfvlI9zR4fGrenVVa5zHAUCXdErOpmRDVHrwDN9
9jZ24yAOR+1BR2AGRC25cl8P+xKV4gMNtYzo2kkUq6NADQFJ6c7AbnkKkDcyQtyT1yjfouoVkN0Z
42lktgTfl7mNdOykbIt3bGN9/MM8TABUE3/2TGLgx8nA9DSmqTNSb2YQvIuM1alM1nj15xo5o/Mn
pZAK6Can/6fay1oFwItE95fKPi0f21ICXbvLPct4aEFEIZx+otReQbKQj3kf9sgYQ84Hf2akxAtO
IiBlKIRWIczT4AouaV+qP3tP4FqaaDRMsRHMckYO38PBA7KKMwMcHwGK+x+LaEWnKlRbo0S+z7sp
TQmszR1Z+YwV65a77vgdnfHq7P6HUcUKIm7eQ+5WUtgG2TPSrYs10mFgFMICUh8Q4MyCGZGI1eVt
rL0/lXQbdSu+rxFfsz4l0FjpWMtk9idtjWGbbBeap889s//cXynpmAHZwqsft4IfJZLIFNwxsQcU
PHKwE9IBhIBUIWwKZ6aTs9SuBaam40miLRZMq+RWcZsui3EWraISS1fs9OPcbafKNtQv2YtHxu8A
hEOE9H0E2d4+6j0mmT+nNECP9HVahvPoi1dVQcdvPmwyvRedG5ml2oMmRu51Bko9pkCTmVDVrru3
/+ffyviuQ5oRONHqi9G8gmurvMpMBkwc7uoUeQLUMv4u1d4J4k61XImtzrHcr+l40zHQ6zrxaESL
W4zpM7Yp7+Zww/xvJiNpBK0u5yMKlkMfQnJh1RHH5I/Ovgb931XJQD2d2chioFHC08EOThkKtY7g
kX+hNwGHzqMGTFMpLzJrzMtGW6jrIlweLkXb9GDDPE6ZerHLRImXw6buSLsIUDaUhVaIb8W5ah+0
fHpFhA4BNlbpxukKHOXgxPgkLsfXL3rA1SqdUYXAJsKhNXUVNYQ7z9gnT5BIiK607kOM7Sxb9o1F
r86Pla5/H4efQAC9IT+1zbG7+SycUJJ2O0UJfAUaBGeR3KhzqI6FmL9Zr9vSgGQtWvUPj/DbjOPp
jGOIC2QQjBeIddZT4royf0zuYZRA0xNPkO0KD5QdI3R3NscMsOkLRYMWEDPPt/rktbCiVwN2mkhE
RHhxTh9bnbO+XJwgyG/XgZ9jqHPl1iMyLIphOAp3yBixL9h0wBIfumT77qHRL/lNLHqznhQpFViB
lMy9EHC0st/9Va5fcYw+BtCPO1D/GvObYzazt8uXuSZtO6sPnaVOBwLL2yaDvNHtxW/7IYiB0Bxj
8FodfOdVWp+bW9/ShuHx4YrmZRHPac6hhdSWd5hVUv4bO0nEOu0+f5XAQt2c0L3GaVwQ6G+jPJIq
1H1WlK+vDyG6yPalFz5CRyswk6iaZBJuARDPjsj/GQEI/qSZCA0Ics3g+PozozrdF+w4MZ7MYGiB
FJMI5fupUDcHwSQFL/D+84q3+X+GgVym3DuDS+pYKXdNjAF7lbRXuc9qncMGyEBEEc2sjGkpfLPY
wvZUn0m4AdbDbKAAjL8yfekOhWBLi3yqsOltZdoI5hxbM41EaZYWvcGcsU5NtsHkI0kvJHZlx34d
FGmi1tqcDVBQzetabZ4QuU6AL3Tm9z8+p9//hidO2hZScjP8SWNbPeCjojOaf3NiAn4v2YuxlLMZ
u8Ara/mswNg1NMUIuqTQtGLF2+7yZt1NMvpEAhcjkEdNIFNWYad2ZGgU9WPedbDpTBWDZCq+fvMi
7mZsiOgvCW42L6BtIRawGRyF+/Jc/shI/a+z8s5LVyMz0MtHYSVW9+kmYLFbzPjmx+v3JnX5m1oH
pTkCg41rto16L8KiTBj3/FNNYrmqa2cr2RUb/8eL+w+j9x2WUnxp7ucJuehzr6rD7IUEYvSnzO4W
/irLr+bc+kgoT2x808SlhhQgFRcCHcQK7JImY6GTq4587EVulEIlNKDUYw1tTkCeWXh3tOGr71/g
SQTa+PVAmapmWeWXN3giN5XdiLORbhYEFWQ94rCZAELIE3iSLqX/tjLd1fyC/wjN0cvWEEUZBs8e
TQxDiq8PRsoGS8r2EkKVeKFVCDoHPaf04niHJO1scm5KG09vCzTidfuoYuiEcSzjJTQVEfqa+pjr
hwwyGn1zBKjp7xF9NIIJ2ervZelbphgoiqT/5xGILEivE050PZsyYIUwPnts0rPsgudxCzQ7Ozhy
5aTU7WT2bmxoB0neM/8ZiU1fIdFjuwjePe+TIsS72jzKLo8GwePLvQ7o+n4qAtegsWqdXGfQbOzr
I7OpZ8mhmcT5inUqnhfMQDeBQ9eRO7RXSVZ9Ggp9PvQ5c9fNe4PPwp5E2ZycOinS8Od2jEtaAVgM
FFwaEVQuztAZQJ6BpZk5QJax8rihJOvzBD6yYj7IYFja7ONK0bSFTO2vSGFDY5eM3zNgW0sKlcOz
z4ox8oo4wL7UPZJj9jtmvJY/GnGChzUHqCvPr6FrpKUWQm9nq/VFBdHh1lcfhA1aWyFuo4OXGNPd
5OQwcAhU5sE6UpmzwRVN8xDMMxA2CBTmSW2HWrF5BrVCtPNCGakwSzTjAK4YWZMX/B9HwZg/bJv7
pNcM/DSIvjlBZfiQ5PWHGyLT3oJ8/a2sM3UkDEjwMl5L4yRGKbxPgm8UYu1Xkboew2vgEvEF0m98
88uS8D5pz4JS+feWszL2VbVNATCSSRC8kolSK9cTwL2Kan64zycVFKAce56NkiCCn5CW/SFvuVn3
83XuLTxnQ0jM7fN1dXN1MMEwlHtalEXNyrEmrBgXiYWfyrUAaEPetQbvbmTPkFOABaONN3hlKrYI
UIOrZ25U3ElJnksMOYn9kHPgqDagQRRYFTE5GNhOXLgc6mAZkHErV5a+mfPVcJiG3PzOlW80oAeG
zyzyGhAQLkcvopwc5f1023w/NtX/Oswj5bIclg1K1e/ReR8kyOXQZhtGYugn8tR9oze/OCYHtkV3
IImiQF4mW2+mvlwEiOreIJzzL1y2FEqTKBOmGsuzJtACpwMuOXhyYBHhmDZw5c4OSMfaB4jz51AU
XiD66BxYou2X6QuutOJtyzlFDd0aw1RzGCRCmDuCrD5yTTkhT+3o+/cuRTHbowXbMKhvKScX6ka3
43JQy26UKguLpwJmI+mmO58Z4UW4KdgVSjFUcihc3z7LebhJ5mcXVXG94nzvrH/uh5uyYICRRqyZ
oCZQNfpdpXn6uzVLh3NLvsPX/cD9mkUCbBU8ZIWFJZMpePrBSaC5/P7SHvhMlCw8oAJ77La9sIGM
62PjlSdkVAplFdvbMVoQ8hYDxCogL4YgUPYnwvXzMh9WSh8K/eF8JKnujaUF8lhnybHHKmLzRPac
xi1fsfR6qXRJNmXQxV92rzurHrlRbzuXIBrwej1YFUz90jR3DUdtl27dxQqWB+QtePJG2UMRK4Oe
7ofwSKxwVCTrkrINSKCb1x/VNZNUopZkE/tqN2De5NOvTdM6bhgxVd6dfZ2nD06lo0JU6R/BIhh+
pQ5UinNBuS9QIxF1DGiqaGwH5PFrJtRURWD7OgprVwdtmYuh6jPA4GjmG/or5RBEf6Eos26TpNNH
J14PCW6dqb6yf6OtJKZaDnpYjMkqnt1HKXEHQVn1nJk2cqgVMZIaZFqbxBU/MIjqTLrwmfT32Pyq
a7wGJboJtdkDKPrVNMPk3/qzIO5rmuM6unbDJFyzvI03skl6Ui7Zk+edx+6mL8K0hGHTNyxYX7GP
hyQJhLXOa3Krm349t9bRl3tpJLbPiJy1Bk4FCEzPkc3Xylk7vu2PQn6PcZbMbVGF4xBGBNeoZ9vg
K3LdvAx1I05KbJIkHFtnXp7uqX0oSQHFESMd2kCwz78ERe8VmfodVsPhMO9y5WX3oS23UGAJCiDI
xB9Ryk32vxEBwKbCCCpgqN0jSYJkIvc8zdQOEC6HjOGvalcevgNY7E4P+iNlOiufgwoK0I2APcXk
GBSv6rHj4dcprWQVxHPhrE4J7WhBPEHrpRuj0fsrWRuZAN2f4uvLPJ12rJB6syR/PwKampvwo8v1
hoghh3fYLyLafF/BVc3wjtm9HLsTyIVsK2yU5K+tjqzQlL2vZQyYbHy9FpHM3kUF2JHAYKJDQgI0
jARolQIBOQzHrrIHRNe8TU18QqZCuwCkfOLlKRy0YjW0UWi/zJ1ihDUJVMt3dSRe8U2DKNu9jtx+
UxDpnw8u5bn8lNc6dKrtR/OSjNjx2OrTTbvdt0bAq9ZluMtJyAJUDYd8LjuKvNsfJjSe3AF29D8y
NgHk9W5ZwA+jrh0/tMqmFFRrO2WWl5OHhPE9yGKQWXR8im5N7JNHpdzAcT5gZgurECxpANnM9J+k
gUISYTKTyC65jEDaDgCCoImGAXqUnFxgVX4DY52dM/gbBK18AZ1sOkCVyBWZx3YAyft0le9GqDjw
/VA9BSsL9q49AjwNCuIPBvmVDEIY9h0iOJdSNn1aGBeDSsDh6iTGUMajnD39b0X8PxClCmZd/PfP
io4kErvAolsRaUHs1g0Rdnh0R80HLsdvoJ1kD+WpykjEQV5t4ao7SU99bMl5gcHlz170x1h7Dtr/
rEjX61BZOIvyWPoVRC0B9usCnJIMB+zXYj6bbO6/yJLPwzD2MnvBgOB8/rYaFfyRai+a4KfWATX2
Hs9idzwFQzgBZo23zjWmGFUJf+lQAHVhBMs/DhUv4E1Pi6RkZAiaVv2mr8x75xchN5PSqRf2biOA
fblu8vqO/uy9g4LISGnEWoCAI+VqQVxtnsHGSoexmq7xU3JGdvddwWLhFLClmqsWc2FFZTiUHRua
9u0ly31BXt6LxjjlYX7tNnxhsy4G4KgUpv+2kMuxxFxSF0xMeqoXZkp6PebOxqGf5cbo36dRID8q
szMees9TiJRP6LUT4Hvf3LT22AI+1eWVGiNxf80uKoVQBMaEg15IB01ag4naSQ+5cgKmL/Wx4QGE
Xtl+vj9g57gLYNeD3W6FEibLqvyTMMTfk7NbSDdqe3gTkDh7+BtZowHILv/38J5vlQ2ExE5eMTTk
EL8paCc81ddmusK/f193lM/XFXJVxfaJ01D/U49uvKTbV6BVA98vG4uCdML58aQRoCFkeaCM/Nbg
zPAMZ29l0mrtBF7BcP766M2QYGmTHRTzfXynenEDr0IJUBqnh4QmGOqM0wpZLw7dHnysxHb1Cp+s
aMz/34tlV+r91sTIAJkHeQNjiAbyiQ0Zsw4hbMc67ecIgbYQ4Hq75gFHDjKs2MwKK+0DIa2zvuwi
vD4Hc7yawTyBAXs8ugAawnEr53RVwEwi9BISzXVlp12AWEMC3CJhRbYAY7j3hB4YITKjTNra6mnX
l0OgD/VF6Z7PqB1xyPLc8zNlnuSJFeCmRBjqq/wsK3DWQaLzJ4myb0KPll5z5N2Gi81zUFtG4cxo
sbi+sASQmmd4GMnZuOhxCM2V1yCDo9OJepsZ6ZuBeQvjxyqF0+Rz4FukyVD1WWkBNXZe8GBXoKZv
EVSJmMafLtrdYWxy0jWZTaDsaj5ml9X4Ji50pRxKpWhtudb8Btr2ngSS0C7Q7TJUNzF5igrT4IKm
xSH02FYbOcbHET0aH/O0oQLpHWnXN48rY+mRKPlMePZzqme6pmQrL7nMLbw/pduc1MYH5bbA12+Y
+dxDuogh2gPL924FPn7qpFT0Iz32u0u6M9L8ZwSa68PPk24rGpAAwvqFxGPL3f49Q3l3GCDs9LrI
N4QYjHUpE+ROwGfe/Pb9XuWcqBRXDvIpwqie0vmpZnRxsQWOT+E0rje6iwLngE+jnQbxP4CfhU+F
UipZwOCKiu1HlABVAVzWXteEdMO2AOh73T2D6vbq4JgYgqLFMsB/O2gZKfNeAy0VdSkIrS8sVspQ
Q4ZMM7buS2BDwCHsAOfUKOBNlLKq17ZOJnTK66pn/ZyJq23UqExXIzwnPz1x1gYAMGfxvxX6ntqG
y6Ai4Z5zMvSIARYg3YaauPaDsX5Dn088C6fdBop3hNmZC7PBLc0O9x9ZYP6aLRVVW8PZXfW7g7u4
YVXbvbcCDcXrPCtIsbVfODi6V6QhIr2H1vqYe7VA71RTemTz+1GI5GzOU3wz7BAoYMMWSzr2Ibtc
Knt76sAyeCKjiw5nfjTQ/jNlt76GUPLA3PLi6zTw/fOjgpJr0aIqWYArGncCcbEtdzL1qs6D6d1z
262hSODhnwXZkogcAZh/C6oTkRAolmsrxIHsy+YP07K+ejk5G2kG1Mdk8NW/WKA//DpwgE9kV0YY
EZJryCIj3YzWmOEffC659AYj5aE1FLzaKCHIU2WGdlMS0RcUi/X9eo25SmsMWIUAcAc575opPxbu
QNljVoleVlzFFKCKDYO7+MyF8DidNiUhcnQkfL9+0oLPEFPEcMDuVa3j5I7euavj2l1schT/lKgs
mkPfsD9ovfx+L5VPnlBID91411xg7/gmKDUGRikA16kuiECotP8G0sZjb1rzCMXugH9U2AOCrB9o
ZPZsVTHX1YmjpKt5OxCXFenY9Iefo3fwhmq98Rb+hted3ZTXjXnENa6frXFc4ClaZnQjH3VBUUHI
l0GMuNbzXffrYkcC6SIDUQlnt27wpWJs3vQNbSi+zjBJrkiFnYItHSbyHCYDw+BWLM4WTrqa7Wl1
yq08WtgQ95JvQkvEfD00D04rONJmSnPbk2XguO27k8LH3DY3GFWCNHzak8QlBnOdjg+nIfVQE4P5
V18d+tchWxmIJzZbKKCTe5gwpPHSgNHEA/D5x14PTHWxTDm3WmrEgnjMZjvddVUtOiK4gvCl5bgL
utCeWJZ445NrdDBjbanUnHMXo+eRU2nyioBEZPCcwPCb3cvIXpAlz5GwQGfMpzzD66T+QLOd7LBt
u7xJuEhnt2OVIyWpb4QCNR3redehj6fMTvheWlBGtdUMExJTlHY8EOmTl5U1IB6j7MavFw+QCS4U
zO7pw8kO74pQHVGTPwEEoUqRdJIj9LUx2Xb6cVL58dlpSRjXANLX4C8JTPdaoG9Rs00sVU9L2rOl
LXaHjULTtViXolB5hXWLHSPASjyfDljrh+h9hbMy92EhBHoAtrg3Npj+PtdVf5nkN8oic+y1/TkE
iE5lKRweQVPvA4NkAxW/00WieihxoxdjWbXwNfSeDAcNz3WtUL2lN7m8AG5F2NXoJGBGeRb/90Ut
EpOaYLPQbxZ4GyKjP8X5n4kle6oIkCn9QmgmNl68Wwmo1urf7If1a0hBABWFBonxhlPJYEpVssfK
WzlPcIuzadGNvaO4iERkbnFBoJHAxw63mUX0g0nQTsbboHcjnkaHmBjL5nzmKebbSOGO9Sdehxs5
hrFGNjfM5Nqyf2kpUKU8M7/R1N/KHkSn+wGOu/KRGdPy0wqVKXMdy8/ilsWNr7cSLC4SZ003joN8
Cz0LnhRqjHLhSMOfUZyadERKIonB0v4Rq4JPqgZmUeU/hwh/xpjAShSY2I9NjaVuWmF8+2wLBcxV
1tiwo8gcCkQTAEyeA+8jIXpQhPeK2wmnWtecIH3pafEnYu6zam/KNudnkX6k1lsfm68EbcxJelUV
krc8fh87mteQi5PQYU6n81HzKudrQEMgt01rAbCCAeRsuTjG1WaHZmTI9p7+C4lFwJYJmk3IFH5W
YlHYGpwMB4DVZdMBcdLJe4nlbYbbmHkl5jhzAYSF4X4/oD8l9q24GA5OhIo+vbQFsS+p4kPegUBQ
AYazn5zEEXjqN7LEOJNWhLbGFSB+AvGw4pf8d0CLRqxf2tghbqUtTvpWyQBaSdk8lKrcosvXCcCS
cO0nYuLCIWHjVRAojquvC62tWcgeBtjB8s2BXW3X/oTUI1tJ6BFiumFIbtC7bmh6L4KfiBaeR5mb
LmLBSNKJ45GZg1YM5sJdneCASMawQBgYQUD+Jqs3HDTqMZfIAInTbdiBbSWakMX1j1nvjfXWADc1
lvqGP1gmI64KSjBNsoJRaSarOqqEtllQDcP2jnPwXdDdy3WaSlR7umwme5iHKis5c44c/WIAo7cM
hqPNK3LsS95Yibjpq52Q68unRBGU8gnoTGjdm6Fnxi1eJVM/a80bCoBZYx3IPVnrFzl7hBIo+9Kg
sQI6dQ1f8dn3ih+chYcZwjbHoX8exAr+IoG6OyAHdCL74yFzaiC7Gfwp+uGjMg3Mm77EUxDg6t4g
gtJWoVBnS989nnssgotWFhI8YOtSl29N9aJmOwO3NK5aQnjr8n6ymomwk7OTsMCitHW2SwTjDphV
mSUSUw/KSJ0Lyhd134m+0xGXoYO+6OF3xmnQ/LBSUfbxd2g04b7qhEGNhZUNn0TJ3G/Ri1JAbIJI
erVp1ozSyt5yv9LSpl205vo+punXGcXDKrBz0jA8LFL4p2Fa+5PfPvrvH2eeC1vEkXEEoJciIBti
iXWEe5e8/gD1wBycddtdJItCpRtTyVH36B4EDWQBGASOc0eN2QRuYsmRXccsNzo+8A0Tj9d/JkHa
0M4nfGkxiAZaKYlyi10oNKil330Vh7E7uSoPP+cv1TSzWL1D2HlbXREdnvz6Xw+eYHk1gXH9BZyi
fqR8wJcMyRECnWkMyFKhQJk3mVjdN4tHhPH0nRc/nt4R6El77RAcZ6jUaX9m07hvOiGGj7loUzFr
4w4RwQZ6gmIWY3dYHQ4CZBalgcqDymX2iRdE5Yzch2pkCwseBgOoSpnktnku25rjMhYcj7sLk225
MFFy3QB9H2vk8Fqa+QMjgnKYSqTPs+YB8yDizwL3+VJ8TO9pTPKiY/Zo4m39n1wFeBnZS14bhdYy
fkdTheN6hUAsojd9IMadyW5phXjMJkk+v4dLNj93/hC8DgwtM+EB5ASLwIRsYCQ08Xjyxeo7Y9At
YoR1/PcjKm8ZA4YTQuVRVV17zNfZU/DfTRDUGcSaO0iWQuJoOlDKZYOMtjmnjVPEPYK7sUsthmrB
lQQTb8Tr0VH5G/vsBbUBmxBleVrL+rCXou50Qsce4HZXwZsOl9sMCy6UTPXvRl36UAMTcmtsgTTQ
sCD083A4YwIACMyjTaxy5ed8G73NatoXhMwhHkuPkVZClCYoeZTrOBMnaQdRZEVok9kpdhWRfdPv
wAxvNOMNGCj73pgcRV0DvW3vXZcmmJKi0epIcMrgydYcqzOx88YZcqjZQRXYu4QwM7BP5b02w9Cw
kULeTWyM30hZqsnaXcYPzL6zieZ/IsU4wVuByRMhnF4p6IXR3O7AKRasbtgbVlPlLKYtUImSJduW
tjQpxozp2HxGx25K1Az5xNFgEWSqIXHRSKDXXOGtwWzeL/qWgIpfybTdulYjNP6swYr12saY/Yhs
eHCAYWEtkre/j68sTNz/7KcMenCfp36LPS7kZyQENg5GeiwacYtq8Hq+hUw6018Tsb4YINdi3Cgo
Nrn2xRGOZQmI0+cLhxkxz6PkXgUpe146mViDImdK2TUQl4l6FANY1rY3h3muwNZgQTCPTuIheeFu
oxe1PoJplrM6uAR+DdciqW4LSX/OIUrK27TSuhjXr8Ee3MqfU0yXoycy7mjIitPJinOMooW/z/1V
vkleQoVbKDHFehe46x0DBo71RvJ4pIx5BH52AYYNKGj283NHQi6BrbLmQIFQjpY6x+6f00ksoax+
HZPZ/9NS/DNRHJTx/Nz8FF8C+MgdkDAYDZsIiPhhrZD1VfopkXvulTiRn2064xslxmClBeeVFqai
im0SZmCnhMWCwUeZTB+ckIywUSL8Zi3zShZG0+8eHoU1ZNOrgIp66bAL/sUqJpiHXZQijpb5Sw9i
eY2s4nGFPAsurbi2n9ZnL3MwJ4cpsldLcoXQw6+/a/7T4jRBMSv7GcJx5h4Rql0WVlZbfLVza7WZ
kbF6Qf12sqAKTtarmP4dg7wo8n9v58VaCuk4eoLiVnjVavH3GBeD5lxbFnXCgLoW1qGUmEYvllhv
K1EBylIyEm0nZNz6lIXvnsY84ZJA0Ogts0lY8zQ6hJ/zGchepBCf9sWBJNxjw6CiA4/gFsxMuTJA
Tl/Vhfkn0HOMS7xFPPG2Lbwethvm89E9IwM4t8y9ykXpfu9xWeUwwrz3/U4FLZbhPj8onwa18d/X
/rbFOIz2WWhdKtaCV4GYwTcyOla4u4KkndNZiiGUfU6+qFQaOeAANmtCjXZ2G1efMpgROvPn8v6P
k3brZeV1KGZKuCMh4zzXMmFM279kcEmttbDpgdkyP6DWiPctpDl3dWwLdFWakCZgGy/FUBuM4uYq
vHbEYVaWhNoyVOrnNp+1nHx93BetygQrSs6Ga9tvoG+rMBjaJmhW0b39Zxn18OSuI5SNykb4Yxbv
xlSVOt917dbU7jpU2QYs2CWCU9sR6weId36+Xhy26UmUcC9EDhnpofmAV3cFAW4fVtuxjliMoTcQ
VBmAzWaCpVDKA+v0F5RiVxiSYKPixDZVoxqrnrOVAow7vE8SbkRwkgl9yAs4XSB8zPPDkcaKqZK1
JeAXE++Ag8zDnTM5YZhZDHyeQTdViMeOX+4bVw7Upb267D2kI0Mj2/tcqTS0F6XFTVs+hXKYc4Xc
x3oRcNVtiyvJFPcgQzxdITLo1H1KBf9vMHQutBzdfLqWJBd7l4YBOAhktFexojuU+EZPqAwmfsMH
1WSt+t6iJOiMb9bpncVmFigG4duJoGpFEqNRClBePnkUb154H7iGETGalbb1T7axE7PuuwHmwpqS
7OSReNul34VzbCDDoz1oeYSvDyLUgN+KI3DLSKZNZKFhAiVigRplNMw0tex3uDe6Is8pgWqps/Uv
z7bOhgJH5O/FYgikKyijxecrqAAU1Rpo7z1MjQWQyPnds6UezLluHMgtg0oJivluGgyYQPQKbzuV
vGag4GQNNNpYq/lZ6uaA1faehySAOVzl/gJ01WIfRwDsycD7u1bVOUj780dTgL010x2Mbjs7Xt5g
3T2DTbTre5A49Zop/D92hE7hrZngtkHGxkoltm1UgS1VxnFEa42AxB3ugzw4QNn/QAPfOKAa1RSH
4njoizE4kYP6Ka+rzSceS00qL8QW5L1yvfyOnCNmKDCmPFlo2HxA+kTS2ZdII5irN2NVA8W1KWUz
P5oVcsPYBRyRUG4522be8HsK7OckRhuA3ZXaT5DAOjY7PIh7kksswSyG6ekMptcmU8jUBocFHjpm
1VV0e7W8vVqi7GQaJrQqg8JvcwearYLqTKfDH/HWfsU1x/nPdHPyaWs2xv1au1/ditJL4Rsd0IUA
QyaCpy5YYOO0CNdnxcLm3+zW2moC/mSWV7GEohOVLXWOs3dyeYM7mQT0pBpxhx5zR7RfowmGl9DG
Fj2eBO5F85ecApBNoD1xYNcq6dTylM+x5GcsYv/uor2EwJD39p/BSQrhEjVgAdR+kwO3LDKC0zAV
2v1fq0ZuqET6JvMYN+k3eYYH/GPuJolGOjmEYvENOK8CthhXgr7AdHEKoUbAudDNhW9addJPjeFO
fI/3bule2Oy0TNyd5qfY9asQScXk4k80BGYmh/AlltS8GE8QkO/EvvymFYv4P0dLdw0Wcl55+zx5
oIcDkSFVvqS2QYAaJ4OpqMvLNbljIQ8AfNzTj01VMXtgBwcVXI6PR2j6dG2IUpCz/uOcrQo6ojKj
82HbDTJUfliFc/yKzwXweVsHqA1DMuHKumDIAJRCTvvTx0CKW5EzWGEySy1hOTUF5rYCWJFk9xLF
e397/L9ua5qR7HkOLlz7djPSHZjiy9hE7JaYVreDfHRpUWg4w9oa25xsC4dVk/JanZ1CeM+w+q9f
1HstR6jH9/E3arPLBRXMsZmA5y/5Gi9PYlZs2zgITR0aU6tc6QUzpoaMLzdqvUaPs3bhJygSTZrA
jzlIojGna83zyJbz3qc1Nj2n4cYluUpyB5DFOfgLZ94mMNnHQgYbR1wPDbkY9vEh3755md6W54VC
qCkEOGkIkcJofe+D3ljknzCFuHwqxbkXJD3HEfjTrm/1J9AuIDWDrOVaxfDmRF5Kz4YfzntKfSL/
3LfDDiHuEnxVApPgKmSG73V9NA3X/nSp6JHNyko2mubiEmrK6m8brUH5QxU1Kpbbt8i5LCkIUlG9
RJK/ppUnX2yY9p74u/zWkNq2jKqiSGzUxJkpKLqpLjpqJrLd3iRtpDNXEbBRdshWzmmvRIOnPvQb
cxkJlzsmoStJvj+jb96dj3BjUti9SuEhE4civatH7Viahj8RqYMS/7TefBRTkynBZUKJahHbUXC7
Vq/qKNV8BJC1Yyd0TT4hR8ZmV0k0blOwNu6cm3PradtuBQ2Pw9Hr8Ya+g0UYjh8F/CkR3QgIfMuE
PrEE/rzsIipc8D313616L5q23lcPuOY110tHrVsMtq4JOx8GUuZF/wMy/6e0j4Xscvr4ddoDF2nI
KR+w99pcU0FZ12LB0t+BoRiN4XmJsiI//3o1oOQFK07IcKnWLsaIJeZX1kf1TqMiZ3ooWgl79vwl
x7/M80x0OAPLaXxM+u+YTsw2mFxC9ep/Q5+zSHUNeBNGIqzLBsMXmDZvUpaHR3D8nadWWrkVxfOi
mCIUQhjtSFgvw6aZ2VPyw+u1YpUVCNgiSuVrZR9myqxxQ7wtlZEuwpsPw6AzluV2UiJAPNXXaM/7
XYIkoufOho3oRMydbMQGdhFQhGw2nXaVf79QOnmBXPVpsg5C5KoG/2cZCOdDnZNDYx8NAL5IEW7t
tMH+vvPMZqU/YM4aOOEb3+QO/tQ+Pow8eCmc6nIEpC6FeDrx3hR/h/5DqF1aZAMJR9TEQmqhEPGR
Y8mvXqN/buwn/3AaB3W41e24FNhcHPpHz4emwu/xycT0IgwjyXD6i8ha2QNFbBWQpFStegpFXAPS
BddSoFoddr1NAtoJUZA3Xg9QNnGKTgvvJs6/887pMLAvnWqvxyNFLfsMlD8REBzXVw6+OcCLfCt3
YzGoAxd5WjQubHo40YrlKQJheTDfEIsfk591jrsV1rlU83KhhRfGE5W9fS2qERbUnUVa/E5jJcHh
CdCaIHZDI+JJDY6wKYN7G8ILOSp+yikHWQ2RmQmPjTgjOtbome65SRMo8kRyuTc7it0a9gUqjl9+
nzfvqoPpJDl322enuA7/ezRgtVTX7KsKcPBr8h5wHtvoMBJFhNOATwaQ6791YNuN/iSRLUaV2UIX
FF414dqipxBwudDvo8vWDUZbIhEBdExlD8fxI2M2PGs0Qwfadd4zaIMXWtgPqMmAHcWtjJrDAdyv
9Rk9SOP960Znacj+NKxjGbW4HtIxKh7Hc6hz9DwZ+SkbU+2NLQ45qHfLD3rx9fr4EBhXOMU0Rmfh
4Zmh5psvl4Va4SE7/0jjF0LxcfWOvgS7MyutKjehCRfBFSv9TVoGGtSFgttANMrj7kxkRT3GEQ0T
o1rxUsnmICz/I/GpAty4KUzvnfGnnyXSntWQ+GDDRYQu+MkhJtctKByzmFKFcgaAHm4K/hCRnPEV
kD5iD0yM1qZKPk4W0O2TRpAhbGQSSwirhy6BEbeVyXWpQ/lyvfigePQ3hp2pigfUxBSVJiIxheag
oh9IoBS1yHWKoIVYLSDDdjQTkcOEyT8seWvo5oNAUHj7EmAkpyRVVBrNPqPcWKIviKHRCPccSlk7
1b9H/AcBXLLEl4cnV0bWZGcT4aVHtvqQU3JyDeRqenYSjhkCkdICxceiqwJfpg1xaVHAOn8Lr+Fv
jWEnU5j9ujHAncLBA63rWtC5nmsXLawsZU7dCCbQ9MejtCsTbuM2F5XkjJ8fncJ6glrA6Q3xLkZD
dkztVsdmxygfaXjTroaJhlOqt2BC+wuslyF0XgmO0Cny9DgXpRCbyPbQJETDy+6TbNGxgtdvJPlx
zm2kKStDWpuzdf6jj4BnPjvpCgozO1hlRY98YfSTGk9rnMRvbBhIYdzvTbKTHwsQkn+iXAceedCl
gGjX8LiopclH8UUkKVPDtuCnHlaacQSF9hFnVF9/zVJjIY/6oVo8C2Ny/n3dLNj7qlhEOTJpC8EZ
HkbttRgMgZDDIZfv1oLE1g4Q5sus/NkyPC5CksVGXBTU/scE43diD8F+75gZ8ZhLirxb2wi6/KEA
0pr679b/ye20U9GwAi6hGovZLsNVPPAdFAKy8xSlKE1lTrcECt7wIZOpKqAsEduiKxivrb5UKGhc
fa5M26J7NpFluPkJk6BA3lilg/b160gOYZISChMtwSX1djSXnRnvF4okgm/6XWFxpRpMJOPoGos8
xdQCCNodv2WQ6Jr5Qk4XkKLYC9S8ipcrj6bIa7OLttbylnYibjV3YPknxwg0HVNPUFKS8FqOWt+S
+prEMTw+VLl3JQf+AYu5Ura3UiCwpVpu5V+5isAdH5wjvKP5mQ77Qq31tlujMgQjUghMLiQOeOhc
z1XYXU/0oh/dAwHkObhhAku9eMnJ7M6ieEEogamgqTqI3hPLhDhV0+DDP2TJNd216ufreFYX1/09
kkpwe/lAfCVl19Q0o1wuq8h7Y70RrK5PukB/aOJIsAFMz2QmVgdUUYC1Hu3J6sF/PJljrCq6ulYP
YrzJuNm++lctVX/rJFBq1GEqYwAUES6ddgl0ys8DV7CRtKPnzXe70KcAEXzF7G9Mal9kh2KJrdSi
6BcifRtGbxDxNcyO8ZQ4J6jb1FAw5OAmtKLcnkbKBqVgIRfPyPsmZheZgUVtTxH4HDeg1+EnSUhB
xEXEQ0521mX9vjNfYUoQWQmZM9bnPLjkXuUh1aorEIEGzGjPibZ1vwH8la64ETbnC17/ToU1zUYv
QZ2oig5x2a5ZcixzUysix4w1n5hZsmzSHAbvr+EbBJgo8uNAsngu3DKD6RihL6M2EQopGYw6AEFR
jAHqxSPCBA2vs6nK73C431lkARSoBVrRFa76pX7YhSZG8NvyItwk7zAPHXAYF6BOZujVrksuJzQ4
T2eaAshH6vLQzGWhAADYTeRzS7f8+hhNivfF7EftSHdhG1Faz/10Sb7HbbNPmwMDDwIqwFLQAIvL
USR3KZ8jiZwqiryeEVc37D0pFAa/F6eRdaPr1rc3A0/bwtdKoKPxwlJMaoFO/KGRvm30g2M6ynNS
sZ5xKXuBLMo46dQNQPu3Ruz00sSlddeKSq11KYhSwrvmJ8zeyI1mCG9MVAPykn9LWPsFDlc3ErMw
18+kRvplqZfoO9442swBOxpJYpx+K/6emdQcIdxutve1XAmdN/8N9GIb6S6AI9Vng1o1mQCSZTk0
XQ68UAvumL6X/mN7DWZFHrG5QaSpfcOTpsZvmFEVepv8+oTy4P9uaCUdjsbU46fZxFeLAYTiaStr
59JVN/KM8ubZosdziSaj/lSNbS+AKH/snAFU1bL0hjUUsxuGG7G/OPZ7LxYCosHbww5jYJ1Tshv9
OvOUiccdFc45J1PIOusPnSc7p6vc/tOBnpmev8LLTXkg3DAafMBQrKCkRvYAisklt72QDaxe5Qmw
MdYQSeT52qMKEN0r0xqAx9R2CqqHyHb0+feEFewZDh79+HfL93A5l+TpDbue8uG53i67988vT7cA
6wVAQemC2qWY+hrCawOUD/sLmefMouUzlK4MpHKenSNlH2PH6bVbhOODZV+Z6gCJXKPuU3+3ZVSN
XSTAOuJAr2pkK9vWlFGz/ouCMxYORgQPzXc1r2XL2eUZXIt76OB6YbVVIto4JJzdPV0l/FI4m5rk
aAQ9eW7DKmBl0wruficNC0zxuMKr/0nclD2/wwlTOv06FCKjDI/wXkWY3FA5x0YsY+gCNzUsWIHJ
O8v5ki0x9a/RRwCWqWIltFwWVT2kKOqwY5envNoiv7QuGaw0znQK4b2CGYr481SIBTBIjEonZv8A
7fyep07I9FunNeo14WmxBc2dlSfUsJqe4OE3N1o+/UCu9XvS2RsHtl9xTyc+YYjoiIK0F98hWQaw
P+iBQ8djdFifxjldKqvNM5VoIr/mQFcwxTu1VMNAPjNFPtBz5Qlk72fWtcOHTiKRjayF/PLmqpDF
6aZzHOdXDz6rAhHBAy4uYanyv2UFblMTp0yIGshPV63iXsJWLUPNLyQZaKTKq0c8aQYscZ6cLVHU
lLB7ah+1Dx76Qqu9lxe8NxvYPjYxmXFFUcIGLmOWEhCfdeMuEN50tFcFsSGX5WS8DPuiWIuJup/+
4HnOnWUDzrjhI5zwDtGXtFZ0t/GQGXdD0r4krN7Jd2XL8wZWKWczl7PHguLolcdIP549wtoVTSZa
iHbiEIBhRiLgEqaJljcuoOHwnHEQhfNVg/bCeWUe/gjyEeekQ20JARO/tLaa75v3pdijrUwy86X3
sdfCT1Vw2Aawj5ILROXX8LyB/hMgg41MfFByqdwY3qeJSiFWLXpcBt0nnyivcTtNH8YGh82XlXJB
RR0ARPMpf7Y8mxVaH69wVkxDyOtrDqTG/Ss9gqryO2y1oTk2zBEA9FR9LzBWmksb4Cp+hINKtyDL
YzDDszUO6H8gtcxEHQnFbdsbJzla/D575PV12sAqfTKPHqiMZQuPiwBYlu9eatOJvryPX+ZmJscU
y6/TjfQWQEXOQxzbyQz49bg6Ttw3tydfawuYMsbujz9WBnL7mrGHbdlRmBJcvvEMc4URbfyDTZmR
TqIDTcH7rWW1lIZzzQC4QEIe/qpa0+ai9dtcxkISFi7O7/s/S2EJLZTvi05TCQQ1GJlUxVxYzFv3
gxau69ZAHWa/s6jkt8+FFeKf3mjNT1NN5J65EQhlW0yNoktbT5SbppDgWZ8K3O613llFjR2k2nUt
QozjJzUOl6DLNwPNBqMssBF6VSN7qKt9J89gUTV7gFWcY+rdA8X3Y3b953H0A0FgBRLaY3HFoJrW
VEKm+kbcFrQL5JIc6Ccg0pwFJOyfCDjScF5+s00Im8UlxXXS1/2AZIR6k2Li5Hv0Csrgty70ATry
LC7NGvavIdzwy9wYxaeXtAdSDAmITaV3gYFomH5TR8R2umFi/h18uGSgCdjWT08hiZv2Rq0MXxvu
4/DEvLv2bl/JzpGqsqjAtRtazkrYvFmsJinebbXdQa46vYhMK2mIbv0lx0ugaThHozUrYZHS7pyW
oYDA3FvamWFmZrlIOdVFxYywFLvBrbsVikVXrF1IZf6Gynh2aB+3lOWIhJtdDxmlo0lt8RM+/1t0
9L/xaCDLscLIt5RAgB8MbdIdFgv1RMZBBtuDio2xlJAeHIBNlpr8kHBCYWGOSIFwHeaMbxawN41+
OrbQ2DXn0JMLmk1Wgg/1rpu6rGfdhVZ3YAupeS14ZrKD2Oy034lwrGg+Weqc6Z2c9v4VsvSKkKn8
f6mz0OXqT1QtSKVK0I6knrwHbT6oyBYKsuJP4AB57OMrF7+lTpTm4Ci4RErNd1bYPoaQ/uKhTfj6
xIOFK5BgAiVMKdiy0VMhzFo+/YT75KjsGajkWo3MCNFgJetz6CJ5e3lA+be9PV9xLkxju2SUJoB0
Ajftz3ZnPCzoWoWt5odZEiAX5IUlWVgWUmIQnp+EJVjFV26O6d+TWVnnMAKnpPHE2V5+iz6ctWYB
RL1DFcUoM5yAXfLmUjFcQPF81Gp4x6f2ReXQ4LwXf4AJnXM7ddrhM0EcX46n+IkUQY0x6InzbvIo
URKtPqffFuuCRaA6LlSrAzxLNtu5rYrjxX/JpFjD1B1FO2yzOF/6z9NZBCZiHSTaa2KAXejvyX4g
5RX1IERvxPR+B3M01uuo1O3cWlPGbn6tYQfIkGpjxqP7dZLxDm65SrAHWOMYpxPuyapLouWKGxwU
bwmVR9+rckrVUQOnOX5BBItLmGbv0ox3aYkOgn/gNvNsWBb1dwJEmwbZj4P2jDtgq5CE+okniwwG
8EIVtY6U/Nb1xoouO6B3TMgy2l6ppMP+8r+1Kfeu2xG6p52qZuWYpCvTjl0JJ0hM6vp70fVgcG8I
ZGcHhY1OanVM90XYWBKcVu1TrJPD+BEbrhKHA3vTgsjV9PM22QVofcBIejvlzTs+l5R30O4RSsWb
5hiADBnUuBhfTIBCxVozkPra/ebhWHmxLO4IsRNF0EwxzNoDIU5iQYNZkViDB6l5s9b1vnR0l8Wz
1Xs2FjjBU1pyIigXL+bWUcOKesNA3d5NhrFFlqUxkYLz8khI7bLDa5jUkVTMTaH/GwXkMeULqmUO
Xg9fJxCD0tk+km4edpgtfCMqdBzLNVvo8T8vb8OUVghJB6JzbmyHZHUFPBaleFidFh2kj6iUJrU7
gBy/Wi6XlhPOER6GyDgT9/q1HScNcdyRjaFtnI2TFxdiQyCaT0OnK+i3p0Tx6i2QKF0LqVVs/2/y
9raTPgdxEmY8Ky+cu1HVD/VCgD1ZdNpUCALULvEHJpHeEj+1RAIgoaSNltN6kj8KEggxe+aUtQWx
G1LYu/lgaqUlJChcHLxnvmzDgYgmzMWZ6URsWFdszKZQykM0M3R7pv2kP3+jpvOx27TeK9991siu
y+Bdqw8/uHlVpKKle9OUh5xTWRQ7jyS9cJuyKyogSVMyqsf9C6UgMq/yr3H7LRG+apdeCMwvaPHP
e4bGajW/YRwoPYo6rVAb2RGU2nyw3b99+1kgeswG2JJxuiIYdUAVlDVM1JxvTAPfojsWA/062ChA
FwT32esJeQhUXHv+LvW6mBezZ+dleOR2GJaLn8J5jbEQ8n8wuQugQtNEuYzlRJs9B7vLDgNHSodm
PjGxTUh+iBdAxIaFtOr5RbVyHaLMm+mee1BjhyX+5JMo76oW/jR/gXu/P3ihT0GHG0aYqrRkQZef
rgTRuUUsgT1zju6viA4JvnAgcenmn06Tc5Hk41mCxGmquFtw0AEEbRq9gYeRuj0wOrMFVcO5BWZl
Oo4ad3C6NukedpR+KeTXN79Hdxu7oJl9YkJjnE1TLayxhKqNIX0FWdadK4HCHTVWfGiIJM5WvhJ3
i3Rojx2Zl9GTD8R9AUoDU8n1OybeAT/71CT1LzCQPzBriKe/MI5hVI6DydvMFOcppomUxU4cvBkT
uJFww4la0T+SHY8HLDpo+KAXGA0Lxc+XfB4fDB9N/804CT8xa4xgMLAwQzK1GKcTNQBLUaI4HKL+
fqqwOUIwluCTK6kmIkaXzGq5Ah/aaYBtPoxhNPCsYG2G+dW0Dq04dt1FVb5ybOVtv4Rak0OdrWiB
7nrBDgafEtZl+9m2tO6gsyyiKqEA1PcoQnmbOIMAVdk+IY0QFhpChPsJTrFrpBIG9rK2c1LitJDq
lPgApI3n4nTDSP0AJU/lndVQr9BIshM3BrcP9QFW9/M7gf1PnBqbyQaBIOP5/GLE/A2HGMHMw7VR
eZ7F+NwSi5uu6TrQfCpgNL7hSGia4xQ6GQfYU0CKH/RvQFq7mIEQsJJBfQrVaAsthcwQrspGUgqF
DynP8wOiZLjud/ldnykhX3Cm+VCwR0dGs6BNiEfNgeWxQ4RhFAXMdeBhMuI7Mvd4mVPkBiHes7j+
WYNHHncIUv75GTfHUibbe2Z5GRILGkdYm8uLC/11c60UwmNpggLo8FfV4S067efT4NdW1izlK4em
qft5v7iwombUq9iOHvCoYIMU3ZVAbI1fLB7mglBmVeOPpa3EJ4iCoAwZnCOcBSnDzSqVXF+oLgiU
J1F1kPMHYprB5+poNxKxC3Bz7VFfu3NYgOkem7s0bDc1lkOBpgejz+ZPBA9a6UazHClzRNSRyRbt
GXUOd1McxSKb5rxqemslg3tMEsrVSAjmKQMv+zV86UaMxtGC4JwxGUTUgt+LtyfbPCnIJJhBdeLO
X5ocj2eFpA0dqTy2oazqyKYDM1mWoVw0D+g4v6cr3FIFjcYYlIKSR/d3FeNO33a/+339kaJ87Sgd
z/wpZgWrTDFje9ofdIOhSy/jYa9Zd1GpCZMGOG3ih3Z8jioW5kpBdGE81LrBswFGfe8IGuSnUW6B
pAw6CKNUUGnBn4LmhyYwR3eyj8jHl3ji/c0nph5wihJPyhjzkxl5XOyE9HrrLr0bfsLla3U9EFHY
IVdJ7zoVE1kxtEYWKb7kp/lJHIUfRMjymcVx6Pk1trT4056o0KIjfKtIwIGuWN+9Vr5lOviIGG8f
TqAHms99qoD4r3cldSQxINrBfvNtB1x1jBDXpKI2ZtMepN/n0t8kdzFcHw/fbOqjDPhYiXMhAC8l
J2zZVNJwm8Vzk/YxJAM3I9xziradfwt94tRrBdPl50MgniDl3bCV5RKsG0zJiQW/t+D3I6MT4OQJ
e49Zp9zYNlst2qkQJOvnUSHg5oAldqNI5VmyTdawYBk9If3a+ett36/4+gjzkXCtQnUZUt4V0Fvd
YTesYQPdUmopMB6lIOz6bG9hQ5QpwS41cE7qhH2ZehL5usopUKQ1OaR3tclxoDHU7ZVPLxiChnXU
nrABqUaMWlyRQhpLcQmmF3ayPOIotk3JCWXNR31/wJQb3BITDnVCe1lOjgi2MCky35SNeHaaOW6n
J8yCho6wqRICbL/nWoqK5uv8zphWD8P/Uj9bY1YZdDT1vqWG1tJGHP8DZpTlk79ZcxYqHmMSKlsq
iyCzx1EV/VQeMKT8F26nzDkcd0fd36F9HYc5pv/FU3BANcz7sOq+6czbaNn2vLz0sP0JLyICWLwY
GQUG3zwGVKvD53DdgEoeMIjDO02id0xipDRIdirvGCHHDfxmvrKDIv3owhbab23DZkr9k15el7HZ
yJXfGgwcpzajl9jXzH/S1+0QKlh1yiGHneZ67hMHgufzMbZirJ6YkBJDFlg30+XW3UiPvkdh20Hu
7uBxMPx5nsX+OfX/6UpaIW3+UIad9km63GluiPK8QhG/QC2ZMNbBZMIzbx6RZ2d+8lywihcTPwkP
Quwx0vIG0+E1ofJ+FSdchZuIFa0ZfLR8DibRsv6ikIZMW3Be1VZ3zk0jHmOKVGoloB1DYvrCzyku
ceEEDuEt7jfhqiUUfBPP835H3/iWFddk5Q4a6B+nK8ngsQH76j6A800E1lEwTbGipiS+nOMv0RuG
/X5CWCgnaxGYQVVPEP7AqEZbCuP7MrEH0uCG9z/7ODgKwe52Mdvfy2Fh2Y/jED2/GFJI/yNDRq3c
J03GBbM60ABJimmWCBSEozVWoKOkBMIPYHYPqeYF/GD5Uf+C8lbk0d+fsUw6j4E0achm7IUpacow
O25JYEkMV6cf8hAV+aJO/dFusrSBn6r7H6pvQ4SjLjX98dAftIbVBMHtH1pB0GtkSfSyLTgdBxh4
ygIKfRmQLXi0ntFrimXAO39o+WneYYpTQnNu0Y4PjUW6Mtcf9MHukc6Qkit+QM7MUmcTwVhRGE2j
jYO0D3fFX58YB4jHA0VjJeJ5XAd9mZAAUIt3S1PjkJU4spYExILUHGYlqTsgDUwhVJ8So2wuzG5P
M2ziEhqSFvm29qMiqFgM5XshdnQgrQv0TNkWsHEQdKqJF2OrPv6T9fjeZVImRuj1MAsEL4jsBM3I
6t87LZOQ14S8+1fjcP8eiuWDW3QB3EL7WDYf8zwt/IgadArMYTvdO97j31orYJHETs9xem+VzYV4
3aQedeSuepr1hf43dDHhBYcRKtK6DRkIZhPRpXCap/0+3xxetjGHWO/adS+vnMBTp7QXiVdWmcE+
yYtcgxnMsxiOQ45wlyXt0iyCLlspWc7gw3v2wdYxJa0rFhZ4XV1+IIFu+Mx4E5bkFh7b5qigY9y7
R1pnjS3HGlWiTsRIXIb3swT5Z+gh9PkzmqiV9SrgTXtkZusAk6GOJI4UFjOV3y9Jz4Mf4NPiwzBc
VLKLaNj/dtESe4/m1LvmiwK/tdkq5tZdUY8whbzXTx6yS1DPjYukn+IBxQq7n6+bI6KFMB6+ZmzR
BWvrGivZ2doMCdkdz1v+sdBwedn/dLjh3rkWHdPcd0Z6nJk35qDc1J9REl31rpl3T2QY6Ukn6qgp
3BGufEOXK/PYgPL9XwlsfgFVgS8nXiNltwIAPjvxbz2Cb8N18hjKukFzGP3Ht6pCnPtG2Hshkwco
sveZQOeMV0UTi7hUC8cGWer/eSje5Sjm7qgKm5doknXSFJuKNDVcYnSr3QOmurCFH/StYOtrtp83
8bDC/niqZ675FY0NDFihAWjfTOB+BZgga86ucXRtZcY0wCrATYgipK63/SPvdcn90Ivkowobk+CC
DTFOsyJqXjaUIWg/yHakMN/ETl97pTC96kyqoKz6z2Ch4BCi1OQRJiyce29cGpgjhYP/dwy+zpnC
F7xRfuR2/eG4tF+j66fI1P8vnkr2RCHl225oks5Z+aGb6NzpL87cNC15db62TzSOQNn8b/2qdf4X
0e5Kkrkt0nFM2JfM/w8yMdPSAmLH1zRApSG+XrSLt6ctaI0GGoacs8NHjt6kvJTTXzFVPywzMNDK
dR0y4UHxyd/N45P6ydfDRJ/i3FkdU9ACdQPGEHVxK2KreLGqptXAr+msXnJCtO+RDZAd/5wL2WvP
79lM8F95W+OBC9920MPHRv2H0mqhdElHXOhAt+Quppfl8ppqVsWZiAfsHk0fmROx1g+Ste3sMbI9
hJr2QnHdRxf9PACsCltl8Z8u+y4/94ENEh45pbpkvIUhc/40Zd1d9ZgNvoRRXyAuqFjF+rgaqduZ
EILw/0BV4vGjoA1zV6Bv47gAE4MrOzfUR4GiAdBEoELctG8yTQVlUb6GMFDNNoVVJiGJwkmwmAnk
eI8QKbVo3d7k60Wb5/D2KmiWNM0N2XJjZwHNzgoEhrl+7cUimZPXfa3C2/ZzRwQLYlUm7ayaSHGF
koVn0laQA4cmotwRrlp0Nsh1pWtnFXGvQ9HS6WLs/b3TemmoJyP6UZTSPN+82pbBP06GDZkd7xlT
hcus+tAvMWJtRkpO6//l+XiOWr+FVk/eqhnGpo6wjisKhWegvFAKbdA5kUtt0R/02LUyk4Ky5rjK
p2Y8jEA6i7shD7qugNj7BkfnyILkuP1hMxFSYpd0ti8f/tc8lbWbcSPRkoPF63c5f1OfylwnNaP9
UMtnAPdtIqVckjSXG3QsXYick09BKAPdg++j+6zxDqENQVzDg17unfCZepEWw1st+ExJx8hsuu++
IqW9pVtHVe5JErFBx/OHuRXhhcoSuORmQN/dZnOah36VoXC3C88ZEQlsRYMiZ4YBHpbsFj4jLqWd
5gfMrLSpih1VIREo/Yze8a13HCWY6MIVqgXa35KoxVUKyG7kJLQkWxaVXI5vJvak8PZH8AXsVQ05
jh4xzle1TJl25h165sHGEcgDynnj8+OPMAs1hhCwoYmQSH8OkB86XmWTTia89OAMf0NTPqBwvnXD
GluCMLnsBRFHem8tjQ3PjXpE0KGIZXA+MImUAwpSIYVRO3obj02DPN9+tZrVBXmMuA4ZxsfEWihl
uKk7ohzzN3odN8IRTcKcDveW53rxxPDpd/ZK02uDchqJC2uxeZzk9k7BHGVWdiU/zn/LB0s82ArG
CZoWQva4RMFTJjerhRINyWhu3OCDqrhPldlxmzmbbxeglGL5Wj12fdkLzdubUPfUqM2o8sUM7KKE
3W3xB+ulyzH32IZ0GZn2p05C1uhS9OEbFZAbsQX7q/pE0aMLqtHVno0Tp9+ly/vMCQHjOQ92qTiW
zbgvWDTsmO2nUuYoMHeXryBgXgvJd6UFnCFWw+wuKNvS7FGn5qlZO7mxD8nHKaIFmuU7PZR+KPCL
arrKaxBd5zRSWbohnLylwfRGX1+U9qZ2qOHwGgpghrPPpUm4tDdVilw7+bT9lVKqFyifGChXe5us
RNZw9wRFCJSjHN34yZdBErxBcK91LtGaR1/7FOsTd6xeyRux0T07NSxpL2p5QDAAwl8VTBtfzBQC
02nzeCgv2I4rh3AhXZePxFzSp/ELymz+P5nyPF4n3iA6Ge51xv5siQ8bMKaG7AJce9txdphqjOAO
AxxQJNF0wP9VStIhQfXADOjI3PL8fgR+uErc2a0xrzaLP6z9fvSDs1OJbaA1xvabtysWCkMuYcTL
ecqOQNrWs3lQoLiwFbpZg5DqWP5Gk4z7e98oMSiF4LzIAMe4nG7rGrPnh5bnZFYT4LACv4XQgTYE
AcCmqGe6kRS6QFi9Tn2Rqt8cpIooP7gNp2KZL+zBXjnhnlTho75O0clhLHVBUNR2jVdMxCZKmgEe
QuhhPAMV9dAjxGx0OS6tiJIg49PMlSQK4u2iC2SGw0wsEmTYJ/0GmIvkNOodBF9iugbTXXG87CPG
hIIp3SCPT1XQsqxL7Pbtkp+UdBwzIwYY/pUfFlBrp+owlWHDybVkGSRzNFxwe3NCk9s8QEPbr8wo
nGfDjDP2G1mTU9nn5z71q/H/mtmCbdDXvUnHJH8RmpOJDo3eaYKf+iBqieNCbz8chLvimmfdOp+r
Dz53dJ25e7ZTOC8e/29K7FTHwXcBjWAV3GxMiuVC2zeQmA8sh1Bel+YcFkuOjS+IrvASvweuRQk7
2Wu4M8XjOlB4gtTpzEkjzv2DNRIWkePqFNYd9Di4O6ybNjs44THgAWbpaD46WnNxItV7482HL9X+
3bTpwvR4XcOA+52Qw91iaa/RhiUdjnGbj6OoxkUh88KRr5BZcoJbdaNhOZccHOsmoHtG4GPm0ZhE
eGzQmp7Ny3S4rZxAepW/5p/Dkb8sjdQJuKvS5YsgZUMiAVQXBww+aIULD/0h/KWLGqj5wi3b67+5
a9b75fOJXEnHU6cowtdzwHWPDF1eyBAgXzxq77bPDPWDVhC0quKRYYPP2HMyKouR1aNQiqsleRoZ
FviGZiyP+ieVXkCIQ5UAJl8y3PWOlCQ5F5zAfYKvAO+f9XKoGBDE7xhlK/MvqVFRoBdIqBop7Pg9
qZ41Kz1KGHE1bsAhpP8yKHpq8qt3svyVRWWIgHoO0thKeDoPPgNhLNyFlNFXYSsHhdJ9G5PUysur
5H68yT0Ydwq3aBX585/0JWiT5Lqd9vzu5/s4m5WYIhzJuTnQmCydWD+CMDghls+BvN7Re5tW09mg
mkFcdfKpgw8B474Ltr4lyulKahL9wGkdINbMlv9Ib/WD90+IapJjY8gS3aFoKYDM/wBnCUpLCTnW
IK8BcGIHTYQq0Pcc5cjaUWPgjbk83sCo3fFkp74xwaCQ7s0yRajeqc0/HN0BvqsGbj4ddcZ4yFyu
27MYJnlJKkC389oscOq4PTXNtvUMqcQR+rjxuoN5+QwDwQdMgTtXTEBCsu7x9bs7/A3N3YzMsqYO
MxXtebbxro51uJl/p0GPx/qAWr3lXffSfgqkjaKvVxFqWnTeKNVkI0IjZpRxh9V6BXvIvH/rYdIe
Byr25plbESjk7ACZB0Z5NKMw/6mzkMYoT1XXpxpuQYeBfaD4yXL6VqFzNAg1gP2OmZUmfF05Djc2
sV3vrcI2XV0uWlPJK0+iQWf+IA/xRzfL4mtQ1qMgExkDh95Ax2vU4GORX5WBi26Opj7F+NeAXvGk
TsQqZ0eKahF5Ic2k2eD3Tjjsno9jfD7ZZineYFRp2/LCzsoMcWWG6p1i5z6Lk3ytE+7O0uRPApEb
IHKQIIw4gMRKrP2V//R+0Jw/MWLL5PKzSC1RHMUk+3j12oPX7bSbAp0AEkDZ/8aYHmWo8gh1W/XX
pQ2Ml9t+5a/PlSda561uR2zAMX1upGR83LgUqSSwQb60GzlR559M6DZe2hp50lEvgnZ1ZnIvh5n3
B+QQDUr9MYB/+B31UFNt5nwgIea6b5XZbi1YS7W/7iPV3NrTs8hjWvrU4dPoAjFVaJHNdlUDDDof
QYikQmAURPLOAjvDzLZ/GNlSakbJwuMkY+N6oV88ZWK4+qNIgQq53SugmUB9/ags4L/Dud2JAxEj
iDcqB0Ayec+F5iKWnPq6SZuJEtTZcLbX3ER9H9AqQjpKrh0MFOaz2HAFba2A8nYOXnczviSKAb0k
+dZTH2rSlz1Xwp0vsGdyBm4l7HAtrn2QNUFmyxV//JMCABAfNpwF+oH9EVHzTh/swx0eQiMdoSPP
NwqQ3YX07+ZIzammkBX5gIyBnwKYGys4P0717lzIuUitR9/LPwW921lcPg74wST+p9wPmU9MZxEI
l4yEZfNKXIejx/LcCRS1Tiz2QHPTBluZJg8zttOLlCKnmQcm+2zFxOmOivZPA9tQN8RvcWh64o7J
7wK1+ZMmR4EgzOEP4EMGSPWkFFIbnjPDELSPTZrvTdQZpUiEejISmMLN+X7HlFw2RGQU45TqRMHf
MozFdg8rVBy+P3UcnL0R+MWX3q9nQzT9H3NUfcOaUmILMw5mYBI3jYzmXYkRHhO+IwuAw5nD/oHk
gNrtkCzVSzxU25vo+wkc7UxKFuFb7ONnRt3GeatV6eK9J37c9rehxJcJGbohGi/x2J5VSMsPdc/U
9vjRwPsmYBuOMChTUI5QlTVjBb1jBu2ORlXp1jTH3QCxAxjm5ebUiVmFL2UjkSN4uHrGQOdQn56T
14vNIL3zlOdsEbEds7vyjsK7YGCtlLLR0DgxG8YNn8nMbXv0f33wj+KFMOiRMLDimbB+60bvVn33
A5HgICLNCIc2ufUuJkKeZMVxSOBOiGeg5g7rpOdCkXRtAisJKhav/ACHtJKSEu4V4Ug/NXEvS+L/
Mp8JSgFV+l2JljaN0gv3HATi676ssQ5ey18qp3l1edB9YQEHYRWYtFwMQSPuS1DJNVpE8L3jOza0
WX90GpFpDxUG0ir5mQhRlc5vhSdRzhr2gEuFy/BXXCZRIqb+BGez5ba0mg/pmbviDSRudMJNlGfO
V5ShbK4GD4qZzO1cvTN9vpCnWAosEXIK+yUoaOJeN5aJftpsbIQey1CuFYcFR17Uux7X7puqfl2M
K+/nS7gbfpW8N5SqZMepoi6zY/bF7k4+mGxU7OPksM3n/LHt/177xOgqt/HmmWPAZTeznW24r1aj
3ZB0oy331n3FHjJQ4XqqfCvSIl1MHegb63vYLZ7fFvXa42cwq9avyM6oer5ek49IjLUgBe0mTWAh
WStTElj8Guhpj7X/RnR0T2zXdzpD7z6eD0G93bXEvKH3fESFjNyRNT/BEmrg22LXuB95jduwIP2u
OSTdVK8qNDoQzwoz9cxTl9pYGzJiMqF4p54CvkgtFYE8eEe4K4BDMeLh1UAH7B9Nb5bfM3HBfrsH
Xy9mQvSNh3FOBFJJJ3927xUB2QxHyUi8s/IRsR2rcD2RUMXYSBW0VJY6Kov8M6K7V0DvJRczyk9b
6ANp9ggX2IakXKH0KL9VQReOuQzSs6CpjU2I43Ym44xsyHqI2LCH707ydfjZSm+QSN7lGvylp1Om
OStHs01VUwbiXbuoGAA44i2zeZwcbmUhwJaG+nuppWBsZReNOg37OxQJq5nneGRbDJLFIo6ORdoD
KXehdiTxRTfLsHzu+I67z3IAPH2IwvW1d8xb8AcaIYOBobPHe+Gg1zUKmuHQIZJkmzrd7Di23Q9K
DKN8mS4Ujh8/4CD1DHeey3EEBX9TlGXDnEoSgr+aUAUIpQlpFUG9zatdGCjlFP7PjdFbYxTx0b03
yh5CYlE/iThJYRokVgyafgoDp091d3AYwK09/Z1CDezE11RQ1xCalY6FOtpjV0zvPr/Gx7Vb5959
LQKHxp/LpFFfBjet7I/bNcrXUOSRLpiG1K/2nUclDVcvDQBSGbBshnjOubmR/V56tgBHafxeYDKk
vsf9Gwsjch6z754uUN+HMFoQfammCCakIKp3VL3b+YeyinPRawcXtSdwFoMQW7qewct8wGgRbc++
D38fc+4Q6Pl+FuArhYTNx9aNIuD3h5xM+1xifzUA55R58aEIug9LUts+sBrItCXz0afwAbO+z+qW
vhVDp3eiuXJz96qn0DaupKD/SJe/zsbFKMDYlphACTNfyzvbN8n1xFuRGAYwdjCgoUnzXItQjdbB
HHBjiukf/+u2p1Gtwthcb2bZS/jSY776NLOb/bouPj+8zQzdoDrlRIqZRVNIGbsOVyclVGVdV5ez
2Enfb5TOIuEZCIB95R8KxRZJzbr5e9TyKxwiS9OA9RRJWR/0gTYayq8QYm5lEQwkPKoxEC4pz1/V
H3Zpy1S3Xf7kbHTSLISePQB79L7TssmXoKFQSfqdEPGMvPIn2KK6AmK94VYMhlr8IOUmQqeMxm9r
MjnXY6PRVIKwETDFP3Rs1rDmHBa4PrkSj6sW4WovkuRBinLKnJMrUwSCyly3nKPEefReuAyJeI/W
imEg1ItWdUH73BuNfjslZDFxEMp0tOwsn5IMqHxqZoBKzCBA6mJFt+Js/6PDZxmdXceA3aQQlNMX
EAv8lK8Cqluq6yd0EPGh+DBAMYIMs6uQRo+B6IfA5Qbi9jEhIL8nzqH2Lw68V86Enh02dSUKbVq9
7jQEN/MStOZVAUQ92jcc4jOikKGP+UKcJIJFM2d9+ljMEUa5RBizT2LReYNdkl476y+JQRUwH+Mm
IHAZ+NJbJyVcTst4BwbjmkcLJeJCLv4XM68F2m7z/M/SjlYrY8//L+7rXgYodtnWGHMYM4gCA5+8
pSaShJ3AZIplZaxbK/irld8fcMnmSUDi8tvfOH4N2BJ75oR6S7/fXKMRBAabCrjK4c0cAlC7SBPo
rsRF2YFAdrAdrtyUhJcpQnpoiCq7vK3ToudQCDWTMtdJx7pD8JwQkH1VSNux44zvTiq3WVdmYzHX
QzNotJLWjvRb4Dm5rSMDTTTJFQoj/Pc8+KUpkEPhkOQl3ydUNvzf3x3dJtvXuwbTaTWm4WVA9Iyn
LQOaTnbYQmIx34THsRzcyuXoy1wLcNihRvvEJpRBrTOwTHtSiZBWCD17Stz96xc5e9keF5aUDo6R
0IocJbeRkMQ0fkCY/PPBSjF90nAn4GdVF2Gq6MMuaRmmP0zbvYr4BdCiduhjsQjkmrbZ+WWbh6gl
lXQHFDAqfs8UGZ4W9xE6+D7anEHA4J37ICBHlmupYo9YnavtCDCyHHZgKhxqhjCQqGqpF2gJbUEC
3taQ1F47EBScm/iLXEEP98YdVqbORHeKZBzbx6cZI8sjkNxxkGIcBvL61oBEY3JSaq5r05TW4Zzm
H4T/36gBTBgSXgWfvXXbAmQ2isHOO2lRBzMfnBWHM5JtXw/dKlia2qIkTcA1mDGuiaUEclIfqbyg
ynbiFfm/O+FPuxn2pIqppYcWB5hHVLkCLdf3vpHGVoFj/EMMpulDF10XkCpdpAxuRlUZw2Z7fTuB
PJSAMYX9ChOEyQ6xGmM7md+IFFfRJ4/3UdD60UAR7LMzuPXScI9YjpSJBYZlXHufYj9dn8T2wMDr
BK9jLdOzJlHsgv9tOubf5ElKT+6cHYFzPGAI/CyftAkTlsaiSxIRG9TexPvxdFBDhtRM203gk7Vn
T48sPkYm999KlrP62+PVZ+9ppL8XbppXqIXoFh/YYtT0uVBerlp6J7xzw7sM+8ZBwr3owWdo8WMO
dNWvt/+6GZRNQsYBJ/y6jxLGKo262rMVfn7O1u9Y/hUym14fQTbw8rjcEQXd/9ZyvVXhv3T903aL
F541eV65X0hMR0MsF04EHi4EyvEBAyqNP5hdazakrsWPktP7O8itRYUpD9lxKyCwR2F4EoughmYf
+yBwWe5UzIGKZhgLKPVbwGef7EcEufwc90NhdXxEQq+MIOM6DH2YikdMfQdJwyHpJA/4NbMo/0Bt
ZwIi/FlqP+tqEyKHXD5n77+lXVIcTNW+0sjuputE2EbZE7PFE3lBOYgMNKVhybYQLIqS5qG825eI
vONRx3H2GsxAJwD8q84a0zka6hFAZnr+zOaFq1TDwihpaujA/IpavVqhHrmFXeCuaKLEjQK3NhoI
+geW9CnpfN2rNs0ewu0pJOu/oQEhTu6xlNN8beF3TYVMzBTeAAl8lgUNylwGQ+9+iDBLS2k8CE/x
bnLjGfihc3KqKIfpCEvajUWYIdT4MNC6uBoYBatkzRYwhj27yzscYn+CXjBK7D3izKVFR2R55IDx
J1rG3cz/MQJpiCGBnFNJk09ctGZDJFJpVE8z/bz3EhXaV5AdNahDhTwqNAsWtgyOkNT/XhLt6fYI
Vgal61gNvxYRVQxx0/BFbJVPvecpXTwxT6VB8k2czb7P0JlKqlGft2oQeaLGd7/4j9lapkKSjPPG
W1r4ztMOTztAg00DNfBTQ8ZKKAWQxpB3yzwpG1HJZyJifbfZvhni2J+RlCT3uCtP2p8fACQ3LGmI
kdvZrNmknoSdTjWLx9XifHy/QBcH6UJRddEygScgCn2pjYM+waYXonokzYciWTLUuEGEj3pUl3BV
KDc7XUTjjimb4wuu6aaM5Bnt0tnKUvg/0pyG2AIPA+YDiSPZ2BzF+66fZjbrj8wYlrnfAreNFbP1
t8sMMMicoDttFAJt+B38QxNTHU0GCMy7ZdzrDqOwfy0AoS70tj54/gdRav+Ma6sfMsDZUTwAZihN
a/ryztp7dwtkgUddenMu9WjH9Je3srvUfv2I541ZYebX1t/sN31hHrbgT6fMg8mmaVzJzokqT5ut
da4V1q+hf/83XD8et/A+xrunpqxoHETKVAMl7rzV5Uqienfx1RFe3GGjoufD+w3LfWPPaDG8/eNn
JX0mdzwqUHBZU9o0JtsX/ZvTkEGp6InlQFw+K+Zd+Zc2LVC64AGyrozCHhd4sdaamGeUbC9DXYAI
5PBTZ7af1PnsdwjVnRLmoSNrn87+x2Ag24uVmbeqOSH0SrCj4x5cXL6KatkRQttz7b5TcxSeX/Jb
bXI0FeD3IPjr8CB8f/VgYENba6nFtSNjeleucJryN2sEtegcLb8XIQiZyA1yc703ZSXbPCjhHpaW
87rSFwT0TV+mV+zODLkuVsAhasUo7QIRQ9xculnCCFyz9Q8tqJ2aLw5LPC5Jz0FNMGA/DMS4aMF5
1XjhRhe5JbMevaZk7PBPAbr5ZKjvpmUI4q2uoR4ISQq0ajq2QEHQqO1GojPyi4Tur54dZW3DX8yT
B9xmPdkgjCT50vLn0oRfx6z9fOr0lNpE/cXQSoMgtKCMubLwVKJ9NYgViHfrxEUAGYqux1LTB6zh
1pcxsEyXVNAs0jOUDL4s7jGOLX4K4EYz7ggRsgdgS/3x2bOBkKaUeGFIPblbuVeGRIsJKcASpfG6
Ju65ISUNzobxs/AapDghLIKhhHyzfzZzz1xbq0FSjTJR2MJmZjXVhnEMw3WEGrbqba57a5Dq7ym9
nBHPfjpSV/87MwnmpkEK4/YwmF+rRH4pGXxsftv3r0nVob0SzNfgB7bHrJIZsZJd/pS2capfPBR/
uNEcYvgNnZBcqNjDSOlo/P/AAVhphShpbQC3iy3l430CT6Jd1z8j8mRZAvqAkZ5q+FrUZptmgIDC
PI+7AS4CPfLsND7CKT4ASKWtSvjfYtVilFhfh6K9tmaOacBbPa182EzfJr3QsExJJbLs910wL0qk
2abGHuiZbHJlL/SMigbbW7RqwSKxScyhRRWnZlsyWDJpKFv8Y9q1v2tUSJGDgtu6AdQ+aWOH66Ow
muI5kHsli03ZNArM9xFXdA6bvyjDvQlMrMw/05EbzGT/OoQvvpo51GcOpArokGLx29ydmjk4cGjb
E8PoNCjF6xDv8RvQcNFPUNUU+5kP9bj1kfbHtbL0O122m1lPZYWDpUUwRmn4uUIK5t4MfZu+9gQH
u/7NJv8et1R28IxKnbA7/EvM0gt847oP8LiFvT41bOBR+70eA2N0W+Scx76o1ooxC6+H2QrzCYIv
9v2ngcJRk81z9I952VhwCvLZZjcQnIMpkJ7lm++C/txxlTPtD4gH+J/i/3pdJwlZ2QLpEzyPNybb
zYOQd/0b1ro33vot0XcxLQRWYEpe/tb765UZ/+9doZnZb8PO7nz5RnmNE6MLXRHErbHMEc7n0vLi
I3f8OE+gTdfnxhyWMYY/cltjy4m/IetDEy5AFZM2/TVF44ZyRES3luVwTvbhFATMn+i63+Er6dNn
10y6mKDgXEHnrSK6vJMOsIX/LB18FlpksB2fXTyk2wbFaLlxP7H9sT43NvUUOpINHXV1FkrHd4uQ
T0V2t8A912Hwy4oEpf20oRMGwbLcMhEHI2dHfegaNja+9dyv90cNopnoiruayOEMHOfuHUWpIjVM
CyJKaTOZOsDxQ3xTARA6vAWES5tVNYQuvugQpFmR+rfBFbhMW0xKfhVhYvxvxmHLZhzs7gjQHe8V
xexnenMAuj8bVne1WqfIAbquTR4zxeeGL+5rEjRIcnzZ0R8uD3Yyfca7VsN+FiEFvRme1dxIfbkf
Uk56b6O5hGEX0VECw8EvjCqNZ3iu+FdO7mpvoGMO0RBUgnsw6U/VqItsiwFPtD7h+PIsLBnkb0Xb
aWrZJERzQTtIVkccD8gIhST3gzHGAulB6eVUD2s4T0s7RC/bteM0OYNCzY62qRBClrckdplKaziN
LwJjheWziHmWLXv/EmEzvircmeHZrwseqOspNGPRn1IN6o3cuAFtFGTqcT90UVYRHiGFeJhKRTpt
mTu5pQ92+vI6FKjsw1i6iSvfxoa8yiv386uyTyn8pHzDOQGpRf7E2sjQSKFETad0DfUKndjNco4c
czryzb3E4mFppFxIWW4BLZIGoiKh5sAK1p2iaNftBEIAHfuBKpdgyzvwGgOC+jn4EYurgsMF4m3h
kgnAuKR/WubxBz9rvLRyc6U1OFDszJd6M2hm+nLGlZy1QyCMLBenjk/hjR1AZWfPKksFSu9FB7KO
g2Erhkoj9T6LgTcoKmuw+CVJ6rPdRP4GSKt1hCVSnrXu3D8edjAEsro5GtSHCL3L1e9zcjyXfKXx
XHeAsPc3yMt4mVTB82orEwr0CPz8Wp5LSEuLfSSW0DMliG4f+r4PI72XbvdE9+PYe3eM8K1HF3O+
jbMpwADWU/bqchVf/wD6w/GU2AqcIK5kTbwYW9zUpAmRTFIk8umfyDRWbOUEGm2dt7Ov4ShTotmi
inVIXvFrlmwmfXoUk/dbLTN8uTe3Gm4qRoRsTOeN5DNBqMXA8wA6z9GlVKXVbrzL5DbQes6gqlsJ
P95S84ksbIK1pCUYfbny5agcBiYIfV+R3NthsvubmtcbncYZgbZ1NDI6BqRIURtw/oQr+jUtSunl
o7e+htbY8+yZLnUbKLfeSlwBGyYm1Avs5L0099PB/zaw0nqjh6oO/T8vFz+yyQsqb8fnPAiIWKU+
xA//o5tn6ASG9XREmqGabIs4xMaC8BvgPt7yd56s1tkEQ9+emp95ONaC6EmbC/0MYiDrCIC3fKg4
FDaIY3D5xgdYGg2YPR8O1cxcGKeJ23zl2FuurrLRnRRroh6L7cqUdJy29OGfwy60DU3XZj7lva0X
v5+UOVGYxEiEFKsVdqASwmCpV20QZSOHRosdWIkgtQroreAPfrlAgZor0MMITA+G9emWvwpPLn1M
tsI98ra9YV0hZ5OhZhY7N0LK3hPic2dXOzkCXMIA+0vwbc6EcFuaVz8Nx4HH1TxzwEJQoUTf2rAT
BOmYcs76VdV01I9ZfQu2VYOW9DsuJt0/BTXU5+DNbLMpRgi5exK4zDmQuVKWGLFgOX01bAANPuax
i2G4/l8RVu+xsecvSlZTwZ6nQw/mcVneP8Vfu7LEto+akvSz/W1KwUlYkIfUCt2zi6Ye+zQNoxzg
CbTsMejNvS374G5h9r5CfkEogZf4mSTT9/u4PM/OvrOZouHkAnq5e2HfhxzgIg2t5LECDDHM0G3P
U2kZQoNAWhtJj/1P5AedNHHIoPdx+7S9aF9AJ9+zn+5DB4ZVQSf+uRLiuwtv52z2rlpmWPsBR2w6
56H43hlykIt7wrXE4wuyn01Yepcq1VZdj54DMaN97KSP1+aDzuomitiglgTQ4jsuCn/NxV+2lA+y
8Mtou/FWXSCTE15oZyeQ89fEE8lnQGQp/Mps+/yOX2nFdTSw4VWACGMlLpkTpk0ph6UIL2fEnNa4
cmXfvDhTuUAqxobZ9XoCdxqZo+H6E0EX8Of0eUtV44cCL+3ocahjKONdCIf1o/5cUMu2ioKO/FtZ
phDFnRwoPOzkOHAR1IqczNIiWD4b3lm4caRBHcB7i02Z5L2MZEViycrbE2n7RC8Km2VS6wfILwfP
u/uEv356bFkyS5G3GS//BspSNnKNdo/fxz1J0yoxAgRwxqBETxVAYi3rpDgm6OQr21k12NLMsJto
3DRfprggKu1ATMupLaaNxDox1xEqhQ2W9C4IszfO7yRWuFW9653DEaZwmu254Fb/ORfgdGBZ47Np
Teh5FFvpDEo9CiwgkkrmS0RlogOpkfOeCUTtCCRRJDwn93iHWazf2/3huU8gTZfKXtzeG87KhIoz
0PDnDSGrBJC/DVrF5Jh/EMTHf9TwsJsvFRD4higYA+K9hG1cu9rxteJx540Hz7R+FWiTWWazW8IV
+2s2ORAXxpnVI+vSrzDqxR5h+81nR6rMVMaRufCxG3vAJh5uD7rpKwEpTS/qmDSUc5jgrMw4wjsd
k9ShRvCExXQmR+h3Ks+f6WZXeQfF9SRDO/S4JkbJr37N31fyFIR4jPnheU//yehzRYVRN0EnYZGq
DVBCUiV8VRGuAns+wADcfdDLBNQQYsZ45VAXHIsc4+wnRcTEGnB+CDGbDCXBda9TboyesIQcmy0p
efL+hjghoUzN7gTPfqyAsHPlkJxHG0TKT6hw80tDDRMqFmBmatDaWVFQ+prg2yXWm0689m95JWLW
cLrnmpudgi5AuVmbVGFEFqWIwzQcbGwPqzN8mJI8gicakJ3S0gKIOca8c3XVBzOAEWjpvBxN4m92
0wpySblQf0VqynG3Q33TVS8zMPwQ1cKPBswpkZDNK0UDpHHjosLIulyXmKJ/Y5gxpf8imEad9EBu
Djxle/qdO6Aq/k2KPsAxaNV2JkfdYW8h0MEl5OH002vTFaed6ROMF8Q5TLNTXSZytv8HUpahJ3vg
AuobBaRZNDH1RT6gtPQ+zVTE0twcZd3/7vZp7xFcMoj8kIyTZjM/vNbEaUy7bv1YujyHnU4U2NlI
eaPun9OiSBZ7407/L7p6jLxVto8u6z5oDEbh8jGDyeYr/BuMwcO1OFVGBo/tuWqQ4XPS0ACcOT3j
ABFV4xqXKm4nJssO3dIzkAN7OoJllKDxjQU8gB4YvHcvv4kdsX02qIxZpH5VDNxGk9k6nOd130E7
2EVLiJRm0R+xLtKhaiFcZE/B1qZSv/s4tX/pFh/56hDGRrl5A+60pFwoP4UhP2Glde7YOeXfZlPZ
OqJMzALE4pb/rkMwtQfwiYsJ7thgVw9wDbx9Af7hPAf0FbjzGz5Ja+hgUSCxGekFhBsUXbG++1eS
QvcKblGpSfQwOIdFW9cLr5HXgC15gwZqpyknOiqkdpPKYFjPEApC1mSrNTFrl1/QcSNFwXxEqFBN
CzLTKdA2zQlVPp5nSRaopNdHdgEyUuZmYsatHDKTF0vrhJC1s02V9jPZRfX6+5EcgdyBvSz/dy35
gzeN0Up3DKphhUhvw8KvesrY8WV+zNiqt/s5+zMXULTvlADTeSzVLaBWn/nf9MBNBMC0XJ6BZyF4
xFDTIUykRs1y8ddZQMNZHPPr27aUGaSOYAhR6PXTauvlvDWm/JtVg55q5OA0DwUux/fOtI57WaVK
QT8d2aOEN4U8rz9cvMJEcWiIugF8Vjzm0oi23LxLjy6spGGvPlDrfhatJvWOP7mWa0+TaGbZbb+a
fIzOIMg090GztEq0uynC7ZakjgPzYWMbgwxBuy6d15Coak9iXR9bYUvOigNr4dLRQts/zbPqCMz4
i3JtnTOX29SYGfhNt3OIIOGi/of2o+LOhQE0JQLkIKiqgb7BkuTgTYoPp8GV/mQAtW5x4MLT+zY0
AlByUFN6CJedmWY4e6aC2MBQ78/NfP0PPelh8XkfcF3A+xs1a93RojuKj6ehCQ+bozDMtVz1qkmQ
SSuS2aakv71wBlSJEawAIwryfBtFYnIX4+qJAPvltoII295GnajNfD4LXbK9ngiJCsMNgxik4d+s
u9MZi+/MnhJAxr+TwsKbzkY7DJW+UwDqX5YnY17VgdqDwjOB0YNKmuyqtwy8uNI4AovCh7gy+3xb
1wsEJhGpUlTkmwW93OGh31p7NRHl90MHq4Qm1QRr0oBUDPV2E+xazNvrKSPMRZFwuPHJ8W+icZ2q
zMPnSLR/iDzlesZeyfVQuyfNxDGOFlly0KZ6VNawKEV/8Lp8y9vMR7P0DORsKjwMnFSUM0fzF10p
XEnCwtU8Kx6G8kZpBw8Lq5YlYcTVa8RTRBchUDIx/NgqcuUxWMn96YKYB1vCLs+LgfhAunlSXhdR
8oZq34+h1xxg/pe3R187rZJ8aubBX2pvft3o+CrV8dfAna5RV7XwrkZdfRFvtF2uGWQoqHT/++RH
CNv5TiU6dhvMgUue/PBP0u4wcNz3BebbloC5icFY3bWF7n66c0O9YSfYtiHqNQk9JX3XvJ7jWFi4
61JinZUMzvpT/o/wNIvyaSzwICN6bIxiMXyc0+4lQS17iI48r4izhL3WeW7dBv91QyaUlMady49i
jMZ8VglO+NbuYGxDNKKbMu11FwLZ2mHbDJP6SJ8q3nPBAiwoFYNEzBmG/T7jcdyrzXTRV6qS771A
cjbNaKXL9pW8mhMVbIvs7k20g8SRMdKwSzA/zdflp75HXoefUp69gfFn0O1WKvrQMVKEyWCe5U/v
jjEbvwXu98SS6MV3ynwmPzaKtkWuCFturEE0nw5YBSVMnsclnTSeI2VCLG2mY88zXXq2deZVJiLR
0FX9hHebMWbPKn1crAmDJMpYFAhiO4PUKoL3/7o0BcKm+OlEtLXgnP6DvuF9iORO//Pa/kuyuVMQ
wUwl3eaCmg56URvVr3FO2qvQTdFLkx1japM1babncDQsU+m9SZ7JWx8Kr/+GgpAc3msDIC+7PHLf
kyURf69tgHcNc8U2G84ocv7Q+g86LF0VEo6WmY2Z0GETBcaYVQAXAdJM6Ax7FtUmRuzI4ZOG+8OF
wR8fu7Wavquxycnv3Ois7o8iFBYQHp91LmAokQFCiXesdnfx4+NHxVilQyWCAc53mvTM1IzE6Edg
chPB3UjhQbfWlkyXXAMWq48H8lvQtQ/bByLCANXh5tgl/gebmO6e6kFe9r/xqyxgMtGtEUHYzZR6
O1jLzV9BDMckVVqsdH/4IwivpDvG7cBQXv+3vQc7NnVCRVV25Q58iWImFOi/h0DE9vnxFouF3ZyL
VtIefiyBjLZO4fo+Hpy6FJZp6nGDuF1XwooLAxQNWZPohfSYHK4pBqMGtZmvbd1Kbpshn7BJwdss
DfFdDfjNWK+hhxH3Z8R/gzLqa/EaPtcV1dbBaBJjNIEOtZm0MlR4LBZTJkVEv1sajiPioAHwf9SG
Hd879pT2KZ4CbHeEdVxgp3KehqVj1LLYqZlBlNnVwxx+f00ZdBgWLlckiHFRHkpI0v+eVEbfqOuk
nWPbdzNA+/eTrVBjMTEN4tWGdHPLCFfOaYCrHpbJcw2O3BSqajX7s6ivWaT7zBFgkL00bUaW7GKV
M1jOGcoViJ5OdOpw/6n+NjIMfVYGVItRPmvvtZgVOVjYAlH8Av9CTMRrgcjrzJ08Hh2Nmd8Mi/b9
PA23qegWwzBh4wFx9XoAqY7mnZQh+4+EsvE9vQFzVEyRISVmwXo6JNdVf+Yc7KS1uFGwCFA/pvtJ
Ieainme7aVaSrcQoqmPZgrmcWrk06qO4XxDQ32niarJNoiNu4EssVAOWYva6pHHT3NdxLOx8D7MP
A+6+/JPzLtHgDRLxS+RVSsC3ma5A0/6uHHcoG3GppBACIJerZsP8Vo8TRIxQ3frBifVOnJNK5JP3
WBjGboW8/fC17KScvbv2nHSbEWTvtmqojQFXih97rw1FKduRQ6KMu2HGyh+eSF/TX1l4p3iC7IZ1
jiSU/8Sr2YW0bmJQZbP0+nRb2LfH/jmOp5EdIGeXhR29k5oIKSy39px/lbsKxGXoBaRJfuejI2+t
dEPueuuQvBdxUreq5J6Gt+nHHA80nM31Bcw6bzjCZEnXa+sswhMN9IUQ5W+RmVcxlhLO+O5RZ5j5
fhWINnapZt9ST+fWRr/lOKeJ/UBZ+/+o8QZY1IrEgQz1MSI81yLV7+XUllT6SUT9ulIEUF6QoDUd
10wAfurNV2PiG7oaQz/kXnf9qLbUi+scmwB5dr3h5VREn3EILH+go6lmjdOxAYjOgYUVJBGExt47
0BeQCDjkRabmT+1Rbk/movw/OB50QUfYUXQXBQ77s4dAoMps2z8z7D5EM8br5jXS3T6rdLj2lTWl
LbXDVlNHYuidaYwaUBSmTDoNo9UcA56eIJI35qHo3qXiYf5oaJpHZn3CTndapxGOpmEm9zD5ktXF
aN+gVG7zMJRf8xn2220jvpH6PqH3Z9DI69LUOJF4XMLKEtAlc71pN6JMjFT4L1RqV7NRTqSNQsdD
xqCmAm3TXQ8QxQbAuKrTWQFV0AJbQvX/C4DvabQFShJSe28+LyfuAl5i9saNgTeNFfNOB9T6Igh3
D9tpxIz0SGaxNIETKDXIDSTd5p8ny7T3gVf2Z/dxluNV5jviCdwG1R8vaqznnzy9nFPzmZB8xrVB
48AjPyHxZ4SMuFx0SaO2Of7GrE9QCLr2RvPXkRkHYOpzc0cedoyRfcy6guNiNFLzoiycqfDiFCiX
pSV1f12p13nGVh9ed7xru17cErCYySiak2GY6Udv7hEtM+bHOLHyFWsY4+79p17IeMI3Q5ONlMtZ
TFeH0vgiv2sBeRUnUo+89cHQtHAX/2tWD5D5weodqxk6vQ0dKsEtJNIyf0u8/hD1VI1dd9Ipfhdr
pNPBHveHL44QX6204LgFqinlmUCOW3YkmmZ9DmA/umPeGAEjuw8KOtIaExqcKNn98LJDt/TOASjr
91D6gad8EbqBPoEHQcBkxgFSKq0IML8JnS4hjxqdV2z/M/nnUWfGG3NBklWfKOHP2A7qylR37AGd
BEk5+0kYm12/jDT7cPCQ9zudZPFkXZxtpMXPGb5h4EJ5buJTEiMjF9tzyxyKryMByZkvHFksqptG
Sl9UZharruFMWA716AEyH5GP4TR8khH6nret4hRQGOe6rpcmwPKfZRJuhDXKt2DDSiO62dtqFPK8
4KisRwwonbquRStGojfg3qRmgcdFFQUBFMCoyDuG8osmzaVpSpcSaYiNJeST+uUoqY4f7IqUVO7R
CT8Xf9JiaU5f0eYr7T2hJzXXY4+BVNz3quqjMj2z/tevMGvbbcfjb5NvQTheODgHELMeMTAjMBqs
/zCkb4BwAY6CAns03xxa2Qf2HCN/pERYegH61n5CEz7/sa8C8LlDvpxi0zHO7oQEb08iRxPlmT2k
ZEmJV7XDIDiq3Rzc/dquFEPoEm3y7Kny0Y2sLk1aEqNlDzKDvXcEiu/BheUF/Cfrv64QwHttcyLu
Ks1vIefBRDJ1w/mO2eYDduHQwlTpMeFHbrr3+iv+ev6w6jlTXTq3xqeXuq+zRhdLXPa5YsdzVPcZ
QHDW2BozMUknHYqgBHHa5Dax461pmLbPWcptIDUMVszjyEE/7GESXAJ+Ex71QVzSJI1ijze1po5c
T2efS9qEkWsfBpWRBk3JWkQY3jjKqeZeefsCdJcGyez7dG1ibJcIycYSRqQ1MErxTLI2qE1dMzkG
PbzA0h5xC35LY+rQIRA8uj4nwcTbPaqBOLbC7PcZ1UaYMCILRZaTRu2UCj5GecbRO7YNxTIqTnlX
O97eAPFSkmf1QZrUeOFU1WKd4tkQXCAn1bpecQl63i73MMG1YpZUrOsLH4fXKFqY2+hzjPAEPW3Q
4weFRxDQ187yv4tpwKzLvfIU17zEgp5iUYwDSpsnnxdf59eV1WvXQiqoOYkQPCl+AfLjv9GznUWl
QCCk++JFNwSyYvwVC6HTQ5qvW0MqhPzG3IT8q1Fca4vh9wV6D8IPBzm7aI2LlZVADUBctfwF2Mtl
uLRvAn8K4C9n2juUQ77e4fk5wLKNkdSpo99H3MaX3zgjfZrZiSb9M42fonjRGnXizvCaOaQR0eZr
f0yMUXaa0G2ZAtsNYaKD/+H2tx/S9lj5VU8wMucXBMbLpFQiF0VTy8nJ0kygoO0IbUon6sXYjykl
anWyHMiYRU4FgpwQCDLe0T3TjFVbZyIl3AF55n9hBHn/h+9lOn8OkCFASvQjJvtY0WxcpWQbS+UO
AIZCN3f21RabpKgtHiNN07Gz5j56+A3GIPTXpClbm6U48H3Ulve14mrK3mWrPL5E9gLltHv6nD9i
vTvpKiu3pPOjMOC6a0+9BWUZbSkzj2grD8UIFgkXFBfOZ3AuLlEWX1qMCe5VNrZnWQJTR43bfVdL
KY4kfugoEda5KjRst1D8Szw4fUtDg3g8qr5R7BVnuu+b+Uh49MVH1cajoLmNwjz8yGti+37MEoux
Z+RkFy9OIJRS0cRQIWj0dDMt2YwseuDBkpwcAbGhDxj4gVV9uOokVgnK+y7oTxLm5skhagyDwyr7
xxDC5gNr8s/dxLBCoT5HoXTnpBXWwdheqtXQb/KoyYkaL+1TOzbsV/qf2UxIYiKbduwhc/Xj3Dv+
uWwVeJ8IS9R0Wl4bPVHnZ6XowEs6ZluCxkJ6j7U7Ec90lAVV0hcWCUNMs4YqN4IM6PoiCXo4UXOV
UJBaxusK/CqcIfHm+o6kZS9SjCBXvWeqkRfnIJ5IVZmfmy/G9+sMrxY1iT8+elQGjWXkkSvMNpLP
3SC6P/Oxducp9o7einiyJMV4ffvfTyyN0ilvpdNxkXcUhsx76nbMkgrVmdIlixeWej6Cm4hOUP7T
bBDb7Gd8AaYb/IyyuCA5w3JmqLWvuuLD/RAjpciCXXPrVgsE/mbkzXInBPh9iuTASp6AE8Kk09HA
c07crNTzBxsOwQ+aS5C9o0A2Lx9nP0kfXuiSiAHm26Z8+1oDEYqSqm5TBHI91llBc6zmTZq69FLq
3rRQlJcG+/6Esx1J9pvs7zWcr4mTxaPAw+j6VAGDL3aChxL7s3o6XStEQ/jSrA7Hj0t6VKEtpGHR
uMd2wRxfpx4JZ1kl1aVoLIZgUxDLYx2A8zZO89Bo9Hvik62rxW2Knbh6fwLvzL8Dguvb3cy8NVaP
0De9ZLF+U9/9UdLQTZ3voe0+bRZIYofBwYO31Qh5773fgZu1Fjnvz4RBhik10nHmGFZkjh6Kb7L+
TCtP+vcK1mG35XuYbJQxdG2lX2Kfpy5+WBPvSV/N1sPgqAqMQHvJZokorCYTB105E+mMmkw7yQow
3qT6lEl0mfnZC92Ysyk522f9tkZw7+HZIrfef94iW3RI8tOeuSQT4Wg5ck1cMZTiRWY4dfBMdxnC
cA03d1zlPlFEqMPM+mGyydrCxsw3pGnJpYwvO0y+NZqXfY5mc0QxfNMVh9cFf1+yyfK7X2USk/2I
9C7mhqZpc1TgOJYDRFtpm3eWN5SH9jn03lkYuOn6jKCIBIjfJwZqRI4d9ucTrVicmmYC85eLf/dG
5itHFZ9SZTV9Ze3F0MGDY9ReHXmFAZ3yDF+edrZ+e9N07xqTev9rBuQ/v47d5POzIIU918jW2IpB
9C3azXwI/gQ1bx0tzrzOzoRFJIrAFfe3rZnsRa8hMDZLgQWr/TvAadNfBmnpPU1h1wAQLXtkwqwZ
AiYmnFbUvhvtmMM+CuLAt039E0ByvYuuoT2w+rxZDFnT70Pdl+7w0LiUDd6Px8KpND4dexxe0TIt
E1UyBFpnaopngOxmXb5CcKOUA4k+Xcj7gtUtxToXgjivhKRqmIB/pidveNekU8BwF2QJyEikKl/4
RHnbGbu2M5MsTcd0rLB6tXyLEUIu0v8vMv/KopvV9b98xOuxx0ryr0VZDQmkpqviPaTvmjEHrA5K
Qrmn5F29SmlPnMquvuVJ+FPokGRmlJpK3J85HGgjYmZNOO7tQ4Ip6YKinY0jeyPflQX1uuqQzdPG
oYZ9mme1Q44zkPsdVe7JOnqQX/rJtrHLWlPTMKtGW/0Ae71axD/tUlAIygfwal/VzYP6fQUvRXlo
F9FtyGPEWMx6GKiKoEBWQFIQYc3kau3kg19/JautRl2WED0tcRfaWGt3yZ0KayhUJUwS/9NyfcVi
omWLYNUStHQDKtMV/3F84wZdku+vjNfZGWbTqlrRaMHViUgElspmPyulvfCoiG0WE03eEfCm0ARC
/lvlcxb8zoPG6cE6dlgZAGJXbMxG0ujiyzSOm53ENlK4Vek/ZPRJPUHs1eqgZWVLBr7kM2Mg9/nX
R+tjCoJnVAILJU6du9GWjFpRQ5fPFdF1UclP1yRqY2QPnAzAGA773gAmIWXqiC9BwoYsj0/ZTHKY
FqcxeFjF+mlD2/qJjNxn5E/MPeoZ25jpwFAlbiRS9LNThSmE94H6L5vxpHMK3CXF4P/WWqDYpG/m
VCjHi40x88m+UPPdyr+B3wXcQ/bQt+o5Hi3NFPl7WE29O2v1UWqWhmnMA8FAtFFWUobXXXDKouYM
T9uJvQN1ZQOEW4ecfd3ut6oaCBJzWqxeKMkBzb7p8lVdWV7Ws36b/nDX4iZxzZ0YmC0yGJ/LKxV9
Or3WDSA3/34xj+O6DVeeLCyOMREBEVLYzDRhaGBN+KQJmJiw9xl7ppqfvSknNS5ADcyJoMFbOgk6
kip+CYdhj5BJoJocQdYH+HvHyCY2KjKAl63YubqoFPNV/RvAVQkXyY6h3B2Hco1zo39z0IfRR07B
P6TA2d3puBbtPlvwK9W82+mR3PusNRrxsj9YCWpjSMerDbVG+EwlmhLNP76uN8lrI9mGEbPZvNlO
uhSnQe4uKYAXI00g7lOij1NXR53QFrl5eUiiItLRsqdfHqifDNtKaxoR+fHlLUOM5bjjjj/5sNmy
VhslJ+7yDDRf2g073JF9rx8G/Qb9i/6FGKLNY0MUy77P67YufwiKtc8hJ+dRB9IxMrqQsVDM+oB+
RVlBzfOoF7QhMHu2LgVpB/PKKEgKUO2TrvRonAyq6dVV55jyo0Jo+CiQjsr3NRZSe3KDsrDoL6Vl
Md5m+rwx8sW24c0nzoFDmyNDaQMqONEoLh2+LtpHAGc97IeSDD43mB6XijsIljCg2LB+5h8RPhBr
zFcMiR3QMlWdziKe+5YJmGMWJv0TXswezDbx5U496iux1HLAfdvmy8B5ppuAIBvWedgCuakupPIe
thLurKvS6aj98Vzz56z3/p7ihl+Bi+/ULkoZnZrjlLbV/UPs57OujgZdQpH6Sl27u/53GyZuFplz
IUNukMXNNRb1WImgP8WIBlVbXONCFIOottij2A59x08wSPVHSft2Rp9PDXbyYM8Kunbwq5KzdEaR
LnSPEPUJDokee/2H9unZmEhiIOrlmFe+hC/VaVg2v9w8PRpB8KLg6XJfezLS01wfivsnzDPYo0ju
4TcGm6tCzutz/9zMJ+iGrX7mkCJeyY5QdQSGVrVlrkf8OH+XwVsFT0zRGD91TzzpSt7lCcwDfkC5
XePtiO+ixK8Vt+aXTmMggCnbW6SOdoYP9GEGmdGNCb5DKMOJZbRdC2ZcktVjtCIfLCB1deoLWR2C
CJN7dN82/Q+F1Vr4MuCUbb8bbgR4RgmQjHKP9GLgDnqoWwGyx7kXRnwNGNJQTXjkPFYFaFW1P0rJ
xY4gMTRVc6hCBiKdYlAAsWyaqlTAZY4XqDTOQN11XHzW43tEHFk4u5hNsTYWBUt/FUhtxojwn7GM
g1ADdfWySCrk/Uam9L4/0nHDGZ+iG2eMwUMLihnrei48fLxIQvclnEWkK86v0nWn4JKbv/uuBsid
gcCRThN2hUX2b6RI0Gqy4uYpV/tda4maXyfPuadhhhnsZcm2u6R/MDv4qpKa0A/Fke4iGDpKKykA
WpltsJeN0ZvPOg6LvvOVWiQKahpT70nsrhhqOu2V3xOElFmU1BHV8SZ/+AIrEhgOGrYxq/a3e0xS
xGtdXfalnrd/Bh8Z1aBzF1BI3sOU06AlAMxBRs+9D0Im/X2VbZ28k8AqNRLjxc/Us++OUODpV8sz
ZVWqzUu1ikyOVk7s6wIhm6h+E6vFJ0bUkiiAszL0xM0Qy1RnZe+ssbwI6Drh4HUoHW8QnUY3ddTU
1zuPOg305u5wTewvFr76DncdtUl/v0PEk2kwoq0eTxX576B1Q/B//NjriGVo+bhcG8yeqzKvB8WY
SS3s4HrdM86W3dep1KjAQrsr0Uf5OoEtZf6r8b3XqQPF6RZGYf7+BWxyyiD+No2lqgUBFd3KrWw4
PezGitw8/SckuOIp7y+F0QYu9lJZZBpQNhHYrwXKEt5tfUG9URY4aV9RQBlImiv+ju3ThssWwsQ+
IdbDepzL54zzTibyZYDKM/OVK0DKEmsJSNzo+8lLriXODFnYgymFoQPogqaiDVd0qUxy7i46oL0N
raoVw6VF7OfSP4BVAcF9ZlTE+B7cBP/C2ifP1tCJd4mN48ACmOJQTjgEprFl3c5TWiTKojbx2guE
Tp1rHrUwo9mJy535sUfpz/OM8dnJn6zT7Z7Z0flIqsFo28xpe8QxAVsOjx9nItgYowTfborQCyS/
z+i9IZM2TvepWc4ZLpDGbs8LELlM+YY/yIOCFsB+WfGdiA68XQPVaZKWKMdqR1Swaq77WKRE315n
krXLz3Fqq2IKqiu2AWMaSbjdCb12gP2dchWpW81lMIlvRWaCuqQ4elDWOiVcHfPmqe0DYVajkWhW
jqgOdW9nF2uArJb9sV9Ql3hRSzQ47MH12AvTHfoV/VyS3WoNaFvqJdIHFXslzRiyNS7HnIz+bL3b
X4pCtHowyDPK+iemZdnMHlJjWfTzSpOQI9Shg2xo04pv78RFjN9DP0fl9Mrp24H7AnxNO0eFBcZL
8HAQbhKxHpXqIJnEDywB4lcVWprcGBVvfVW6w8zMkY0aeBH21Idy0K0+GS9qRF9XxbvZQ5bf7p8Z
dEL4fsYrhgFIZr5Qvqh3/Os5+S9EUyi2qGpzLnIEj+MxUtgCE2NRuD7JH6lkO47Ru3inVeTOMQ60
dsfACeuhKHF24J1n5m42hc5AWtAarpFaUbKDhD4ZDLOVIzNphDRUgiBGRdZg5qmbY+P1eP5ntPjf
ndrqebOk9GdLPMCWaIZWNrAOlBwMH1nGKpKdUxGHIM2zD64n+iG/Qm+cM22taEZ/TV9bkVTPaurh
xPvrECl73xwVL9UyNrVf8HDyYsH3pYuU2N1sAvPexDBqEtzzciA8bWLu5U/2r+Pqctt4uqQzUw41
SWyKAwuGWV7azWKSDwBsoPSotRc/kAclMzSamWb690Qn6lVmg4rj2kQNy9zMEVXg8+JWl3XgRoGZ
KJlmTz8aKdB48tZfHGd7+zQoySeDDUSRKK50mRxaMPMAY1QaYgfUpjzmj2U4zhyHRWSI42CmucUH
umYBQa1dIfusODr7xfEBH1tDMYhfKuohHMvhRuNkzP3pUYCgUWsQlLvW5WN3HTGgcdVIROkqPh2S
UKcVm6ohm0gsK44LNj/1sisKX0yYDimSZlWIC2I6UQAhwJcFaSEn+w4rQNJExqLtRQUY0PgKMwU8
HquUMS8M94aTkkbCfjJX5jKN8bVqv9vM978i0hzJy0s3podvbgsYwaQqmo6nba0hUlnDjPQVI1n9
G4qBtYO7WOr/dPoJnuHBV+i6KPg+jUlCeUC6fdq4/xfoq+AcfCLjKqqRufzcPGcHyhRL6l91jWIV
p5N+VsgEcqHNuoErnqosV83xWPSgF1HIkbBu3WTeUWfhiS0rzy2xOvDDgcy8f/Rbyh4cIAuwChPj
sz495u/ArFNZlN6iSiLFE3Kbsy4tRU+iC6bunrehMK1oB2JVNTnt2iGxZzYVyiGVccuXAwVYA2+9
1cd7vJpfRWYU9RZVUZ6h+Z6F8Uy3dFhE5R2oMwhBPea0VBc3aufwT1O7S/7UYVphvoR05xAa9Ine
+0NXcnRjUBLPMxFBjYmn3oG78eiucMgN9fCuAR7t2zD0whJ89mav34x3bRyFDe8Asc2maQ5Jh+oa
cJdih56iVMHUqKfaoZWYMfMyBtvCF4g3GOOzk/r+PgQSJEixcx9LJTlyAwFZgJHAPxz9GG4KYwpt
zbkRJq3JVgnzKCVMZzjrVLZaX5zVPOvvxYH5RbMB9Qu1ciZt57ONeqiqVXGZEYujbr9YPxugl4pM
onuNTcLRTbQyWYFjdX3x6QvZhWzHsexOJykso+mMAiMdA2df4gtw2dfA+bETPItEjkxfapI2EuOj
4T/fklqTqiKagncXP8Eveew4Vk8K62xUNcAXyBB1EvwNJHo52tybQhFFucRhESYzusQiF07yb/Lj
EyujyXZiwy6SX6LdOHiXCejJISd4rS1iscsGzvmizMdblcf9PJPBpBvGZkc3pU9udrQQe39MLiWb
vh6rXKWWwNRkTDvgEk6edQ9HLYag5xIJT/ZmLRWZHBniQMroKX1dJGxGtWeEehjDxpEVq6sBQN++
q1C7k1u86oIQOGKTfSTwblyXfaYFdmYsUM2W67Qn7n4NvfocA707DUc5/VGcbOAHZU5QB6syoWjQ
lzA71QX+Li9BFTGeMlIckYimjWd+p63cjdwhtq5cyWRZSXNW+BQtyHlkeMEuPnSb4WHWtofYALOy
/8xzEWSdTcq+nS0ZOz5cr9alv7UgjZmWBg1cLzqrp4G/I8i2nr35/irbrHMijMIFr70J+ENGuLQr
RaPB5cxQmyT0fG4hpJ60WjqYl8+1xZlEN7rn1I5KePzh+sUVoy7kBeFWxhZihUJf1XQfgWKxlMHY
UokN+rc/RRHMRifOBuUNaXcg1LwbYainEFUWY8asDRRTKkd2cngX29/nX9IIF3wyW84UsOdcmubO
PrXTHyfQJDO1ImZLyJUUGO+Lg/iXlJdqvlAdow5vHogcA97kzvEaX2fWm/avJvi9UkdcYZ3fhpcV
8qxjd/Iiixyo+/t5/stQ2dDTKUN7v4B0aJQsetw1ZqJbMv49pRTiX95i1eX4cvP75X44txH7TfD3
I1DqIDOYFutyMZYeql9tzIRvu1zw68NlgWyxicCl+96sLfeNklyopmznX68qVupmtlcz41Jdn+MB
xGVcqLhVQa/Z2hHJVpRH6IBdfwehkx1GzZdP3ZQEHkx4PdgoJqjnRBrVsb1rvSuUVjCaX1N4C7Cj
bEQF0bs2Bm93zpEzRB0OKN+QWV/sgBrX/qfqWO0bZKJZRi500WeHwARakS42h0uUUHOkyx4Kvftk
PR6JE93M6AOMz+4plOeKT06gro1xJmNWZaLdzso4fW41W5CEdR0zJh6yp2BWtuzP0Qsg9pvFVZEI
xoGrVBrstHBbxxC4rXx4K4J+0T0CzVCfeFFyfr07n3gdGi5WEQvYPr+WXrXf7CiQmfgsRKtTl6EJ
ZeCwxw7OZn7hG6Nc4VmiH2Bh+CjBZ8hCG/msNMXqnbtDWzkocoM8hC8fRE/aac0Bg4W7LIwiB09d
lbMZKnHaQxzY5O3/eS9nE/A+jfINefjtxI7vUl+EkM8mUCdTr0AqFDGs8YmngYHx9UqZUQgWwN4+
VaiwXcmZJZqc4uTpYxfUGMjpfMzJc4NsGAXmoXmb35NgLiDi+/euCfZ3QUxBstN1iUQpx2fO96Yt
pKCiH5tJyBmGJK6yHqjacZQ/fjmZLhY/4PwsuKUr5i2C+G/VtzQS0Qe5v+pibgDWQ7UWW5xN7kQd
EWRXmpqWFjeXF1GUmgSN3+DQT4NzlKv+P45o+0t1p0qCocs6nU9H68p2gkTG9tFkFTNqyaDeBre9
kzD14FeFFenhBS+jdnh7Ytjy0hn0AaB3zIpH9noL7ncDVzGaiYbKSHe09xFyj2YPYU8co8OtP5ZA
hqiuuAsVwZOA6W6h54mHLIW0oMB83uadaNf10bKsNykS6LF01hqOB+nD7KOKQBC3VB5zmkGfVAHT
3WknqGATUAPE4bijg45Se3JfosFNlgxwePVrDojpsZvOSCPRqithf9Kx1CPLwt1ZYWH9axbsfWAK
PV2o1bBsXirzTy240ND4C3hA1VKtcDDAhgvaVXQfIX5yo4sl6cU9+zVh+EDq1v22D5HxDlr/MO0h
P89NzNTxPCkIw7/gwML9Poz/fsx4s3nKJgNDbBHVey1IB0oIOGp62NnXiIK8w1jaaAsueqibseKN
MI31sycLbKrVgzzjIBtMzYw6QUTcOE3RhRKmdY5yd8qisHOChPqy4NPVOuTjLK0azUctrqQcolSC
k+eLtIdoy9wYwvw4CNyU/FLDjfhHejsN7Jd6MMbnpVWVqCE4QwfNBUEoAWSMZSbSZ7h76MqyjkwH
qsuKMc1zN+BmjGu7kzoVPTEBtKYy5NmXQU8vMl7V1zR7Hu0qtE0j7mUlovhy2+fUL0OypCy16Ygn
ZeRdxHcKv69AdEuvM60nbpY+JYiRu3oqkcuYPzYmJVyLLxIhR/YGUxTzqjEN9T7XfyHxfyIk+sF3
Dyy7/af1BGomhrbFmcH5sfb9d30chjGDNKQwl61YwpxrMOQ1lAhqgG2FRFfyBa3b6DLC2rEnpmEQ
BWXcwDS0l06aqLsdfoRqSdJJ35ymt+/yuPHrzsUJXwgYCI2bGQNuHUp34B2HeS9Gsf7zNa97OXeC
5U1Mwax/AG5NEOiHP7jzK3uNDIJWgGUxwt6PqEIQymEvYzEgUgeki97Oyb1Exsx5CitN43Qy5s1B
/WWOz0sSPfQnXAxjYbEfRwsErwarrl1gfhQ+CoaXwhoWpazH5hvEOAUGkFOyVnNvCT5/cSMRowOe
ikWtXucV6fEwSmgSR5E+/FZhPVC5G7d2hpgvYfk7/Wl8f8dFoeAnMldATDY8OPY67gr6DKWtA2dM
+p0uF7/3wBS5d72bzZUdxVxaNQ1m8Tt/81HA+23b1Z0YW5nhnM0pxQ8ObdXExqrcztDhLyiSDxVQ
/LJ44oIVvx2tfyPJ+xru8wmk21O9Mez5++/umYH04hnpIaJJW7n6qgJPZZU0yIA0Ms2YN7KBnQpo
UNZVE6jM7cP9z6JqlPnhx6RhSa3BfL6IvVPAbxICLS5YRPPNlh/+4atVwPkF2hTvmfztrakMUxhX
udXYAPWehOYzXWH8WPAQx8vhEVBouQ3FdDcgCwStEtJIJWF9XdUPGDij90FD0W1YC3VgiUU5Bibi
Ka7uV41DSR3WXidm6mQX/P3Ma0uGSyO8kSfqkxa1Ps+YxtGqMmqw51PzSo/GQXWnapRBCBTKHZ7R
bl65yV7eMjDD0JumsUqX0SFgcqLdbfPlp909CJwPTxuKbutHtZV/bjviwm/A4ujyUw73PwLgPU9t
riItjok7YmNvP48OO0HToiWpEO5w+WqrvyOCF00/AWVrWOS7vFnvCt6ZTOxmLtDPZG6mgO1adM+p
m/l8XsagNb+ZcQ6U2hZH597R3DS+ti2l9C23sJ1TkdwrLnHacrZdRurMgYnMrFB75xfgET1CP/SX
y56vqs9eWlDZzFHniUywvaFnungopS9dU34pkqFCz7rtkuvKyPXtUcX0rB5oZBE+XEVcFSWcf9WX
rZu9o//dSpUcGDlBElDT0YKwkpGi09n7bHGLhfw451ECfoKtT3EhOoO59gs92OXuwC5pjn1a44eF
3uWmmZrUKwQV9Atwq+N3jjCezZ+5AlQcT9pIBG4fDgfTNVCI1wbYNzefxqImzhGkErfSt79Lppa5
VoZP4qGHRwDAGPotlllNe0YNsqkc8mWlcc1roMULHTkfeolynLRmq4pAbRNrQISS1bSyuYrmdcfR
TtThIjL+HmRDT8fQHFdDXj0kU5crN62hHeM5fP2Ib/3/uonV3C0XE/eDEFk5v3hZKavDNJL2xnYR
QT7IiEGoWaCR76nSGMRod5+foMzT5fER3R6Uzng02xx66/pz6Vw8wNr8D9MHAO8gOaDwdUwF4Lzb
jKaqUa8XVGZ7d3F0hdJqlMI3T26cmTKGEvWfxTXvS6o1gDYRqtO/mcGydemmH9+j0kUwYurTjkUE
MndRSbaGLApmI41O2MwZiLB+lqu/iOGi5b3fwmPmMviuY9Qo5/++MBlIxI8MvIyG5NXXqUqBvH2V
0byz9G9dKHKizDuQM7vtuphbUh/8POen4eJIbtpqYjzzPXY+DpqBgrBUui3EHxh3h9BX3tww7zYq
Av4/O6feEpgLCYGrIY26g8NCVhI5AF6DwtdqnFaJXUvJupl3BAFoiulz0T7qL1AizrgDe6bCnZ/I
BK32zFZdQLswWPCH1TEsaMIdwqIcXoffk0fbMdS2C1iu0ou48BJR7lnygMwI2WVhAubXzTx+qNTe
WuN0g/chz1P0Ow9QuRE6egyS3Pcikyv8rceVsBIf9XF/ycOgdujGDANwQm+i3DoFl6s2CGD8mby8
ArhiKUKxtOWY8BVj5M4dNkErHQGGpYieVVy/USFJ9kjCcVxwIVFZ6hW8+sy/fXN+8ElKT+llPkje
druCyFjeHhZAeGZhX4j3aQ2kPnVfbG/PHWZM/GkIPpw+ousNW0PMRDi4Cxt0xkN7RoJx3E1yxEB7
7WVMpiZA/tC91hKXlAkxdEA59ABT7WSijJL1w41aPPmcKq++RGyaG2dQmbevWmayEBLiwGdEhHsj
sTR9F8VvojFVvTHNRNKMS4pUQ5g+8CET9/gAnpooXc1ZRMQwshpGiFBzHnJgkEPYC+mHMLlQ+tTp
AEo7gCGFELd9RzzYnvfS3uANVY2FAZxUoOIPusL7mhViht6EEGG3cZQQ/ErVrEiibtK/Wcvxi8mC
79bV2jfHht6bm7gvOjWyKHBwsQ6XzfO4tzxf0/g8x8AB9cb6NE1/hG2WjkDNHA2tfmRqn/cuDOXR
MP4XKzRD0cAcxcWsKL5PhtpGiC5zruxtdUIO95J1Edlui0SP4sVt1djl73MhEx8CjSH2SsgJIxnZ
Qb4EpqaPOTiEoncMbC9UaSxhkgB4/ppR1513n9noH7JpAnqLKdwmvxqV4P1SlVLYdf/mhhaFNeOW
I/J9+BJObK9GEQIeuSH30X66H+U+WYK7UufAg0mUUG+b6+deHKaMNSKDLIIjzAVnHR7H7W8IHB4H
EAMjvPAt10jnYraZ7q3LxczzaAq/CCpNLJZfIyn276Mri3cVCep1v0/diSgUpTZ5VjlB4QTxTpuX
N0itLmQLx4IeE1GfSodxXSu3qiyweme9dhsBkQMRFYoJ5PzH3PfMgCvBGmnHGQRYhETmztXAN4YH
l8CS8LTzxVfHLiZy9uAhgQLwrVhgFKRKgAc3qv6jMIX6rJKNTE5xdhrnuG4L6ETUju6wHMrsawXk
RDVesRPlHIVdYhB1eryjoOQEbOLc0YkGr2L8SU2P6sTN1qe89bxF66tI+ZaeZNi7YLdfIRHuP/JE
bQAQQGrBRdMfH+KD/LWAz4MueHoIV2THZ/ZpRyqK67n1l5uNdMXKqv5Tvs0tZe3M/qeXrJI8OyGM
6UhLo5h2cfiT6VI4FU4hRXckgMiYMQtcHHqTvpgnE/m4GmDa6WFtt73hkWT7mzKnXfyn8eQG1FOM
5FRZ2yoJ+sVSMokWZuxMLQN+D2oMkjRIEN/YTY6hnT29XE+UlYJTQcgnU9g77zEeXouFY9F4+pw3
QMeIvFCBrIfiJtZnnm5+jHolEJUJN32qkmBTa/ZDaNWZGgn9AZsdX7pxpJEpp4Yg3q1CJgapMDzu
V+OL6iO/YAcg3WzhaV4StcUADrFpNu2PN3PpEIIweql7FjAf6NhciSfYOjktBJCp+EcURyMqWlAR
1woqIea0kLQaTBjNbz3e5ICean69t86GuGgLxVLHkqDuZGbKUwALeUlLlw9ARSNZEtgLUWOYMUTJ
XVf03xYFBYM/EDgfCSLwhr4AHJt4YWLjRXLgJMCER1fAtxvdw1eU724NP8oUGEH7/4Li4mShMh4x
I2FvgVm1ebJ83stoOAd0+e5pZwRD9z+5g4ULgdOVqvgRqmo0WoKQuEhTrupoQpY+lJORc8aYt3Ii
nhg8zZSN2jsF7zMh1/UFeUJHw3eIEnOl+JIEt+C/AzfmRd6JX2YDSITYDlHhJzTUt4ZCmCZUyZkg
caD57O+yQjNY6jI80oNbULbnKa5AC+O4uub07/BTJNz3tQAKjLgOXq/e/0ni1WDzBIyxJsDKojx6
iM7dfH3EyYex1+YstYtl1rgOY4RpCl0Kq9VwZvueSsl4obFEcfKB55C3FCvs5D7BaHznuZ4nAEqf
XnqjsPQS9odZiSuRGM9HqrrZyjtyfCIZq1fWaVLSc+tsPth0bZoq+F9uj7ivxMekPNbNjE66ADA1
i+NQ553WNi5PMOAW8Sy5BXfDZBpAqS1rUqm6tDcsIoWM7rmmzv7WvwFTUeDt87dErpZ8Wfs/fdAJ
cFQOOXfGgnOHPKcDnnOt4xFy+seWP8y/XVY4xzjc8Hfa4+VWmAWYY/+DoplisnB566W3JhZHETHK
/Idx71Pj5mxOocUxQeunysfkBU345qIgcshB6GmsF8plg7Vxd1MAA2F+ylpGmlR39KlgJG2RbDVh
roJE1KPBKv/qE/en+SvXDnRaD9/q1mb9KDwpVRcYYZsdNiUU9xJniwz6TLqiufZBC4ZYf5BsdH9g
59Eg/RQh96c9TSB6r7rhz0gqzp63y9ZLBjm41SflPmOaxIqne/Hy3DEhsmiC5rlMoumhXAvF8Gpl
LnPNVenbEh9rDqZNcup9cq46VD6a5pNaijs0g1/CubFm7PxlBFTA/7QJRZH70Q1bjcP/i/vBS4M1
CMvgtoEAAb6Z5Wp9hJ2az5VNc2YjFwSK3iM/MtSfWp9Wxskzg/AG6Qxr8HIt5Isih2Aq0Uhgopup
o1Gd24LMuwCiYd/QXBqJdrxccq5791pCPCBmgmjW2qxlqz+rzRk+yjpZPpYE8f/kIAI03ZwnPIYm
YV0DuqVuXql69p/iguaQRHCfbijTpB3DHbqcLMOnfZwWLsVZup90nMWg4/QokpJFSVsHdeJpTvLl
txcJ0qJLcD3NDMNNibRtVsd3fVBPF3ENMk8nas9R/eKtXD+cl5XjD+lMb9ZB/HYaplFzM9vjM6jM
ZF1MUGcIoNw50l6+QoZ6upSDka1mfdoiGd9Cf7s4n2Bi+x+lNiYUw2fyzXe0UmSaI8YtL1fx/UTm
lBVem95To71KaM+cjAmtLiGjc23JuTpgCCV795nhSMiYRdMntDU72xihgFPtYiwUaGcPIlJy8A+D
Y2HuEln6qR+I6slGaI5sSvqyGqre01VJq5+DA6h2z4WUEA8tjOtAgQO97O8G5Izbl8bd3Si080wQ
bvfz59Wxbx+BH2DbvIl+hmD+bhRQsajWbL0M8W+9FeUXq5gzahgbcQFUL3PsRm6Nu+FXyIZkt9Dq
t78RyQCb8jmpbgc0fTPFl2xAlxCKj419TPSdYYd+D0mPPJ3mTzDkuks1J4pyHImsgaOtmyARc4Wx
7CYNvcsv7wkG4pbds0kVGZRJlQxVKOgsxgPhyLFSTPgxh6vBEuCrXCSElDjU9VVTjfiBnAbT7fPS
y1GsNA2PKGIJgCoyTnikVtBrNTr8/MkYUt5CHhM8vhfgnaAPM0nnZ4RVmleLz5jhdbUH6Kru2Ggb
oEFPLgmN2mlbXJkQY4VMcuH+/WyPjgBUembe5Is4gTtKnGiIbt6cU0uvakAioQHgqWfwPlbnpf+E
SUdWWbSf1K//GjsyEYPUHNp/aAZotqc+E4KNM34P77NfAwvzYj0z6wqbzBN5crWCE7G4vD/Fow1b
fEy3lQ3k8WSBBrKqRUaCBSqeb4QRIxVT5pYKRcApoei8kjFCL/LnNcv13mHO5mc2XJ9X83ncgckA
xXsZlMKZ1pFy///P9b/ilw69l+qid+jQCuWIYxdXVO2ZUghgkShx7eiGf9WzCXykbIYUf6aDWZZx
YHZ/pVm63bRPbSYqYFJH9iRuKYND6OvM6bLzEsO2PCIE44RAH6Z6wWHDyjb4xmIgdjiyKg2iMFog
iDoBXuCTXJ4qccw1iXm3/ju0YtgPlYS7BZ9TMMDzCcmKi9tNf6VdF9ldjTTZtbCmOb1irrxTQu7X
T/pACix7Rvex4u5LVEmhzO+I1xGNbWpd+5MChAyQdMtCDvCmUZwm7dZclcct4r4YOJMQu0bD/9BA
MN4hCG5YjDK+loamNgCJDUU4/Dso8MfIvtag3+zMEb6fVMy0r46WMPQrPh4Zsu3pCE3vtSeZ7Lfp
4+N7DKWB3p7rHCxvh/NWx6bF3/WVshVeb6pfV9YLzjeGCXGLgU1dfILuA8uQ5IZ4yCy5TdOdf6cU
blr44wK4DyHgIcfhhJmBYFoecGB4CxmmMqPVQVifgs+vu4acfewIqPhuuLBtcaAGEUWtPzCsQ+cL
zG7SZKpe2MvaNH8OqGxdf6EOObJHOhHwGnuRkJYQGJcTO5eJsrH4o9PL3njZvesVG3WMHszGx1jV
ebPM3vbHtx4wUKoSgRq0pTs7htKwNV09r10/cHR7yHJItEhuoJq+d0jK/VNQudpoiVO/dzsEHyKS
KHnbb4JNIy0BmDb1UC3qm08nmX6+JLQ3T2ipireHfR78h5fTUAq0y22iSnRElq0AeS899aWomB/K
6WhIlLFCONV43/FNtDyRClhwA0wN0atoMkLl8fniRRvDu3oXmMDu2+RS6uzXiy9NIny50QoeLV47
hr/HVjbT6M4TUNMndrp9B1mRMdlVGushRpNyNhGjx2jionh6odaN1E2Z9Tpi57vJ6WWq5BOLduAu
hlKoFhr+OxMOPzcB01fk4IWvQrXxu044ozJPcUxNrjJfSbGC9NDEZaNwrAGaFxgi62f0A6mM4Awz
8SzkP+HFv08eT6oD3dPZWqYNOrVJ2oO8nMGPPYgKnd6b7QYhbqO92DhkR+g5YpNTFfBzKFeRSaTG
q8NOXpfir0QgyoTucNhHHXVsd4SUKaIU4trp0KpGU4vKUndMC1nCa+vTeHOXd3EaJp0NLnAekWhu
xZf5OSF4ygvDxwIJloyMPstaQXEPehd5V8BNmJp0igFTsplJ//6KTcZ8PGg2R/uGV9HN942EhKHI
mOyjap5FIVf8jGgVMBqGYMjqdMSN+jc+yuklVU+GYrzhT9PbhTW2NaUi8XFvktHNL6kw5zy4Vyf8
lcyxw217m/1/8QuEaCc5BCDDBRmVjZi+7tMRFhyuXDAWve7LhDX6hr9SRuJ5Lf5czpWWcCsE5oD4
KmeD5nEwZUIpq7LOq3uLp2+IK3BfEKfxuHgfUwjuFcvlkBtr2fXjUebccTiOFfl8qrLZ5v6WyI7+
Lfx/J6xkiCXjHz7xKFedDC+ASKfFzo2Xj+GRtLkjsAVmI8LTRwFqBzpJF1EXXSYfXxi+IHxtHDms
o5VYCH1rzeaQGfKiCipZ3eBNuHQtQu5IAbBsDaX+aRmaw3xcXT9g7j4RB35UhzAQXfYhtL784aYe
rXc6br7CVYSFlpfvS+9/pYJwpuOUxvNGBICdJiP5rAzvOKVkm3vv3mR2WbeKh9nvqWC4BY5P7cLR
q1arnXdO6moO6QNUKD7RlyhzqKt1Ckl9faVzzAcjbNM5UWrk6ST6MFT/yXYi5O6rMo077lBWYPfd
6gC2lTouGcBOVbXmHZ3diNR+ozcIucI2T8MAU2h38Neyb1gtjKaBOFHGSPczsBlO9TNNAcq1Gg2a
0lZKf7dSQiwfVSMX7WOZ2FBNAfLvsXGaTjwgwxGS88hpU0TMOfB9PPDx+KWSIsERApX+7s5J9UqH
VeovXw13ZsPUmf9RCq/fcD3xc/BBGbBUZ0SN74IhHD07G1UzubAgidAqyhSPPjHp8hneYmv+7Bnp
gtkdaX4AGHrN1cd77nDbxT/W92Gy3/HtEjYD3X3CR/59WExvDEHsDzcy3aksVeWIan7uXDuFAwx5
/VP5MwDK08xIqiQOCMpKCXckzGyI7BAIf9TkQVbPjjapugjuggeWFKqDFakhmWoHp3dIBvb+CSML
5B1YRjNAFIFlDXExEp4DlY17H10uvvdTDRpOEqd8zk8oTAfu+7m32arU7Z8pQocwHhhn8LWOqlL6
Pz27zMMOxeZvTUsSmwEPnhp6rrnD5Mp8Xad6zGjL9f+L/6D8/upkfZBk6ivSj1s2Es2rdHuKrl5K
V++g+YCg6fD1xh5C7G8D8TZXEIFgz6C9KGgCpG8tbQcrCE3MoOcefmkQltQ7NGg8NcR1+KQVZeZM
kYTtSuJPSYAavvC2rIYKRwqx0sZf3YI3zT7TUcG2BrM0gFJcmNFwr+pi/JlL2W9Ytana9BoNO3Bd
W8breEaSFHP9OVfDHHC1gRJqfIQbUoG0+yztFTyQf62YGDsd3G2x2h14plpowGpAAfZHK4XrdJbF
aC33tNgCUYrvNHUEkh8es1WFNMLznfpPl2RTlGi4cKV0ACTbdfLnaEbRJD8hap2Mavq/H6UxUu9i
KOYy3787oW9KLZEl37F/psq3TjTYxraEyWhjA3ExDa50ElHZ9UBo7zRMAATeGWsoLg/qg2TxLK4H
5403HVd1w/BaXN0W3f50DVzW4jISvBwx/DcuqpNS1XO9yQBQGmWnNX7X7lBFI7wQxwl6MMrMXUWZ
uaEMdk/PrV/uHbSLiP5fF5UN/wV+mKZ+aLX+UISoUdiwr69X+xdlaixe9SxdZXPTU2gb41h143OE
BsA3xxaUybu5tSNOX2n5QheBEi0bnDkNgKdvlbaOewsvyRV5qBho7u5R9Ex5/nnRODbDHnJtgnE+
FKQhrQof5n+7ozKaZOcH91R71bw8T38y0k7zP0q4KYy5AAqIkKpmArPiF73JNEt0CE3Jbn/3WVCS
mbyu2dYa2euPZEzUjE8yhJ19S15iG0rnEhVtv7E4Dpf+Efkg54KE0jHpFDXYE/N+/IMAe4JAAfOH
w+SCSO31dQMRCNv6QJ2+ZKBO3179AVWvYty3ooW+zOR8GDkcrWXjLAAonpNhFfajDpFBGtH5S4E3
adrq2o1K/+lezaI9wtDqIs9aJALp8z0UDKMosDQTufLECcA42NvVpKch/5QXOLO750jGE2mEaXI9
Yxb8ZYbCIAA5h7dPY2bYpA37hE6aT9nWHfLsFpPAemW77/a13vf4uVGj14qQ/aq+Trd+4Ptn3ojF
Da/xNTQKMtIces49C4Zryt2QSAOqNQEiDFqjKTqGiU83Sb0CtHWPi+LLjAWwMIQWX6lQ6yDfGsqg
tdAvcg2Vt8ZaoP6tJp6L/UjK+XHELt3jN2q5ZMkLhX44ERn0WRdDJT59ny57rg51uPVWQLZdjQ0H
TY8xyzVq6+4rDStdPIDzIE79loc/dQlzSYZic0d7tWtIl6AKlLn9LT/ksNEy7mlwMUZe/JR9kfx8
J+ToLTy2BEE0lXfky5DwBQjZn+arbw+020RUxwN1Z6bo9pSwkwwTAbTiAJ1n1JDaHEqQjeZFinD1
RXVZArqmDQGh9SueHW6oyTqTs6eUPhmqIrrPpOp/VK1STdQbfo+rM/FfpHi2i/hQO/Vwd9+6ga/c
10ViWHRIt6VfKdk+M7v/SC1Rr2OA7MthI11zwIHJGomKLucsHB66Tght4ywyDnp0YWIbuHr0cC2S
DQl1STZ80wgu+xN9Qq25+m4/4dj5fUihM1S/8HNTKhnUYLCyvsjIeLvg0bGJI971rtxUgB2CXlAF
cZ7qbie0Wz1ugDwLfcO9EnHxGftz2n3iN/fAA27s01Br1eHPNSALMnlP301oAEynXc8gdDriOB3D
9fNUIBiGZUp1ABcEFfnmDjZnMk0s8O9IQ8pPJPpSxbEZKBf7JUEEn2xoArE4NAymsAICk/r1nBQ6
85R3548fvYs3GQ2k+2j5ZYOvT7BdaoGzaVFiIwjcKBnTUFVdi3jCB2ttJXD4emDbmqxUGi9lzZGI
MJ9t93UOU+PdifY8ot1hD9nr1Mn1asTh49/2Vpd6JVBwdhygZUXvGWtOsf7TVzF1xSUC8sbd4cgX
JR7NQCQYMo3iIyMsB/DxD52wf6Spjj0rKfBwmomnKguxYYOZWSbYO/BO5Pw7G342fL3FnvuxKTcc
JFPBvmfi6kya+pD19lmTGB7aanwEll/8bgzmD70RwPTjswzRznmIXK46lfr4Tt/5YZk/KHD+1UA8
OH+vHbOUG7lg+EpxmKjwhJvYItpC/6a46vQv81mTWYoc3qqehi6JBMA58LuDg5QK7ny2jpxc9v7i
608RgaLKOLh7Sn+GncPN56Ec2ELtxodqoUfuzvkLJYu0yuORRD7ugUWrpxUxlrsYvxUJQ5Bpa1YD
YbTRXYNbJQ6r7AFjutSsBFfrjKKmGaq2pwGDQ56mZkl7wNsxifkHgPyYaTyfmd3Bm0QLpTOqp2vv
OLuDa7EkDPoi5KnDi0K9MbDGPrSFAoD25J+BHLRKAzgbUL1KuO9VeKRV40SPzpgG4si3apPC4OWC
UNx86kkP9DqiGuACfLTwA6Cm6LZ/NiHN1rpTfTI3IPx6OAT7jf4usvVOiv2KRxJTvGvFvzRLMj04
NXhchnCZPa4FB4PaARL1bhQgZ6eDxcqgn9GF4oJIb1sNiUU5NyJlK9FtGnpxGROhssEgTK6jt7R+
vKs2xfH83uqzD5PnuLYLF/7YyGZtvqi9Idrh4e4rysAz7uyvaW3Gi7iiJLVUtxRTwDS/56qGAiPp
IlB2ywl3oB6wUTrXdJJlw/P8/fen1zkJzumqE5jG/XoJBIH4hH5wxoLXnqulWiIFcghobiiDLVN8
WaTlMHTpempyx3o9EJ0yFrM9j4Lv/55L2vAnTlZvu+xD5LPP668+2X9FMENBOz4c4d3TtGk02xSc
392afGnbykQ05UFh7VrfX0rZWOdswpNK8zRrGpsD0rgcio+yAUxs1OP3bHHjzU1AoNAQYOLH4qlI
j7uZccISgeB+D67xY8UWxX1xBjPTDoXVFMYpQYk7PwW6rqBulSDDEA/WEu6clmAg7iP2VzSdN3xC
GOscdOz0KEEZ/xTtLZCT1P+dRyb0jv05uhwzhubPYfXEv5893m3vv2jo1Bv5/Sx0WFQl/x/ec4Jw
OB5YIIQAGD5iFTLKCGaC7+6kEfe8JmWBdTNSAW7XbI1hWy7wt0BnynAa4Q874wjjYpQuEXFzdv03
+ZBL3BXitUkehxehcsnJcZQnB2e5xi6LYDMwylMa0a3cAf5ZrG62HiyUCUHmq45UO7Y8bkCEkVOG
ayCJ3zpwArpo4pvHS3Jy4RCZPAgyjJeAPEJ4TxvXg88h3YWqWkNxzynyF/DTflf7Bkd/N1RnW/8s
H7hlGn3fheMiDpvGwlRFUOi63PomNiJakhGIvKOghjbomzM9PlocaipYIZzqXyy+5eJIOP7hggR1
CaTKyyyPeLT3n9lFQiw23qmklm/3GbHLdZd4OaybkvbgX4W2h+DwxH1sc8n55vilZ8m0kewkONeu
aXNWn1iFIz4nmYDCQs8sh4qfL4+SzuABvW+srgvTDPBO/yiGJveUihPyYYjs2SqsKe9s9hEgzCZU
JKURafa3jetUOdJvbXMCUz88wZhSV64YMswf/fqDa4/dsSA1BLqZJeqPvxsnQH68HDOV0zSolMMx
xXJwTDTSw86Ou1SJjhnW3Xf3gn70ivMzkA/n38fD4rBsHRU7OPWlj7h0EI3clTpMaeqipUUWQ5zG
5k/jT6OQ35QAW+35NCixMft9kgZ2AmEtptz1AywGiCQfG93Th6xy5qL7IMnx02dq6XBSbQDuUV6j
77bclDy0rXEjCyf76C7Q9xQc0vQzfOcnMRDoERnB9gMWJwlE2TQMNlCFVfkSGSjcsj2TPVYDVk1x
RRXPRaDIMT9olP9yXKkMszWGalPVw44wUnou9HCCrYJYKZ7WgQWidKCNBiafLbun+Ohe9XZsxrUx
hPvik7XYtVpHEt0xEu9AlW+l7jKBA0xl5hUBpU6MK5jWSjln1YKuSbkynrMRXDY1HjeOs9OHc3vs
/eAn0n6biJlHctwOcvEH1GXTtU0r2AZ7DtwaIg9IYb65GTgOdGit6Lpp8FtAroyOhpNhN3sfC+YW
vRIrmPvpv0PrhMmNtaTJ6UyhOHnElBjNMJEFV0R7fYPTCriuMbPxKX2RIiOeURRPmIM/pNM52/cM
X4TFCicjC44HGAk6B2pP22W5nR1CV0qC3rmvDT5hITi2Hotw79aVN5lNSdvusGaq5B7U8t/ZK7zS
eNsxmQxxqJE6iSjbrkExOxrjesUBs/fsFAVls0vTk4Kq31DVu0T+ERDyiMWjZ/A1J9M8QPGH5dWG
lh1zgwQP4YEBbDidcF7tbukPhq6CRtM1LP3n1U0qhfreO6qgz2Q5lToq73REROKpzNycnhxHnp9f
WIAHY1G06QGbo09YCHzwT1t4nTGNLDLjktfDrGRvChjYHhS5pkR1VN4JmNfTWsBa401Nxkc7rEUz
ZKiqNz0ahMsmiZmGAXdU95uCeVZ/YnYo1CBgPd8dnMLs27p/4UWMu0g7pE/c3KROXUBRcZk4RcRA
yBSf6zeYLIGUbfpAXNvIBijkYd0D/ls2BP86BdwskpHcD+m3tKLpWtGsoKIV/0LIblo56lOFooPO
XddLenUoXLUjshnC+lu0TcrPRI3plcUSU9PPluda0XSJLpr4kDBkczm203k2PT8bmuoqoaqGxRWb
hO5FkqTR2ztNosGjhDN4D/2AD0yrdWi4m/WrPI79zmiqPWqdAtw52rqNUGRNUsmKs2/LetF1kHfL
0N7hJK2CiBggvw95pVV1Ye9aCXKH6yy0ULyVlgVNamzobM6DDQg2AsRfZU61LsufK63+UAdnCyvx
A1rhaCovAupT/9w5gDapv2eRpSKTezHmtqxRi8lTju0Rv7K02LC5wDYDLAHLjumeu3D8oitr+mhf
UXJxvB4A/I5RB236Qlr1twDg/ILsnae68yHS46arEf0iE9NL2E+LC0IFxC1tvTqSQMvocSJG0EXc
clfQ3UfSeUWtjJjTg4aI1EhA9CAhtzi5Fb3dnVsGVKxu9GQVKxXlo0sEipqErmxJ994GX2zzbV1g
1BdNKVkp+UtUFr73kklJ2HKdgURMRb2iw8KpuLnTKhNZIjpsJU/zrzRt4USTQQlwwD6QxdF6MVp5
ynTP+DhDeA/PUEXGv3sP78EUDXC7yHM2CozzJFgD2zikjKqIZTUu9wEHEfwzS2KdNtaY+CdHCTo9
MLdgCEeXbo+efGSXgH4vpASaWvza74p9ugw/7C4FhHwTVBmw2Q1Cgcski8ZxSFQxvH8nO0XaA9M9
IdJ9HbKCw284eIGIO3SWsC+O4KSv9ohd65ImJBl0Rxk0GB9gAWYwhqbnu8pPvbtUO8096cpi5FKc
zMsLytzrpo84KBovJ0mXgm/CCBrtcvtNrBOH8PJG3ip34oME7zWft/3im1jiPOEd3Xryzf+eBFFA
BcZBS15fxW+kjtYRooBt7iiz05//ieC9SK8nbSxMy4PmshUyPMQOL0MkFNe7QS6agyYJU/cB6P08
eSISDMtzzLcQ7Sd/IcSZJy7fzJnCXT6VK6KteE6hQjFpMuls98rRy7ytV3P1tvyzuzbcjqQfHKIH
WKe2FqfnbYjVrM/NvGCD6Erq/Y4CPt3kFBOC1hzFvw4DUDGfSMIHpxzrhOx2edcD9fEheepGi4Sb
JNw1mKVk8J26BT8wRrggEhzRB+t21Zqj2RkKVdfjbka5IKgTt6UUmZN4y+b0JRSYMovY6kui17iw
XN+ZAj5HegUy89UaYgJX/sieY/avgSQ8xTeyYvg+naa67fwT8E9aZb05AsxYNto8FrYPhYmYMsMR
/Y5vKA5oh/gc1TboiggtBBya4i043JQ6bUcQ3IBLUM6v0ZAsKndk4kqLwB5COMsqK2S7NzfWTwe0
ZzorcyODi/F+desJ9kgkknUdGtjD0sHnGchQMJ6Bg4mZU1D5lVElIw8v5E58uar5JvGU8IOvPdbG
YM/V1uDEI58aC/OC6CBHZ3QKEW0IMpV0mqIhGhWL3g26sfJ9dDK7KvD5zF8+a70RJ6eOl+4JHdO/
29ZHYcwUIDNF8hSwrFdBbBpMxVkXKg5b5t8UP7Po7BiUVLJLesp6eBgeSYiwgUWIzB50Qay6OApk
l4/ywTbxmY3MehY2XjXFUA3VV4Cw0ntGN9iGUmIQLYqbnDE7FkZAOifT0vaxezoNqEoMpeaxMwT5
71fDKXGhHKQlXwGdexnIamuEpxbkWO6ZVvBPt8mf8MJjQU7Kab61tl6HyrSY+swcLbGDZNbX0o5S
ZDeqJHIXMW8M1j4OWr9v7qiFcUHEaiMhLQPYytXuRM6MFqj3yubKyGMAUhoFBjpDoav3K8cU7KYD
dzIUVrj43bMIsj1l3oEihOcka1aScOJtlzxEqpUjsB727KHsxZjqsXWxHaSpAxZhnE38ejRZFpsL
8DOLr5GTy8NARgbiw9DQqJhws41hJs/yPVV+H5r7oBwt+/Lmnv2nazb7VhkHzUO2DCaZCp1OLY95
/I4QnlD/UUAK2Ndj5SuQjtI6+7xwoczuPwkxLA8qIRZ9mh6SMHIxvj1VH51CtTEUZ4OVZJqjQn5U
8dOyUuLUrgf330GUKydUJi8AFF3V6cG/pgvLuX1cXshCLmiwIiNVUrWBV5BZ9DtKv+dLRuQgGySq
AEsZBnUrWlC+T07S7UQkPW6HpWtTJjDY+Zw3kxu1FQfedxWi9XGtQcQtmBYDd/QzH79NEBdtu/bR
cvroUrNhaHm7+L8ApSeeAvrxchyHfa9ueRW8M/MxcrUwYtyEv0ulXgW2ivCP2URGd4tcXClWKPsI
QOeduaxTtMobpTSRmO9aAkTuKIGTY0cLxtxSqV8bDAXV8gFGFRK6s60GsS8apS7bsE66ECbwVcc+
EYE3keRTEK4SKR1sxOyxmtVbAp0Vvr4Ncn/c/2TxhUbjRtF2vdnmk+rgPTFCIZU89Ptuld2bsiVk
CTN14CsHomhtXMRN8+Bs+gErQ0A6ZQ/1sM0dU35NeQGnAPDfDJ9xOlICepbdVYTtckfEJ0L51rm8
Qkf+O62DvavIDa2TRc5eruavqa59HxysRDxpRbVzWR2Ih6OHkNpI9om97aQt2CkSFgMBeRS81zNN
GQvtHkQsDG3y1oxPTB0dN5GlUWcn90NKKOTl3IEJXDquWKoTZEqDtGc4KWGxGR4Mt6JUKa0iuWDP
XYU4RGZtul6XT23TsUdd6/F+tInAlyzg9d7OSI+9X0Oqe4ACwHi41411aVuV83bG7vNUXbqx/MuN
+hC/G4fJcEudG+2z1XpfJlksCbO9ysmfBMtLL1/cvKIC4Eiua4kFbZgXhKMJmp7Lgqa+FmrNbKiw
MOLuDpiOeElmgEGckJuWCrlhhbTasxsvd4GG7+II8/JOWg8yNBtmuDmaN/l4kF0/HpqV2v7QOOr/
uwopJ36+htlIE40weKGBhHjAzUYqOdnb7xqxhDtC627f0zSa/n1f5X9r+9z3JeANmPF7y6c7tIti
HnlINfji3ty+iN7BjrVYYzjo5rI6ROlBZbxhF0QhPvuJtUED4pAfG982fMPLuW2se+878yw3vw6I
d0mK/Npz14W/sP/hCKvQWc4bszN9XpCZ5QVXQQ7faU4chqXjkp2lzoxHKzbq+E9eeI9fiafHh9XK
LbJSZj6F+uPaIsEW/b1Ke051W5CgTEJ7bRO3J15PTymg6bx7SlhtpWGRE+84PRnFWewXyhUOcD1q
C2ynmP5po/X+yRTymKhQTZAM3kaMt2Kg1Fxcg3WTnjLG05+KatrwhE3zh/dvyAfEj5NZncpPoS9o
+8pWF/DB+BsX6xBgOowAW5bZRmZtPAvvEfRsldfsx+BiQGgOC6PnnYEhC/dA/jdW+fdoNGM5+va2
vzZSyvUrW9iRbvh3mz2T6Twmo9dHXywe5QE4jFc/ILIQ7F8oTuaXgUYW0HDtXqemhTsGNA5FOd1M
4WKjfNKz626Ko+7de77iZyUKhtkbgSyopEupE0UDm7xKM+KNlCEx4B2T3jH+CPZUUdb1M6oSUhkH
vMe2t0s3ZQLtwgbH7Po/shFvyyM+CduOx81X8kCLhkPxpDEtYqWyI0M3/wv/vAgFwq6GJ5lIoRRD
FxcYqwO9GMoKtj8DgrWh5gi0jWL+jPVrMrC+n7zzJSnMBR1FuR8QZrsoSh8SjW8nj/rl2YZAyrxD
+oTGK8Asad4OMxN7CQC6FZ+r4mtU3EfzxEfRbhN+3YqgJhHD2/3Wo6Edct15kYeQFSi7QBCHikmO
/3Mn5D9EN14OavvGNeZ0C02wkTpn1CzdK51VwL/kYmTjekxWlHZZwb7QJ1Mwt3u7amUVAaUo2R6G
n+IXk4xz0lvtdeZ317tG6nBSvg4klwZTs0wiLNfMJzGkIRsa8Dd9wvk/irY86ojT0EtOAa6TEFSd
EdASk78p3CGTC9kFIkabSEz+4qJvNd7v1ASqll408eSGWM2eJfFHutZYBEEYQoUsxBtNBq/unXGZ
6zsEmfy18mYVzPtuj42MWyjUNGUTeU0N8AqIZSiY1dM+/lHjDKw007JwVQ+lG1U3aDeqxUcO4I65
LYHOsc3cC53SAMoXgeSk5sz7dpwwxmrAaAnsuAy5sA89vO+aiQqAZjnQdK0KCSrT+Ow216zDtnCo
1siMIr4Fek4Lif8/s0yeGGz7g8mIGNoSH9lqFwoaJv5VGAe/6WlHs+zk5GGdRyRkFK9TTim7HgBD
Cc97ifg7xKHyYCr0ibnk7YGM+Ht6kj0PkDjQcy9YDOk4Q52nGjvoJR4SaFIR2YHW6ZM5gSSe+xt4
DpoZRVRlUcAbNOFRGbEMp91pnoPcyr/zQpcTtDxMsb/j5QTtbGvlfjIB2QZ/mFOj8rkKz5UN6r9F
KPGyFkLSt4lrwHWNlEtU4at+bPED30ZeW/AaLmsu9VXefGfmkF4DG3zWNRDL08+ybaU1gstdU1M7
sFHJwDIgH3HkmWc4McE6iPpLyeAAqVXzl9xtSLtF/L7HSQlDtCoEi0Z12VxSJK/m8P1znwRTvbFv
1HOxeguWcMWC7xyy0vzNMQQ6vzHzyJHbY06OuiopH0/3w0zxtrfriNvqvrklACWgcbwwNjlUbpC8
i1nUlDJV9SltqHIAZfK3zhatnv8SFSZQHZ3/WMA75xHEffrfMYEQxMLjeSoZ9il6RuCfob2JWOhb
eXXpxe87AgfUfKsl+b2QwKm9Ml2/PVFpRxscbb3mXUMjRTlD1F1jsI/U32kgl0zfeo7X+zDIQDB0
zHtEaaHzO+aQdDliXuB/NV5mkn6D8KOxsN4fgUN77y2TYj83CF8gJUOPktP+GGBHocL0T69O6hHW
Fcxcjcy/RA6t7slH63H8PRWr1aIRcbNdiJqPKaOETkqx5AxRF+nyJjYaGji5POHNwliS6XfLpPCK
FzDVz0b2BsqDbpCWtcAciUvKcD/eRhFMsJElnL5B+0CbWMNDhxdQ0T8BxewLhwQsPP3Nu7q7Q8Kv
MAjRMote7n9hzV9UQMlwCa2f4oW3IzW5+MTIbsB1tUA36uz3pjQ+1Qop4UVWk63JympdnEyHhnYT
4Zpkp+NL1qVqsU4isKIMINYXAka9Bf28WoXUimxbvFE7XaVDumxlMzgETR81AH+XqrY+XOsZfn0y
tVcsbVU6yPLKVh2iO37T0eeSby7N071P3PArC+3zXQngU0gOA4bOSS0UJ1m6q/FByInoNBgvhzLe
AcM31erYYshz7c6qQR4biKV3Od1LfTKWkM2X1NIVg6a6m09QTUdlvNZ+yCFltgzA5e1MVagCGt+m
B5HsThoGH9dJRzawE2O14L7OwUe39QSYeFDYmXYwe/dNLShulXv7tohnzsYECTXwpMUXmfvsfFxS
G8dVljvNQdJsiEHA8sXRwArI/5twoM42686uUXrKy5S4lzqR5sJPwuQCu+is3O4pA5TjhqsOCqCk
3Z0XZqPEVa/+WMWeP6G4EWSBvYHt7cukoUSu982oY2PCml9paahNUQkyRwqaSPRW+9zUe5G7U1f6
wgTz5jK9rPI5s/J2y+FZ9wMcZt5W08hLcPzH6LoykQV9vcGYgBRBEGqQcjx9U0DL6xE2Cy7kO6KQ
9lPy/iHjott00SsBqdplPwcYzmPzZxFzBrbdahx7h5WB8bSF8jQam/VfN43rehbhbHasAGU7oI4D
zeUCelUZg/yWP8rEvvZk1MV4vp9aqyEIa1+2zXJDxtmFl06q+poOQ14elgR+4uS9PT8r7ZSa0L8+
R3uYYb5sx4C0yqwip5B1PREMr03Qq2lKGlXWo01bEzIxWX9ySLdgLgcqb/Ur7tqxDSRmVDcvy16V
uTQRsDX12AI72/sEtMOmQV65IDeovjeKt4ztW9vl9n2bLy8s4MzoJIA0AHxlf0I6LXQwMX4GWFPk
7G/RlGGaY6V9P3QQEqBMLF3h8t0X9/+mEa6Z9+zTucUwvL7J/a0Jg11pAIyS/FKPPgttrtaBEVrC
gQFkb/21lVHdQthjzHsl7/GwyQYJ4yr8bFY/W6qigdVQUI0GCr9krtxkGdpR48nh2T4LODRxFKAa
WlSQRdRKLT/Y71oeEg5oM/mQHxWxqquhRwWhloupGqcP/2s7Z4Eve5aTQ6tH4RdJGuOiRlYny5kD
nb3HdU4GSk5A8+twTIk3UnY6x+K3Um8q0sGxhAZUx6z19Y9k7WNycfw2V5PorhKWSTvtxaMN9UQD
voeqvvFef3+jqKNo9qS5DtUgiFp+9KShljMuvOiLYthgAuwaz9pGf41IKsfZwRJGpLCe6wndbfPZ
Fg6v8gYbIk9PbWAgVqlLFsgKL/uEZdbRWcciMVr5I1x9+6x/sTH2hRUpvwjIKgTNkM5EteaPd8pE
WYeck6/eFBFjw78dayvDYQ1HVX/y65p4vJtQse3yv/GqrJuBPjfzgA2cy4eQZ9oVIcqG1qVRVXPR
ZhO+b4yMJEkx9JHGOOrSlT2A2SaWf4TAGE79FHXOq5BjNvvsp6RyygSNqy2aRUP0oJLjHYHWXoZm
EpJG0LeUd8KGt+yjtrnu/F2s7WoN4R5pTOOes5YdlqhxQjK/2FhqBD0Kcs9aZN60PLsHTHJhtCY2
QjWCXY8loQwx6Q97VQ31ovncFK/GHN8XDtfo8+Z2lX4nv5MMtH82N3R4oPT70XFvHOMG+TqAFSKx
L9Zqe01x+fJxxcPCjWYmnSdoRR03+9G6A9nE98U9gX+uI0OITVkNbkUYS4UArLhW4RUWbnHdRuCi
UgbCvJ0NSQhtna21Jw18qFVqyRt4vIITCq7le5HI0NaHfUiDC5eZ6yfXJkBM6i8+AftXI1HEJjwz
UzE+0SeI4idsiHK2Hu0jkifChmGXfV0LjOkJsReFGcAb5Cy/JE0TgyC4JxzxCgfK/Hotr0anaemZ
tBT3JwJdmdNxKXfv+3mp6zw5qzkfm79P21wBljwuMHwf59ikWIPvW6jlLzuaWCrbn3pjeoA0vV2d
EE5ERmbaE8Qd+adauMfM3Ym1tIOk/lWCFSPlol0MFAYUfPulxbcohcWMu3ptsQtEjYL2Cu/c6RJr
NtI8EgEmBFX41p9akBv+tDR1a8d6KW6CA/8xn59GrJ3zRTyHAlN7AK4ev0RlfOJvRR6y7FGZ0fiS
MiWZvN+GQ71K43xvd6ehyjEi06dJq8L0ibXazfFfGvLmXX6iMd8Fzs65b9sNoGBlw5O5Uw5FlfEf
AkFuzm8Qq2+VmSRq3Do4Nqe92YAl07yxusFhPbpirDBVSrmli/03N3EK5a/vWbmeDu3vrMTDTX6i
QdmebX/E2a6eG+PYybBorFROcPZa+DC9ugaCQxljDK5Z4AXwjqTrgVTKz1J641sNh3OxXNPth8ST
keItXXgAoWtnSzmqCndpg+7SIFTomQkcvU5tBEWC9/1JQ9JIikUCDzE8louAnlMspiX+zYPp3TRy
rjz8toPcvy6v+FC7R1If9C2PfuBzQpOea+MMeKH3+iMmidPhYeRzkvGsqcuiXjvs4vUkWlrtjPaU
92a8EBK4kc3JqZEuPMECyhbm/UxuylWuhRwOC2AhJliupNvHQhloCUK2D+7VU17L0ZemZtC8tG35
yUceTLJhB0a1I6HZvnsUrcRePZWd+ZlAAte2GSOI4H6hdMN2kxRRHAlAUQ00C/A9HWK5WFADCiJ5
7nqq/nDK+0REaX+WkknZnZwDEAZ6DKvA41BCde5bucE9YDi0lgnH0k5dH9enNOCyoSTULUz7jXSA
IPc0FrXUSM/JvQNLzSeevaYbDQtAFUTkgCUvmuQ2vFCNGHB/cUx8jYXY90Iwma0KAPODSJpgF/Tv
2GW8HLzsuhxyImYbrMv4prbnpDgKtlyUc8ThmtqjvO7UxjBkk9bKFoCyutXYAswIP72Go/IHjApq
SBLZZMNYkc2kAFI4xXc3WC5wQ9HpPKJ4M40N9My0VVsvOegERq+a5V18APBui/UuWr0I4X4V0w2/
j+sQ/wyoChC2kvqukdYrBSNDMNBHkI6QDYBPAX+Mt5GGye4zSg7C7jmUCXldpNO94yPpoyi56UQv
uPFAnqD8H5lV7HVdXpjHgWSGwgeR2qOsdCnBsGwwm7swX12vqwelN07c4uJObpz+6VJbi4jyTuhC
GzjsALPx0yDCX4OElRTx14dTnvhBdM0AEFedqiqw7wzTcF/0R8ksnp5a8tNRLPiK+WhvlFr0e1oj
MVbSyuc0NNBwoGsgzTE1yVqO2VkkfcVkEqhNbA4bgoJmrzEiU7JgJjuMQgTuoSmkqbfCS7cERudP
Podu/TmrvG4VF4PZF2fKRRW4Ol2giM1KFZmoSBx7SYTkQXOTbxoABrT2JapxjNGZ9GSPCjAZl0/B
97ktWEeO/v6DZygK2iZn/nJa1ni2+XqvmWOjk3jU0YCg9aObloEPBTE4Y2b+h66GjMkJW5cPiKCr
XedZxwadqaDXMu2A148OB9vTc5iKSmP+rBKulCjxPBRBP7GDgvU3EeIKUCXbaOr1a9h+nWGADRY9
aIiwUwIl7sgzbsMABfxsrmueUQknCAfIa3hP4kXGtEeleackxBocQO0a9A+dXzAFXPZI2csFFm0N
bwYFVzK7genQfxBDRtswpr+NrIltILBWcOOhyID8syezpOkkrHYoXXYiPZ/teX9QMmi9RdfQeN+w
52E3rtetekcKJi6VVlb5tardCjF6h1nhuVuWlnNc8PSYtXqZQxAqbX5sHwQ2LHN3FmgEu4iIiidn
2/0e/fUC45F2fMFiSO9YSgfCGQHLUUBLI9dZ5TwpDgQ0SFUsLpAHDDJycP+BW7pl5yZkU4dGGqRp
hnIcTBiIxxjGKk97Q4J4UrX2Ckc88qWoDW+AADX3DlJzP0i/WE3/pE5h44DTFinTfMECLgf34FVL
vHIdc17BOyvfKeeid1fNVN0K+L8w2eLcVr7/G6gILI02sUh9H3vwT+rQj8wDD725amttisb0y4GY
wpKEav4sUtpyov1/HfAkhvxfcQzMzDLnLVol5vCEymfjAWl9aTEZVIKUjRu0ID4+i/yz8d56DNrN
IinlFJNENG6Rj/QP/+hmcIUqYi9PaSViTF+jkzR1k0poNOt9/M6Z6S4T/XzaECjrXApO4WEEy4CB
MOJ5Ci8nNHmvYBlQymz+wKegIlsttu7QtOV41s/wlLFhmLONC0ki82qh/8yIHRPrxLOSDWhnVyHL
5S2cnU46G2YjEyC4KZTfCkFZgLBDS6C3yHN3pgQjnBw/3RT01t8dQhN6hrPfTxhz26/aROz4o8ze
Cl5aqYk9qYHT+nthYEvWZbhRjdG8euv1/wgZGKa6t+gegUHYr0wwRWxT2tTp7lEsOPVQBEOI/4Qb
AhbYBK3G4aWP4LJoD3q3LD5Hf8AuzPgdIH7iylkLwqvnMKRd8ix77rSyUBwf2RTt6NzDxo6Jt2qC
eeifnqK6H93dJe29NYvs3JjBzP2Z8mkbJcWXmrqkPCysO1L+SwpAojDJg1jJS7qm8B381jAAqAlp
cMYQaZ19dAOEHrotEeO7K2q2ri4jWjGd4OI8opCD3C3sJMT2Oqp0TBmZtCYkQ6J0djb+9fKtTLrq
ilQv679hr0e/K70YV238YduT2coqmLVX6alHkCnBYwYzg0IGIsSZuZVIxTNTKWtat9YO9I3cAuzY
YhWDR6cc54j77byoqGXHI7L1Y85cDxG6qlSiHeBMFrnyn8yHXNXaNbnOhrhlIwtT7anYwXQNFQQK
3YPgDj3XBdUEcrpJapHoxRiZVpmissXAnWpIz1u6Daqq9IDDjLNHdW0V7YeYaeyuPJbhPAtE7dho
/qEPm7HeA8/yoBP64w9kys03KyqCU8k0KOcYrT0fuIfVjmVG1NQAUMRGs7Jkbb1Y4jZV+BkNEUjd
VptDMgzTwOGWix+2+hbQmL3hQm1A//Rbds9LbZ7qIdJ34maByDdB15Wph8jJE6qchi1dBKX9RYiz
t5wXtEDM6FQM8D2CHUL/yeZzxINpejlobc3cZkRMilUpooH46kYnGNaE32E4WQ96gYdefz8wBiAm
1qmqHm/OUryMVqATytRLIpKQQkFkAc8PEAgDR4T4iAIcRl9Eqc0CwHnnUlEtQ1FGVm1LlhGsT8vp
T7zM7NY/0Jiy3Eq80hEHA4HseoCJ0b6Gbv+SCWr2X1OBPO9vMBqb8Tl9HOV5rN/EGuV6S+xXTCOt
aD0qaEkyHbCFKZqgMIDrhmwCO+AyrvmRCV+JeaN7olaVJeroNVE84xRROByQA+eDysjyFAJ/2KmT
/Wtuv2wmuoYC2yVs7zdUthSgL+EROuLPNzPQd2qBFxYz7LgMD1xmBPJmR9W8dX18QCa0wjOywWyc
9tEaX7eQiJ+A6F4N+CV4uR/vGU+ipq+ythpVpeUP9rHAbdBooZH2nbVzqzC104ECxblnFe+XSJ0a
oHvpZIvO8rgS4vfrlq06l/94iYEJn4CHYfoQxfxF1xDnyA0p3bctN03SqyLd5xkUbRemEeddCWTz
UQyKfxxlP+EiqGoeoa8l2fWRVzlb2aVjqY8datAaClMfZCOHLLKWBuZXM0pVGSq9/2Q5bFzODS3j
aqgOXbIjwkV7byvW1C0WNcJ9tq1QfU7Glc+mn51TpYyxsx0GGllfHnoqSrN4Ry4aEwKN6Z7nQYIT
GQ3gVWrIzI0CH7eS6GYCs/9FMfgWY/Q0gqZLAtjI4crStr6Bq5f3Q9/uVEHmb7w0yrrYyyMVuLHB
Z+dfc2rhXrQK5R9V7Al8aNYyJJ8NVRDJWXyWGyePgwboF6fkAVkU0h8thhOomZdKQ7lyePmU3R5A
Gxn3ErCXw4kXOPNCV+ektVvIRE/Y7+n+7kaCHOHRirTS/CkLD+lg1yuGoogGwAozRhiZml9ugEZ0
kiUVrDzy59mn8SF5C8j3EtxE5j9k6AHMFlngGTpEOYUM0EXontnrQWzP72Ln8s5nUv49Txh2EURW
JretsAt6SS1520hqeLNWSd47nMKmhNLrEkQEYyaWvlloOmJ/7XIaCvKViWxvVetW1XNC9VJIWaks
7ZPAbSu1FCvQ25kgszJ8UiJp8tHW9gVzaR2hz47GVPzVmqJzxW4jq32qt7pCAzhyQ+LLBJIhP7Uz
7+ZJ+I96oY+pWzv2fwECyxVDdP2xKFiYWscF7hh4uF1Tvf+adlHDCc8LzVIKtz6B9+Lc1wzT7+mJ
OqqiOKitdTelXi/EXRZKwe1rcfkRqHrOWjWKO5Mt5n/fnIbPXltzLZioFRO9pXhWNYN1WbHF7vus
cuPqnFZC5v4hXLJMBqiedc1oW0fDvq0YF+bWQgo63ss/sMh4phpjiAyWF1i8Ruvb07flnnKNRfw+
jdlXdLfL4aFju0kI6lGFt4/BGi76AkDvYND5pk6y0jJpA5hDATNNiYpBHdaS7AEMvBMPkOJ9w3eR
+jtNO17Hwt+cicPrHVKJBRBIioXYg/WBMguSSNSXsckdIEUxklE7nD7JZcyRPr/BsM2PiZ8FiqbU
21N4iucPPcRdU1OQSgOFuLCYjiL0W13xv6MnuNk2xVSNDcanvfuTNctYxOhmC7f/FXwb1xvsaGgD
BMHx7E6exve2LaSunE+wX8l/eI5JrWJqGQtWYyO7iPaOh05nd8uEzON3JqexAjfBCQZsGajeo2LJ
JY2lLnr8K9a90/Abh1YFvQHoDhFOGB5gYu+7+19U0CueVeSBQgO05YTzDBmTgqtRgfze9h4zPeAP
uZey+mYJ+VggIokXebuxh2Wh2dcEzCRvQhcQzSEpOgLcr07+Q6xAoblyOCTDO/6sy3PRiTc1OYA8
xfS2lzjRdoWPseYKv5xm6avfIQQsbuChysMduswOOf3Qq0+INvfa3Mfs6L8dtQ7NI5T4aGBlUdtn
M9QG5EPS64zUjcOxWDVTS4lv9Btxx54M0zvVUlRjPRRzCRY8jc+hde2GKvWXTS21fjgawM598i2L
h5gDu0cPZWBv/sdmMluHtuhs9Gwai+g8zIKUsT6QnHITSUCRbA6bkiiLNkQBv3WFJoAksOAFBTVX
ZcAaoRSAQEjcWEtNWGE7DhlaKq7FfPZGWg5pL7QZbkSc9ZnZwa9EtHrZ2Wd/yNaJ4nwkXu23zxt4
KQnoA5L8yusqu/u7pVztCCWZ1+MilpBXs3YABe1KtOiVJOLaw2DYYf+9u1KyXJmPexsZmG7g74R2
FT29vATR41teIjJY2fdQxvGD7UXlqTYoHp6m5oXW9TiZI8AS2TE+JvwXeDogkAXMi0k8rLYCBaVg
WlU/8xku1Qvd5qaLG7pwHkty2rrIcZCChImw0+RiHOKQHDWJ5Aq+6nHuZ92v30o1mZzJozriN/Mw
wIecKx/7s+WsRxS9xi3btCPY1GSNrB0bp7fUFn+BNQ8EmK44QPN5v8bRHPAzDAIgjor2cHKOI/cN
pBBBqdLOGrnFvnyQc0H59PSymKiM0yGCn/6uuHM8Lei3pkV9/vo4La1INAEVfpL7sE511t/hDDFq
Qfs56W+LWrtEWJ38xJKxFC2PbSPsqtkXKu1MVvV7beGH/WEytPBW9KVu3B1fDTdAH7GZVL/+QSK/
FeAeo828WREOCKMj55wkom8yKIVOAIeV+SQYMshdGf8BmeBVNU46ak2XKMogg77dEtFvqaesEN4o
HcRmorsBNbwRsREzkbu56lXYaG6WEqGxOwefVXK3ICTX2mRFiYT9CpCbzY1y6xyn2es07X5u6e+A
jHe7rBGlqz7NkmYI0DMHNNJzgEl8uDa1QILScWP8GCvHiPwK4rquNQetU5gq7TTmXN5eSNLfAqlz
LW6INcmUAJ4EAB/lWomqgrU7ulg70sqSQbqDk8BLOTVSwNL3lY9NK6D0GWnfTAtspvc0E4Pkwdri
uqdRqbvVh2J5jK9sHqc3bSu/lZiOlTWCGEqRidKe1m4PUxhRENsSPOX/ui4QC6kbC1/0Araq8ayq
FC6NBaxQk4NR3MLD+X5I4kUjqoYmH5WWbaUdCvaRSigmiyoYcHOq8QYqZABSVdbjaFQaiQZHlAGR
gxom9bEm4vNhjeaenNo6zPQh/hMXXWs3saFAwEtOCOzwAPp1TWSp15AnBpxdd1Y96ZYUerI4S4vU
315TlKeRDq3YxSiadIHH+2B60cTORpRH6BuCaPB/5k7ajEr2iKZRkxiqW19uz/XmdsM7o/TLNmWK
27QgT6mfPBQP/RnbFY7mHNdgatfzLB2n0Sve9YTgj4v5QWJgTZOj69q3tmk8+Lej4ECrWr0Um5ic
C3hWyXIHsS5uM9gt5yweLEKrvV7I7ecLKYMMGqN1piqwMCByOYRZTOyCS8qQqgG3U3d2XrdzPZlM
eug+2DIr/gZoHvDQh1mH6ftZ5p0N01XuwQh897WGZALlLGLxftcA0sfr9kKcjRaANuptiy6PxnhF
As9OMINNtuQnTxpov7zckO18MAo4munrqA4HJBt3bW5MxVCkxiqz0HHV0WEbuVO4PzNHPBFQQF8W
4a5fOvlXiLb8zFt+CSzUS8RSjhqkliiutAydtqHeo0n1HEcwMmXBGwigF7PMrGp5frKKWj52NM6c
+eLEM4f8CYK9yO5Pvw7jHeOj6HbI5I0mrqlDvKr74o2thZRY0sA7Z+Rz22BT72mYo/QfdudZSyIu
jLs9N0PMyUdK+YbnjoHtJdPD7mK39Uy0JWBcgO+mU4gkoE4OojbTZFt0ysbC98FRr9AV8Ee/uUHI
aZ6K6XAkkyCBAipt7VgzTRnJ+ksvu3kWu4CmGa5Rodptd0bqToVG6eXARYsWQzZUo3TCHpf/Yfg6
ecg/ACOmRfohcbKnxnL7+H6cCaChP9Qo6zKMGHic7uNSh//im9gAYu4+vyVRySsKV4ur8s8Ma9if
XZ1yiuJ2Q4wSTzFUp7rSiLUlns5DIZ/ucrKgpyPYS1RcvL0uPGtKx5rxYBssh4o1TywIdsH6mJlD
2M/1apdmT24ysmUg0e5ziz9BK41/YHQ3PYP+SvURLEO/A0IBNXEIanYq/h5HoO64qF3+h+x49VMS
9udregW3lnHbzk2XO+u2Kbafzm3OLGKU5cVvQomFJHBP5OQd8xNRp3tKz8I4avx29o2M4G8Fyg92
XMXjzfd2jrTzQDRfH49xOhRn6bLThswLl5eKtS257EiQ+BbSD4ZHaQCRUkvgphAl6JJmRgSSZaQx
l9BX+3LTjYtkQMURoHerjfOi1Srd4NeaG2HSXhdMVWBbPzTi5gR4ahxQg2ZEJmpLRPJdQmFr9hlK
lp3k8kZMbSztWyEYo7ZSizabQzFM7GwRFjApWhoWjwwp0zTndnGwaS/h1dLrOiajf6RJ9ykBYvEr
PWJio6/TQYMgvAnSgF6AnZkZ8jbR57CLoKsVXlg55OHgeIsm50/7AaJhvzBb8F2FOkoGrqjgLnJL
riOlhQeqoKUEPc1K+s5tdWdnEV0eEAcSehqScOL4kvHs/lxkttJb37nbawsWYKNAVPA5M13IV2JX
ta6iSoT+aAQD8HSsJquX7OxihvDIgWWSb8lI97A13L5DR9H0/4TecOPOaBsCbxANijjDxEaXE8vH
jkoijC4OrGCtjPHlGMw6qng31vEQCUf56uCooE7tAGGmGFzG2xA5P9s4rtWrO6Yqy3qZh6xqTNMs
XmEzVQah5M7PSiYXW8zlF+YgVbIDaslkmx/FqwdVyKcGsCv5of/1mM+YFt3Nl9OsWDrck9/Pp3G1
MGQ1mb4uSfrxH7XU9FLmRyNT0rJ0F/gUEJflAIVjyQKZhtirtmlD+U2G6ydm76t2VxxjYctamtPc
geh7lvhVDB0iehrpDxY+QStyky1z2DyszNOs07hDyHOYaZ9+HOEupU5H1KGps02qP3lUKIZ6p3pk
bvpzOMHpWHRb+cp3InuouQGVnS0k/kfyMsLarJwHraRjAwMukL/1jVOlqaAPeEgN2TY94u6hMT42
6IVmnntF7bhbSmpNXVBRm4tNWk7yjHT9tiMOwHEvQMif3zquSs0pzGiFE3aQhDI9vRhahGkgKeoT
CaCTAZ3aQijx1r+s68kExT/p725h3CcSm0lQOsBracB2lRMpldqnYZQ1t02A85+bj5OuoE9/R9q2
kCrG8KuM+0GyU/IS0o9LFTPdqghjeqSPsJcx5zGKiZw8lyTOdMfLLZZgYhbxYoxkWODvx2gFD00n
IZz+LeQoeb2JStDuSvn2GZOIB9QkQQoLzfhlwDU1TqmdQv5WGyCmia2m0gtY+pMBOOw+DbrSgXI9
XzZQArsvpePTbW9PY131tlAlI7bm9CRpZ0GGpDstR9ar3jxJhwA6NI65hofDAuVijzRLINutylgY
JwzzVqEIKBPcREY0Tx2L78+AABtaArMK+UliUhGAUrhHlzV/69svTsSIwVo5cuy+RicrRU14wNqK
RiauJ1b/sN4BfJSAdel3owm0/tgBsWm8C6AQRhmpU+sysk6SYxnofjGOU2lnTflnEZjNmhFPsXzH
qXD0h8CgeRMlkKVuJptr+jF78+HLVTfz/GsZp1B2JEZClvnVY3fu5jyL9IBE5VpLBuJCXZ6OwCHK
ZrTMkXce3obG1/G9B3mwrZ7rH81t/O5J5ZnuTePgHbVKJeqh2NjKB4KsjkoppgUkV5V70gpmR77Z
rbZaykYa/crTYAJ07FdJvuj6PbJqohcbbCWJ/1Z5U6GR+ShaBWX08DufLTqzZrDjLHUCxoyLGhty
RtZIAk8zBQloVKdiv8KhkgyAGW6EDaDmWoFQ75ljs5ULU6amlyrILs+kEBR0uXLx4FFhxTD26Y+S
Zpzohod9lgJvHvJiNe8ULbFQx52U1Y39KycdAhwNRz18s4njbrV7RTZcharR2TrpyslmJsEYQ9w8
OIop3Y106bBNZh1nEGIo3PSvVdpTE2ViztMfGvChZqEnxDPOLrm6MlTyvdOtthJQzrcgpm1cUC+m
NciquhtUGwHa6M0/PfNMcnEKLHdwWjZSH+HXYtvgdjyBvHl7HilfjIf1t/MtLnLja55Ix/1RjILx
R3yGZSGgfYhMgPeqxFHKUS3IgbmTd05kZg6ZqJMLImGSM0W4g6FkGMBaWNAZSeq7djS0s4g+hiIN
qgWroxjN7Q7Tm8Tuq/TNML2Jn6WHoX/eW3acVZQyXNhj0XwtgZ2brhkaBNQ6mUw1iMxNi72Cq5C/
yrA8fSNnO94YJAv6GXApS9aIQU7NoFrcDujA4s4OVauJ+eTjlRkOuaLdgTRxK/v8So3fa9yWMVcH
Nqv9qzybbJ3NkhVNW99EfWdU4Y9FxuBuT6/uisWiNuYHdWHFVdeZs9TnYA6lxUbgVpldq6Q+0Mnc
GoyDlsgHaRiZK/ZPw4a9O2W5YbfK2tzfPBzw1GQP+0vnolJZD0CHtBSOvGgCIB6zXREYsOGxmFt5
lAS8fUi54HuFjxV/JiEHrl+pcAnvuVZ959dsvJMluUNPdaRf5dkKtglLzdmdE1bpaxwchjfkAXLw
OBN6UW0sG7dmjB9Mu6g4+GncLe1VK9I6HkUZzxEvbKQUclaTzCoEhqHjBGu+l2+pzooRRpPLSWzS
AJNhAGpzkpEckIZVudQGIswUqk5QbiWFgg9y0TrUFaaFadSdGNYwSH1dJPv/uA+rnNVyinNh+gPU
ApW+0pg5df9Y95gOKx+cK/lmBFrKyxsh5qnZFnCvzZmXcycRwe9A5mhYQdwHVjJtNy9eYKdNcrCl
0bhyf2i4KgvItzZzixN3gv3a4fJb9n/kkQSx6H6XGhIWcJ7kD9TiAdXqM/Bx1ICK3xoYJ5pb/0nd
pTaICSmrRd19mv/7EadiEcCXZoohU0hsoME79NzUJv5V2KN9Tzej+/t1CKgRLkEleJ91YsqyOfVv
WX+rwcWSmml0s7uBttZJciEjt70jTCpstub9a6sojZX6RUVhNqCRNv0h6u1IUbavkdRN+NiQIXoh
2Ow+0jKIbId2uZFxBF5mmFMsq12lQaDxQRIGVb/Xmt6C3aL0CociSZu6N0xv2hCmskqrNjBKTMs5
JrYTwznJ3h70j66EhBa5p95cWd/iOAPNP2Lpt/W74JK6ytYFwF/KrEiEUIUF4J5gOIT66ZRpYSJS
91LgGHKjc87zvyEZZkccAf3VdBS5d54XiXeDSlOYRsZHZfHkBiWIRuQ/8G+62B627kN0wum5t1so
F0rbHiNBoVzgsqMYqd4zjHdO6URYsZc4eHnNV+AhCxs+SVUKOKojZlq1aXxCHc1Mfe/U7V5qIi4i
vndkiw28EJDMPF/Ygi5AeM7OdpY27Nk4KZHi36kqVU2jllmcQf2dHmLctSxzZJqC7578CCkAlaSX
C4qKRv4GTK1Eq77IeB3EaEfNFurKsUxU8JgY827E9Q8ppcruUAHxpUjHGNpuwEFHaBXMki/GL/WJ
RgMJr8q4fONA5KcXWtKv3vS5cWbdfMO5Ry8zA+UEdAzK5Ohle2VKij6pZg/LvXghldt952A1TsWs
0ZDBnP3X+hKpw67gXcdLnwpdRqcOGkBwbN31N8ycYsOcd6wzjuoC6iMgROabXw3oh64lWc05VONb
DjozF4NrE6kq3wof6MjlvDLSbU5vvvhQohydovq2ZqYGSeI2IfntKIbjkBxvUwpDAQo8yId8Cv0l
Nlfa+SgW+nqEKTh/Mt6/dTP7gukkSJuiK12W8mkIFIXammkD825tOfXaD6UDE3NR5N1n/zEMv2VY
bYjUoQtH0qcYv9Ex7MXcZB4/64M0mqcgavPqYkPxqY7foizWIgljsYXmysxH63WWnWoE4kN5Ayhc
2+tsJYTbIZxTBXBaZK2m8y1fJmdzG1/vfEE22qI0n+jTWFELkXCX7MVEhmoZx51dEqcVzX0pQuEi
XbggGeXxI/fEC7mR8f7R6CN5Tt5P4N7rYkbdZIFfobKPtrCy9Eoca5sRWKJh6heH8oG711FdGJz7
KanOmNH6lcJ2YmnWWmmH2g1eDn/G1mVC81rdvpN3amAba0BPwTKN4OiPia3vSq/q8eFRuKeQCtuM
W8hH+wiyYUQynvCkgg2lmi1yDnPyqZGGTBzYqrwOyIqVpKdhifnwJB9Zs7d3B+0Yx4rPlsPOWZ0/
UB/OIoYPd5JlyVQN/DppI2jMtD7VwbVHYXZ+C2G+CtpUGmrbmwdHFBrZOPMVlGqQglfwrdeIUQ81
4D8OVtARLhbbpvoI0+Ceq3OKIpG9bQda8EIXr6R19G30dsx1NQSx+2C7Dsdcwos2N1JxpkOCn46z
YTpOL4NOikEUw6DTxZdqVvy3ug5lCrMec0eAFl4ED1li7co8xXb0zr8hI2xaFsJFY4LacKnUTrd9
rt55R4pFJcgv/twIDxB1kuIeFbSmz0RkDcJ9qllCXHEaixZ8V4u3VF6PlAmWcOJp6zoC/3+7y8oR
Ww7u5Rpgxe09xsFVWze1oBK8wJJI6gZnsPg4SubRgxZg+7D4yXhzUz5iInMis5UvSSG2oVgBGWIY
CZ0Jn7PdoK6J8FKfRDTLHI8qDPWkuFdZug047HpplslH7gk/dTk8x6OplZ2PwMArwLFpT3A8kO7f
KODhUqBmIw2+kIUaMAS+mepKvFN3NPw7GLtBuHuQPxhRNb246dY6YFF57visqKI1m5riwyZk0WBw
rUXcyAeKE9pvheQ/u/6sbc89u/hbXJSFfzgAtm05NVCdSZGz38umsgh9iCHWTOh78byMJr/FqTc5
RLfiUtoV793VLzT6JqQg3Wdjdn6u5zoUkUZdkjFYPyTInaly7GPlaT02/aOJUeBufrpKP3BxIrX1
zBg3WRYTmj1Qp1IB38WuuMIZB3odat+FtRCb8jIMlRgrOkhS6pOglyuXgpGQ4OHJlHxOONnESGPx
maQL/h3OErEqr6ut2R06+CL0qpmQJpVprxjXrMl09bXGd3Qprf0cKsYkVhNJ3h8zPNhi8vhiiI7G
4BelYX3kWfNYDdnr+N3GtS4vdhqp0J8wDvjGYsPgYXcElQ44buyKLjqBD63rEo+w9pfE657POJz9
dzwOk+qEBpwGzagnwLsWdG7H426Ic/XNj3tjrl2E5sgRp3U2wUXwx8KbgR3nwCxyX9/ijQvn5ZWC
uUOhho36QmUFnCJCQv5BwtMBYmKN4TRGqonGJlsGqbp+6DtSp8xl7HenWXZs6hOopTz5or/fCWwH
HCWU2Ir+JaVkbnejb9Dy7IC6qr5zy+08cxhfBu06IWpuowxsJhqU0/HqldSzI+27fKCm0oY2LjI9
9eV3+tqjoMWGXCvthPAB0RRTMee15aD5+RBLpR5jZhqbZESFE3gdq+zxUHbKv/utuOboKSqrHu41
8z5y/1FJSMjy8DRyTPxQR3U9H3Ar96MFC7JSHE4bVV7A8te9aWGCliVsXkHbGi3SUK/nxDuITZM4
DN2+v/lGpMgEyePUvreD88weqA4Fu3VfBKkdHr/EFiM3BN8AkNKhELEdixQb64I/XB5vMCC7bhLf
xWKkMyz0enJEM262oqBhf80b+JRVF6WWoWWDoEWiTy5s1110UEdW4EjzuK+6RgU3ceS/A/4a/dvL
TcUNAuZxfH9WTvYpcHsx7v1w0utOeZySuihhq8zrF0tD8hzLZZ+MxanPlpcs/joVhREvbPyD/DAT
SQrB96eRCe0ySPtfqjoeZUEgDkYCWgZKVnkPGbbbCrmkmOcoPeYQu1x4LeE76NZi09ZX77fP6kMp
F1sxGr/HEl9WiimNF/C6RFd4KHJDGj20pKKfxJoNfGUGBNrrOUbn06bZLoFdTmabRX0ie8qjQilY
4jJ3H2IxEfBli9Dg932aj/83XeRDGKV+JIABWPGUCNYkkmMzNkkdIRlGarL+apIh6PdmWuenDLcQ
h56zxmEPcW6RegTRAbUUMbPlur7a78GrdOnEEdi/Xs4AcSbosvZzaRZBYaNpOTV8j333Iusp8CoK
irKv0qn8GUmzPrOBznX5zeGnA4/cRD7WOiBsrxRaLlyzUUxerFwrGHl205SkKMLszCCEQYvo911h
nB1qFd5eJxynP75TejAIwcD7pEbLnOczv+ed3rG5+W4nZPXWnLKbsaHsB2A7QILEaaupDRgC9hbU
0OCNNbUED31LiH16b0tJ0bhd1/UKH7REsVfPLcRJzWe8LSaRhHBfjQaP3YqNKy5GwHAVdSQMUYi/
2lMTUnsLm8NNjijCfFo4m8IQux9RGT3GeWECfcpzb7l9Jt0qislnzXnztJH5efDyvdMi4Fup5ikl
aAAQjl2mek2gsLWylqiRuxkok/8DLRuXfzSqZS+1DekXfk6Q63xhpJFmBFPPc7QR3JHNexWS2f0N
Ju6HFIdvPec6gbL1vmv26qLPU4Pd2rQoedMbsgb1z3bMRFvYRY6HNlD37/2ANPCVnxalnLXlaFMn
KCof/Mk19z3ywDU1+OHZ8prQtN0o/sq7ftdUl/Ih0/3nCgTnk9CVb4BxefcoX/aPNT9qWgx0WzuY
mnV0uG1KCLSJZ/MF6vJb8MPwlrn+idmSeZvK6zfffchYvoVGceY99Ciy8Scl6qcSMfXBkU6J4lcU
c5Fzf/FktT0NAQCy/PCXV9CV3AiZJ/Ssgo+jRS1B7whnTLwj0efF1Vgk7OEMv0kV05enpW1nPc6c
SqoJnfSGBfKmm0w3JTzmBPToa2S8eUFBhy46C2sZhWeZVl/HPMaNV6Hav3TMGeuknqLsnS1cmisu
TiAuGFhDjSBkweNEsXLWNrknTyFVjRF8ogPoPexa16kzR7PJpyIbQOFw8LSZoy5YiyJlRjFyfd3/
TYxAS6ciaFMXHuKfmhndoUbDlUVJoGik6cmkuK/+a5bRrAed4cV59WOmt7aO4qvuTJorsD7O+q3w
BSg9yDuNzvatYGSGPQYntDAAha4DEjYIKI+9L0xKKjNRrF8sPLVCNtisS/zkOsHT2vJvEx1RRNwh
ru4MSus34GuysspA4b8SG6KarQh7J6WhDIUkzHvNFYIiKe0xFV2RoxoIs9Kgt2QPISAsSE87HRD6
nybOE9WRgU7aoZLNOW+/CJN2toENNXacefypjmhApB3PsMnqb8UhzmzlkG7JH8Hb1Fm2+N3MP6/7
ukkUUHst9yDVw8d+FCSCY1GM9d/QLTxvbkrEnO3Kkgl5VxVHXDryjiNOi2MWusECcRzYpUoQb/It
phtOWoU2MXR9kJf6wMUm6KMI5EF5/cEaobp6Qav7znRUU06DkSeEUOUFdXcJtFfs8GbDsmn/mXNu
s43eUDsI5sNZyvA9ZzjGI7qAbB6wBO6xiY8HpqnXHeIEcltQoiRdyAiwrjS+c7JmI7kWSiA0gkBf
92pBeyGMWNJ4s565UWGPBPSA65VzVYJpcBWAiezp2H3obLoJTTM7JuTlMWkj+MSib7HZIY9tgbB5
/7cEClz/1+cSvR2YDfhntfMlTga8kYSRgaRWUwjAuwEf0nDKkA8gUgzLorx/LC+0FjT+ZIxDbqI8
cMwaAxG+W7huTFg8Ipk8HGknQv9p2M8taDrafk/HQd5hkKPGYvJ2nlaW3vyMP7tzeCOK6V3KDpbj
48kSEBJ+izTOVryOu1uLxE4pUCttV+jyY6fMErv5irziFOYjRV/ImBFW913t4kwXD5jsVCwrphwG
htG0YLfFq1kIg/lFYuRuLQkJuT3ily8dsOMCXw7umvAOnHYxtA8fvgK4rRh78sKaLILZnQJeQUBC
uIt4uxY3OByA3isklkE1NA5CWKE32yjYab6SSW73TCuLCBdml3NiFaCyJxdMRtaFB7sx7+4gqMKm
swUXVtPBrdhab/el5qJPzH+UckR1Alb7feZHN6Dz+AX9rXY6CJklIXLgKCn+4rgxbydyyenlxTOk
xyx6EVpUoJmRA+gPXoM+3iaJ2cH8ho4rsenVIctiCDsekIiHQSODM5mdPnJmyxUuVH0YM++pzYu4
7fi3S0mN2AhEe+XFZAcqb0VKepm3crFKfl55htx0a+kDpdUP2ZVNeQT63Zs+UHf6Gm5X17kDutGE
fOFpdZn6Y8n7FGIaixsIHtXC+WFIL5X8FytlhJWVz6WIMA+5KBn8yArK3na3p3aSn4BzhHsRtafw
9GryB1BWwW2PqMcidRXiUgajCESUIuiLT6H4mbKcfiD0iGre+2vt+1NezTNjFr8Yuox8Cu2e79oa
jfbn+1Dkt3UQ8FBOpZZRpAXntShVN3VMemetIesFObejjUzeJnf4cSoJSRdCG5YDVo6CB+JdGi64
+pG/Xf5OT04+AwR8YuJOn7ZREk6eVEwAU0bBcOYd863T1L9ANBGlQxv2VGC6yEWD95dTzivu4bUi
3geX4Q0YmZVpX8REZYOKKtYFQy1SWMJaO9w8PMf2gLHjGkjy79NnGCstcfbp7RbR4CtNj3dS3fdm
dNsz1oBLZxiOY/uFmQ8UsYdP9nC1s34kjSvBrmjbdl/ojdBZe3xe+V1ShqvFMbje6fgOZYLd1YKY
O+knPIQ6sQraoYEoiKwgO7e7eAXUvmFAKUKwaRqnrDGFDmJ7DPlRtGp1RsDwzXyJqdrInlm+1c0y
8kMMJcieZ25TWCMP6QetXyl5p/pMqvGh3fYCnBZ8/gRFEJ2AmSMQiz41Nx8WnQec6CtQUnktKnht
PlBI23Bu3C/mcSaj2FMww9EveXnwH6KZ7Y1bgZdm9PI/7jBSFiONB4QiPO1cF3njc15f4pkvbR5a
EkMFhDk64JgDQv2XeVDh8YAH7FzFdbQnpI+cALYkMgmVfRcCsXNgQi/2bTFJjhqocXbOihcFNRwl
iYElylqnG7sfocOLkIswc1Ha4tAwHvkXa6HBQOhDgR7SWtHRsQeP8cLvs3qO+53cWvcCN4kmWBke
OwDT7cd2ziUgEi9rowlELCYhszF+xXTsubMJbObUkxT/wO+njTD89tBPXsJH6NsxuNG6uERY1GqO
jJz3NtlP00RnnGKW9qkfGltO3n7P1zWoJEkuICIQ1mxaBEi/Vi1U0rBo1Rbd80dpUTBYHmN6V5Zp
U/k2ZFV+6ZdStezK2IHwnMJF64zyfLFt9biryetcWVSsx2UeuCxbT9vfUOed+LZmSW5y0uaIhQV4
eFgX4aUGL7iTuxha+Ta04z0J4eO0MGg2M2SfEYoZkvGe+B4aNaA3dmMfG08UnR2/oDwoydWY2FtA
305x+4vv3I9nY2gnDIWbKCPpTwo3V/rcu/gfS44KlS+DmakP49RzM+1LweHJsKoscffT+Wl3k704
KSJaiPKRdqRG8G6fBqsAzQGWAhU9CacVrX36vmU6RuuXVI3Vq9FoOeNUB8bdS2qhItxuV8+GhUYE
548wAEdvwBxhgGVu5Xv2kqwv1tMZQwt/69UYQGSDQJVqNSkTaYiPXpG3F+ZhRS66omOrbLRBRHsB
UqEm73QMcxZU3PYSemmwe/G1YxauzX/oN5IwGcPysZQdLcZzRtvaYR0ZDGCfxU4xOJctglZn9TrE
qlLHkjTLo72wx/6KXNyVZUNEleT8oq6OMvbE3l+CIHHpqwA2UEGiXDQNA2uumd0EWiqA7Sh0keth
BwExw0k+06qBwvUO/iEEWYWTl7YdOuUDQnLYJqEedblwVZj3EO3Rv1fqkom7789A5v24FZJk7IXa
P2zG5jzNbZTIzQK/KoNNQT2wa5i/tOLQft9ueGnCMVU9Wqj8GaW80Y+sJhvCKXOJ+1qoolhD1oaY
/yHZitWnxlrqSzx1i2CgGewZRiduF6oP5ocX/jURqp3PEfQsaN37wdP0M9tNAB+m08aYD89Wz+Qu
ZNnaNW25IwRrYLt/wOs4Iq4ITvk1PCfHE8ZaoQ+JYg3M0fUXQNaG3LpZbjScthLAkaLcY/eGjgpD
tVSKsZSfbDUDFLXyNZd+FQYjhXOkzT2McxybOUCI1Ory/WaaT79zw7rMRsx1s1DL1X1Ld9IIYpyJ
9CGeuPHAQ1VIYjTrBD9UgMlmhrqc2Bx24q4+ReUwY5dRkyHAE53pZw3Xg66yOaOr7KzTgRc1iT9W
qyc/u3sFV5JZNL+0X6e17rfE0kEst9k8WupC5X/+iRUdBqc0gMZUEQi2R39clgJfS6xZ9QI3712U
GR7i172/blA8qwjbeG6sOMufkrfx4cRGHx6KPSSOIt5FsAOcI7vXnqitF7MYRxLALH6VdtJ8I3cw
zYAZ6B0IzqA3zaLWsHIQuvUXmLBAZYFyFjdcqWvb4XC9qHJMLugxa4onN4BgYEMfIcRWGxyGhruE
atfOqJ7CnY3TQfSBq/8160TPyXzoDZHYZVqpHAxz45Qts0ILMjmw1XTSfu7THIlXwNzC8XACHi89
vC9SOi5vW7WS4ZSVprrC/XzIg5ADeBTTwq+lJ+bKgiNeNZCsdq1kdducA7Fc3bpeX6RFR5TKdP2/
rLRBZcpt8hy9UbsfDlOT+chiEJvdFNtDhuadqad7gCkv7aWDDtOIBOuZr1a6XFrVJkl5feMecktd
gm/qSPHMH5ENIpFLIYQ9Q60eBy12aDKQX/Fn+D0qPUr5IcRQ6UOcbIjUQMxsRNGbLS3EQ7SBvjCB
QhrNZRW+OPBZ42hGRTVfpXFMrNKVtRPanRYLVIOMTNXJo1fX7fdLtZ1bVjWUthEQr6+w/aKP67HI
H3PYnLOMCg4F7bE/j37u8d17397YUt3ZarOWix5VWt6BqPRCN8/iSv6ctnU4mQtdbkQdoLt2qT2M
1yjcaPLDHWmTSok84TCt9joEQsI/OhBVUdYK2DbUr4e9QocP6Ai6sCrJHBCMgWZKxs7gsjFvuW5j
VB+ABEwrlWTTPeuTc9sNb7UsXpCc9kQd38U7+3/wTEZ03tzxAvjZ87h/s4iyV1F9w4HxNCjECwKm
jof4h4Pnbn/6YE3raP2tqK3BagkVJmwvCME5F+Yv8pSrzsoKRdcjj5hfFnD8QO/I0GhTWEhoUbIp
oN90lKvX7/LB3+h59Ktku1QFpl64HCMWg4FNuqZo9PFARkFXuln1wOlUaUUDIMpTK4nPFHwBGqTa
HdhllJ2/jjsOvghmnjPxwWCqNHaY+O9iysiEzkbgRLzdXiDhJ9yZbgBSOaMd5mgsZRltKD1NSrmT
mhvWtarxUc0fnE9guf8CW0unV8i985qHNA8/FK3U2WWGNG13g19cOTwXnrnQWHBmTAUZWQ33qsEL
mUR+ky7grFmHrb8SLWejERnnYXGTrwOwNu9ygux2OZqhlcKgu1fzky8UjIZeckuEGO84sMICHEMT
QYgFrwHz4EMdcDSGNpd1lw+V2wfJjjuugYK4w2FHhVJ/URiGabzWPQGQ+nhLntvDCXjwtwaKjfqF
UEREUJL0WJs+fbOxd7Q+US3CMwzfy9weNIbGkctH/qQbgqcJ5Gm9FlkXP06nDDRnV/xczfOfr9Xi
kpm6sirt9SyrCcdgaZW4lHzQyKEgu+YKkwWXbPjBn68mfKkv6jnFuNbEYtTiP3WMD22kSgVp1+ip
PK1Y2iLVDRyTp5TeA0UKwyY3len+35Ta1Mpesq/7zAlHV7rNHlnGm/V4MX5ce8LyNBCFMgFiao9X
LTCjEWBSlhgX7W+sjP0NiLsw+4xLtaTUIPXmHoUjc6kRXey4shW1WUxPp6EwdIAYqioA2h40Z0dq
G89vVeWehDlBSW4lb3tBLPVbufdpxTVvfZDqxgp2wJDtXenZGpXFkzZtT5+R/foL2m1D09BuiS0x
RDTGtaAR3d4zwGks1S1PB+SCakonvmFPc9KEVRYzo6kJ6GdG2pXOfDqzUd512DUjQUwvE/uzISQu
m/Py08cAWyDQmxHRLx8ukWVXCi6l/431v1dndofLYqH60LVjKPbTKnhcuPUYm1A8pE6zFXKjV3Sw
vd1PzDfaPD2yYVv76VohPvdVBXp304iylSDyYI/BHg5Y56VS3L1Jb+ZqVVm+hqSfD35wFVbQ0+Xo
oTIARB/aCnlLnw9Ctn0xyvX9ZI8BwoAKvNXEQQHhkHxuJu8Rw73rT17CMJB5ivC/hLa+mZN93Wjm
+35aciPU9xb6onC5xGkPZr9002eEiyDNduZ+CiIFYuWQb7VARE5VVeDLdqoB8bVvAcUaZ9oDXngQ
ZcOew8geYWYyAF0dofViRqcKWEMMiK2djif4hq1lPnv02qxKjYduqVUB2CAGC7LwUAspy2It9TWy
xTn6BhTz5mvD2S26wwaXKTLjUh5kkpvM0YBnnCSJ15wtxmpNyvnyOpP4ewCnvdohKLQR8tEU8Dyd
3NpqKv1dYwmpaPc4r+2YWMkzkqzNg2K1uinHaIYpFX0UZ1uaJnFYrpvdD06P8EWHKx6IlvVY7cLn
yJah+vDQxwGT2t3OBVi5LESGhStoal5lcq3ZRNWycnXATBVMiC5PVYCWGmdH9B/6gZsuO9B9FkK+
JkQ8lddq3q07k0y8gZsfuJwSSEwSva4/c+EyWbzbeZPCY/8QrPNq4BpIjhxUNwuMuPKgW5Fb91h0
Odaa5oK5Bq0taUG0wygKu8GhxBIlaaNec5O2cx3MJhH+erIgQ9YvBF2S3dQLedOIdS9eMffjlFhj
x49EkNwKy4f3kPS98hJ4Bu0Ly1T1/ozESIvaOPid3xIQ1M19UYA3YGgMt1fUrIlzmeXnC85nVyCH
YI4N9RoQCJrK9pCjmNkChwdt75jg1Myk9K4Mus2HlgFUQubKaf+Rn5xvMl4AoaQy8S7gNBNmNWPz
K45/YEx6pyRwBLXr3e00IxUgE85paxnPK1L9pc0ECmu8Jftqu8MELu5PsSW0+c3MjYaNNT+VykQY
+9Kolb/DXVGFoST8rtCxD0Gu6Od8KORh9iXbLcVN5EBlJepR4bY0yFVz3dcXAz6YA6F5PbsrOOeE
qi0aMfEHm8M1utYU9aIkLjmBWMDZbNjdN3+64H2xgr+HxX673hcfiltQx2j2OvErYjbzT+aW7GQ2
RbPqJNOBJXMe8eJ9WnxkcDd0BxOThDVpGSJB38JsCQ7bJLP4EMU9W0k0IcIXCZcgNSh3bnXs0bSk
q2lF+KEQ0DwC33mMGCesD6tDIOGREkqPGuLJcJJArPEtU7M2Drg0sfNQEj1WeU/DCzOVbjoOfaQX
SxvAam0BVd9ol5Ov9Qqjv/tJ09iJ4IODBeShQgts97eqsIEaF10OlEZQ9fe7oT7bePnHPO1e5obI
n0PLG7DK+Qto6WjyTApI4/5Q3p+2hiMWs+is4ATUSAsBMQLbKQZ5xIcvGA4CPIaqEwd0g4gWzVlp
0LzRTCU4/0oDPyVTf55hbQidDvZr/F3N4A+PcERKYhuDQln+KRnkWRzh548mN+YPoZi4hjUbSv8x
sdgs2l5cSPJu/GA9LxkMymuuLVp+3yHo90GWCoR1m0u4vTkHSNVnFBlbHA9EspUjDZoSmGaxDuer
m+EZVAJYo3IoWNDBYtA4qrVSoYEPZIb+++JDPjjWc+N30oiHkli1VkLu3S4ws7YMxSiYVpL1VXFd
rIIJyBiYIVWCfMRIIEYJ/7srSqDlnrPrKYGROSYoefMFaCyKA1p1CyFqgrDQMtZJW+9wmjkQoXOs
x0vz3JP6MCSsNfUn4SYQpQbwb4zFsXA6lzfpOKTY2ZQHcTOoOwircbmRCPWTsvF4yFFnG3TbPmhM
qNrqpaVgAt59X8Cgtf1uLqDeOQZaUwI/FR7mWPb1fy8cnwUxB2QIfWmiV/mtT3NOSP5AkWjs/vWS
Jk5o/WivVU0ogQ9qW6Jl9xNCdYXaiahKBVlUvoue6iHVxr+5gbvsUxs+IE87yolKCnG6haAZUAMR
myiB5odq8kHx6l+MfUfZ5lUmylIO88Yk6MJ5sppOk3VxLLqabi1uBKM73scvTunCqi+9TrMTc7Mh
VscHmFekJji1BXw9xTgXdBA282dLyxqKishG0qfbsbfvil4Ucz9p+1OGv52E4FngNOi/aIdL3Rkx
JDiT4IQ/FSBJJrh9iW6Lb9lhiXdrmvG7rhB99twlFHMk4PE/vClv7Hku2OurtnJv/dE4yHDrHWsZ
GuDek5EDgr3jo7qE+uOri0EWWiJLz1ngUw7yFtzi1M0VQ7Kp5vqDoE8liydN9nNtIIeK/jlVIHFl
S5wU3K6ANvejTCl+U0KjiC0WQoLeZYd5xfTCcTGKfmWtu3gigcPi4jBkuXJGNRwMVVT5JC492/YW
1EbLIE0LW2OwA/2fgmsKuQLdAF+DeHx/HszKAp0xx4ejXaGxu1haYsfEYte2HJwUf9SLEzFBROtw
2LJJiBV+h2u3NZzlerAZDOD8oWKlSvVsGGQMRlanaoDvel6OCdfVIIH9pNjz64f6jwm8tD/XquPz
yxJjz5gb9w+eNlPwBe6b5wEEd1Jsr8aARDomRF4KdX6mIis1EG5MPpQdQBJI6tEaH8+qS1giEPAb
sZXfuo6Jhiz7fZKMnofpfgYmo+Dq5vCvmFfhOgVFPZJhCZnB+6XVAoQopbpVEHITGck3GrcTZHgM
TdiDf8AssRhPeyjNiVTFelWCyUEN5Oj50gBbiQk/x8Vt8aB6wRInlpkHULveTPRM2k5epUNB9P8h
UWNdTP3gArmug2Gjq5geRRR4px/sR+SC6XNOYlNPXFOXBwUnddOBXyVc+DasykvAniJAX4INsfYO
9qr57ACbvr8lj2VdCIp0v0KmB69Z5+03q5RRPb79a/CeQD0f7x9NRocIAJho/XvWT2CzAwQu2MS2
mb0xMaXuZ6VzQ7DpkpiFy8M9gmBO4Q4k/qHE4osHjkmlOLHEd8spG29ZByZ8/qxX1GTj3uSEmbgT
yvxoxWLIdyK6aoGqu3l+FW2dPQBmvs7mvaTxlch7gV2wXH0tdMELBsXIjvqxIVES/V9TAMc1tp0n
YOB9U9GTCiu4uDNSYCIF/Q9dNAJsroze1kQ5u4WuOWWrlYTHQc6FmMqBKrB8bjvAcWFBi7M8Lx4b
FraBYktaQBFq+tvK+93b7qeFLGp6w0Sjdsn99KN923QY5eSS28AUL9z+dR0f9BsOZqzxwyeni2iV
PHAXEcZrdAE7LVGujiEOBKNNKjdqqQAoXb7wdf9P/sRcO45Ds66LkIPTpWIlAVX1SgY/CfEoUUIr
vnexKtjK+1YgCBlAk6BHbU0aySpzNEIdbbAmubVi2E53kHRodBbXGdtTh+C3ZHQNQJn5w4ZZx9IS
mfRNM3YMkY9pcY9lSzeZ2Gb+rA5flfk25Hl1pKFeZPKbP4Ul/TpCbSuocM7zSAUeQGTvz2mE6NC7
gC+mAwCKtAq40EDQ7rXtgqlP6pm10C0MNHv+mWKHduP8sFh7tkJ1RAlepNjxiR594t9AGITnQfov
VVwZzvUgYjRZ45gxnHwEdBMLTpM3hIGrSyj+mSuwrF9JO240oO2CTeUbHZoA4yjXSCn2Olyqr/Zk
e27bQ4a71IvxrvZF1Nc5zSBv6sXax8VCHa4Lc6VnxAvBX9l4trT98pXvXphv3Ew/hvbgYsl1kTbm
xuWxzZVsC4MZA0EAJY0LhtwMRnCFSHi6P+SvYS5vhKnhxucxmPEtecYjCsqofAUGxejjs+6pczR/
aboZz08t7nrSPRl1m64+OfvdMbUpUj3gcZc2G7fUrWLNff3wi1peHiqqfZtLb8HLJvGEfLtWkuZM
ag3/DxKZW4Bwt5HhuXk2o2O9bDmOQCyGC2qkyRA7zukPVAVSCN3/y1pfypbefIqQ7qVPvqO7dwzZ
vnQSB9LGasE7nX8plRkheTJf7/uxy7nN5k4o4a4yWA3C5DXHcCEmOWExmrR6ISvhW0u7JwZU6p2t
fy4DoHgeufQvsNgZOsUBEQBUoSv2LcSCp3H5aCf38rO2fJ+h8TciwbhvAYYX4MBigc80wZVv8FAn
8JWj+bxWMQ6RkaX3E0WkHuYpUok9FKe5Q7IjoQCmjOQmxUxJYZypC8/XaEkrG/YvF4q/3037Zq8N
nniYenQ3mPg1tIA+nVcynHwSJmMzePonc6SPLvpAbvSU9tqtuURpF4tKwyx1v9hmvuJtju3s0TGI
SkHw4Q8MWND+0qKJTxy+acFaI2meMCI78SzM7U8U9aqsFgNE7jz953XU7/VOOdh8+PzAkOrXTHEU
+fcFyb4O3hWZKyJZWgeoTT1KsjFh3hW+ZIWrA/tbmVwj2jaMWMGAFNfXXXc9kRGSfmTcYdgjgsl8
FLcknJ6f6rSSqHOrVwMfz/yBa6S75vQo96rtQr17XAKyeVejhbWs8Z2uFvi6DZCakP/Ly+/Wq2gJ
jChAsyV1L+UHLKRz8ssaFBmvgUvPsPK/ZFdyWv4ScfCYgfv1TT2zSDnRjFrw8Col3OJzsPQUdAXO
vbNHSZTl/DXHPduIDs/SSQRfUpp3mKOCSwLy9qU8sCp+mfk3AT8+xHsSqXtOWspxljThomajcEES
r6eoNq+COJ7nIhQr1PAW4fkooi/zAQx2HyTej1MBIwyhUGO9jiEwqv3j8jPk/7gM82jX1IFvtmWK
wzNef2EnuoGmXafq6iE99ys3d/GtMmLfz0IazDrwx2fbZQfV6Lwyay9CoiiBcRllNFoDu7Zxgejk
6rrH1y9G8ecbtH+8FPFiA62VNhqmyPTL8Xjiyugvsr4I1TI82XB+267Rk2rDv9h4UGmrt39eYSbf
F30XTXAGtLDLEdueXBMDWZjz2u6M7ohQ2QRWudgVokGrUfzjGaBpviWkN+q+TqYAcedEqHl+0PTp
/ivPcaIXBxUiuP0Y0/9v0++lfzAsm3kkIlO4wkaQPIdnoG9c6YfyBX9nI9qsFZm7E3AeQqnSaOAo
dVHo30aX+JGOrvlN7urx8kfNlZGTeH1lS3HUaSZNvDIfMYgXr+I3KaLE0nzPl0a65j0BtJEb2eRl
M3BUpP/qhT8WAdpJ1/lA88HdSKI95KAIlIIk9y3J7bE/QaSKb7soPRMlQ+3WD85YceuWW+NHJtse
8JaXiRIXWq1ir3dQKyWXueF/X03fZk+m6dhMfqJQbkJo5lsqFK41Ac4RVFaKgW1l8HkvVCAevg7M
1O4ATdhLpauu68KmPuAHF/AwXwOptQGk/xkd0DVjV6JcQE9Dv2mYvCFkjpuWd73CaKh1ADqu0+qg
Ktd0feTUHEpC/Ygd2qCehWqP71CzhMvV2bd7eMHthKFsBRWI+nsfGFfTmHvK+azIRR+h4XLMtgp3
0eGjU5Cl7Ib7fwi8/8LETp2c4HC/neIuuPqU+0rfAW1mW0XxdDSyalrFh2jm5UlXqvkbX9eUWhsd
rkpqnNR6n1gIAoB624ZW3qUGrz69yv/z2ib878/VXDXcUoJ8XUv01e4rIxlqmmE5ZrmWVa5BjKgB
gY8JXvT5Zlv6emjOqehpoqCQb6lpO5+4/25E9godirJL6L1AMGxYlMJeYHZwca8s4HGdVNmmESKh
H7386Cgb9ajMDrZBvuymEqNqBd+N4DHK+FK8PYBGA2cXfEk5r10RCF7uk0vgQ+xR4lO2p/izAo3t
80kMryCSmUv909zrrh7vlXFM+JQ4FWYVdTNOriwopky7e5tuqAgDS5tTMqZANqAGtF/bsalIbTcg
Kp3tpe9nT9meJcBITCJvlImBFACeIWUvrpeOaRsJo5TduTQ2OeJCAEsdMV/0dN5JWA59dZHuH7Ca
zb1JZM8TF2pWGN3/tefUMFEJ6ISoBt1ZSmRdT/Llb1EAFys4bUaR9vkGo+iMl6laeBosD9SXpSnX
FO63J6zxz7NMj63v6e5+ooCqeMkEpH0Fl4xL58U6BxcnEnvoPJ9ZZpH+mmhw8JmPqft8Tl1vmsul
mb72ZJ5U39kmA72/m+IHYzSkfMaDaEwxyp2ex8Z8gW3nplky9JS77aUDXXCMbYDeWKNIwmiJbMnX
1TAJDqXJXmvLr7aMho0taBh5/5uAZhabmWCI4JiV4TQyL3/gL05nDghLbWDF61M13LQQUBQCqSAl
Hn1PVDIBrsxu4Dy2QL0cVHzyVPByLAIVie/yFI2wf1eyZ/GZmKlcBG+mVDJ93t1ZPjfdP91T0BcF
d96+bZIlEV7Y+PRB09K5YJL8fURTtFd0OSU3eWXGEX8Ft3Y8rCZ/l1QO+sh2xoLhct81n9NRoVW0
mz7iAq8hbGLZieOJvZuwXlkNwEH3NuBT0wPD+o6NUDSFp3hXWKgaMnX1jzeTivO+IYtT+vnSD/UQ
82KUA2IopGzvrq9NjMu1cP8oLf56vKVELGEuM4Q/hdZMpqqdnsODUmS7bDRwwr3dwkXUG5xrX1vg
XIFZQCbgk/dgq9UF3ppx9Wk4ghEOjwGGsLhw9Q7YPHWpnJkw/SPtNQtgDIXkOj/r3H/nMM166czC
vPDFL3JgC+BE8rRS3FB3IxbRMsuwo+iiteyL/CAxSBW91KJr4iXAhdIYUFR9OTDUvDiqdVOi9DVX
f17mIrD5PeND54zdqYW7Wq2hxHQ8lmemC0AZF694ORAb1MiwZTPeJwqTjSva+HyUSOJ0ZUhih6mH
QLbQAYbyd9VrL/zppSieB9WoEZEqQ5xC6P27jKoxWgPLOdk2B9TK/7IrFjMuN/HwjQAfNAh4eUG8
btXJGmKOcZ0iY4ot2LPofKxDOdeeoNpBuTSbGkgYyL9pEW4BOFv3ll3nTeh7tHfbkGeOo0RAOVkK
l/Pmrm1eGBNImsx2+kU1mpT8AA8o5XcO/rCAFiPalwioOR2fPgI6NNziX6WzLP/TOhbaGZVHG/5t
NpkP+d40dRggFdAyx2ULuLu6n4Ud5rcH/wSz3DbfypUkOVnwyunJ7ckzsHy2ramVU1wCX5vXRtlO
FBkMKAvhC5ZFtTtlef6T+PYF5QqLoAbjqgzDnN2FrsUfXQAYKAeSHN4d/ujNxMCt5MrtgI4MQKNI
DN5u8rSX3Gul/UdfDt26miTdyr6EfHEEOFDEfxIQavqv2ZhSa5dgOHi1GbizLRTDoQUSTnudYB39
RlklHLiqZ/Qc6tTHV3x/6h5Ow63RJCWD6tl4dlZSFVhEJAlz2JyBvq47h9dkD7rYwC7ecozVdB0O
34mz7PdG5f3eVeeLTCUcj+vuhXDyKP44Ne7cW5DgLNok3Kk43+Q4okfaxUUHPpBXduV/XftkynRu
FQmQTjoW/bZK0F4p7ZGAZkJT/H5Qve4dcCvKd4War5VdujapWG4H1cxZgyFrCSw+RwBszNP13NCo
YUioevWanGeuoqjarG/zZIHaJNb9XKzAux4B/Q7DY842V+xwnkhp6BNrzxaeSeGT5IJvvtBEnaPB
ihfl++iBWwAs1BROvWczMa5bXpzlZkcYDL6TXJg3cvd7r+ycYAtyOwRAr9jMCYmxzXFAwrVVM5cK
pJhska41niFngvrAkLSs0sJD6XRV5tXTwuCo7/ahhLP7XnCy3Ro1zxYlxiMEkL2f1/FfokphW0GX
JUIZW0gvC7PQW5xx9G0SLDcrNDtyw+8ekgQ3Jyp4Umy7TrrqyFe3rAxa/QN7eNAxDYmFOKKucl77
jkRQXIcBNFZrPvRRskTNtjD3+aattOCF8joDujqdsbUT8W0F/PTW9rcvO1gIXLJNIldPiE9Y3Zxw
6A98Djlsy2cjSYFpyCZq4BdcFIBbkX/IQkcD370pOAjMz4KMJOP6n6aYy0j3gM+CBA+U8geBrANn
foD8cD+t92vQoU3l1gcnK3nrfXllz0VBV5fenJtxE9RMGliiWXrbyAOmpTyuuh7kOTDW89j1BLim
Yi3pA6C2TjRLoZSeb6u8du/mAoXpt/skp16iQ2PI1rurKFZXIsn5tQujAceeDZzsiBhhh6GZSme7
5GUlKkKRjFdXfSJ1Xzm15waAnj8TFrxcH4y5SF48EaNo4tswu0RjtQEMXEBiwtgs06oqhCK7F690
F8M1Fj5oXZZRteJf3cKJjmYh91mO1vTlI+BOAK5QRNdwfrC+oZoq+IekxDZpWBsmC3Mwl/2aHEv8
E+Oc3XNac23IuYxAlZ36/58+yhFub4EggUI2yYc5lts70Uhkihj8gkgoBdjOmjgKLYe1pnwBSxIf
l8nqGhsW6rV86R6QgjazQmyVKq9C4VdYBszkZ3HMTOR0UIbPktS2043C5yqIkMGgl+B48ocUeZ7E
6LG/GliN3nmuzdtjw/xxVuk2q22FBFFkSxenwXmo7YyOsjlDT8mgz4PyTxA8XaoVqK2ENxhbq7sg
UJElxeYKIB8Ucbf9cvwPxHrlRdDGVuyFuIJaPQcFIxhYQAhTD1AhvjeJy1MoHw6Tq8fC5m5f/UkI
mWrP7LYvOlGDsr1kIAvmZXowouFVVPJOGu3aX1OXGgGDJKg7CddZDtUO7u61/JeOnSjb86NkDKox
K6BzgAKnVuXljJHASdqX6SJ99rCmcEyU/deuaQt7vqadEtzsrgj75uGRHRYqqISNxC1kHmAXooVr
3WdL3gYM62MPXvm3PiWFj4AHWwpvW6x7J8g0mZFvIp2/hOBwEZ5Z7GpUg7hwv3FdRb/xmuGIMqG7
mHymsm1du/hdIz20Y+sq99oUcxUntadDM2JFtM+VfHHt1azbnwL3Ao7HVR0kncOUv/0irulTPcdi
QRrlL5BCK9ZVwM9SJWoOAncn1xUUMFoKQQ1FCDhFmf7Zw6sZ9KYOU7Ye69YMGI0zi/2JoAvjqbR5
8y7r/Sf16ZiXVUoko1DEnilnCIFDEHz6a2/9TYvvfk2wJg7HEklsmYzOvCX7AAvG3iDZvHccCria
c4TBNsaUzjaI9FyQODatm9REtofSt8D1XjPXcY+CxImp+rVoQR6iDkDCg1V8sOL5LUhc8SkuQQpX
xMz3hPcudUAgYIYNqSZtNTnSURHLMIu5EYyxFyGv0aT1bjf9yjaMA5s8vAeSFt0Oqk2WBakhs7+E
a0vok54it9ztsSiQ9jdUFYcYWBJKMSsJ4Xwsdzla1IQTQBhqBRPVLEaYXKPO+ef4eEPOu5vjAOSr
0zYyyKXOS7RPpN0otuoQgaxRnNz35/OIzZxdPIA3BceOFBLtHbNLB6gihEo710Y8kNkx+LCiNy3g
DWBPxz5X6aNsuQxH8Fb+wYfU14P7+bZDvY56dNUwKjPLsgUcj6U7KqoRcUtDxxRhrpbiSs4p8/Km
7qoOLCNzeZF7StfUnBlnwOILNkN6pxTilTH8Oddsju28Qp/PJiSc4zjpq8v8qDdE1gn1OihcV1nm
SJ7PDzma+A6jkamNkJqxsTEijuC2hzOfqaMQiFOFK8CogM0eMdla7Zq1RY+4fLarC9VOLbxmbc66
J+D76TL+ZxYdWgAhXAAdNwPv8QVlRijs3uYXm3S37PYjuPDJJNSBUKfYKCBz/HlacAA2EWcn2R4B
EjWESpsUgQxzrRMqJulSrRqrU/Dtv51/xwYgeh6dGYf8h8d4dIY/ngabglHlgpGy5MLopTFkKjiR
ILrdD+uVhMZgIBoq9ThenX2mQEO1OeTYDE9lhQJip/Tgq832ztuE/aoodE2WtDDDB97sNOBa9S5O
Z2adjU2KspdbZXzFX2M24xgmndkY/sgrXnUlwqEhKHfQmJs72uYsw38SwgJRxDcY+XMgKuBcz3MB
fGW+al3S1o4Eb9M+B6t/IL2bfYKRwbQWKZCKSrjLO9Owc6VijEnROAN8ffkLFZLoMbu51h8hrNop
ctsGsP7wPXJ1uwEmCdOqS9tBBTWitnAbyaY/9ux1uO3+WT6qiMzSSoIt2EeN2j/uF8FbQd/XiXOM
VWX+n5wX8oB8QXE2UUHn54wAz7f13K+kJbJAKMuhN+UcGY0KbQklZ7zUp0HF+J3IkuTFj4hnSA8+
9xKFVZCDSOt+KncdRn4eAc9h8ZKzodg+QPGtjnKwABE1x6CYtxZjRKePQOKnmviu3suq0TLB/oG8
zspGSxVuAFcT/3fe6lQ7I5NWCN5ybos0cJB0meJQY7oRE8k0YV3WfD8pXhmtQ42i5y0/ukaMa5hS
rkD9iXpcaINt1zDUl4txX52izxpJftloZSbIZSku3jSmI8rqAhuBbCg/B7ipXCA0gmnmCDfN6oQH
8ofwCq04QvvU6YqL/DzneAUMcqLulJqe3g/cnQ7AZVdZjJ6FehMp6dHq+VM7UvQcisNYjUwgyZCZ
UwS7R4MJmeDpDjEBQ0iwi3D3tzMLp1RNwyxapx0oK1AL5wwhHPBVIYQIVs0P289rtYV3+Tw8kQ+s
iBXv4yGJdnwPEzkZdFGY9hyMxlBrpXjC5XI+TTKKzXpWLiEjrCb81Q2+UV6vBbRSwbUfwpCRUhvW
HImXYRLyqVY8vIRqjmca/1rVXDwAb3K1ZXYDmAUP+hrA+BhNgw6CslJvudZSN91NYSAqqUcZ8PlC
MgBNwZ6vxjM8p5rW1y65zIjQKuwW4Rzl7KAr0+O9PU9GiJZr+EKU2CSenF3bR4LZtmVHU9yRA7od
g678iFtzI3URH3jfog1EQOhqc4fOxuvkgh/IRcdP7PHXO315Dkuu4saaJxdXMotJN1gdJPF7OjUS
GsBlx7zg2Fvcgm2p1p1NUMsmHWui7HN/68zswU6UqNXCyj1HWzIv2AGNEPxjRUfbY6MQqqlgNlzo
lkV5RHN5MiKT/NglRECjFdGnmcME/rW0OAWG8HWI15i40KroSpcbHTf2Jc0ovVFknNBbGIlEzpW4
d8s5Fuy6jMMp+ZBbVBKZy7F3SDDpiI4mxN71ZxrcJ0/BEzbC4cGx3j8UaV1yJOUk+lzhTj3yXuv5
2SleNlACKSvGbtqPTXxYNke1YGI3Inc7TesggZRjJ9XKNNntjr4DzFvMUjH9VnP+A+j2Fu+7An0B
4QUeguVRxdw6Ufe1RGSLFEKAix5zu0e9X0zAxLtAy5wNxTwjijlPe3cbkC/M/aPGy/HHclHkTDs0
TpQRcfv2RGSwLx1OzkWRftibO4kc8GIJUIJ2dJLMd4g3WXK91PbEwFZOb1hqsNx3Ht9X/D54Ss0W
eDiWTrdC7Lt1PsKkb2HSdm+fc43WLRYMMKllp/IlTNyT4apd2CXLaaj0pzjWomVadAW0QXA5eI1I
Y+Wu6lXPXbC+ue5VCtB35hhi5W9otq2yN8eoWntSQAghrOWO43L+gNhMSYI50sX+rF1//3IQ7A+K
E22WoZMh5ytzSpZqaI85x3yxxs/tB0sE9MKJuZxuTwPlMi5OhDMooFQc3086LKQW6rgV1Qd4XbP6
gkiOUe5b2IMKwywQ72oZFo/nD96i+UL6Z7XF4JrzvrZx8axC5ccXjW2eLuBd3DAgIQXgMLqU0zhx
XSCUFv3bxFXcG5enF3vaEEI34Q2C/1jFVfTJqK5HnrM+0AdbuBN816rIqwI1v5BtLn8Mp6cyAhcu
ygGDO1CRN0JEzOH0jWy1plCy6ru3os5fEdSDyw1fjpinutN4NDDBJlhLK6yDw4WqJ60udo6UT4Sy
6baoSuvhxF8jsai6gGiC1+zVM22gekgMQlCe4bj8liwvKMW7DzMFZj/H1Q9mY1d39VqPcmSYHJZM
gCRKy/s+s0kr+LcudwuKRMjOgKL/ZnqFPYDPCaoK06CKGROBdATlZJLKB/t04jY9+Z8q8rxmQSL6
tjRqnHL/8lMRqZcRzmIwjziwAdiOivoD81WtXLvo19isEhUHQZ+9yw9VYAdJ2RYvjZqJHXmDIBeX
1zRwtXk3YtdIQfTO3k07njZy6RNkDGafeGVU3TDgS3VkyqGFs/nKHGVZPX0Vw06uDAHXNsxaEn1+
f9BVIT+uAM6D64ErhKv+SlWgsfMpN2YAkTHscdS5iD2UQkzUUyTEKA2vz2jCp395Krl6CFJGOVeL
yW6NXKEndaNSxrCEAk5HoaZLJ5xQWikyA3MS2dmxWf4jMAD8s9SHUlRqz+i+u6ANI1fZlhAh2lgN
1B6uvkTf6yeG7RD8O+ZuUUHlm0phHQm3ewPqjcD+o7olmeyHp4UvAA6UErc7KxSIa3oZrHl6S/sZ
wfAFDTSoKuKzp+GnvAABtS03oliCgy/Iqvdew/BuQ8YUxxKxensLZghhIKWbKx1CXq2gy3MLg4un
yFi5P/pFU5vU4bF+tC7l6nC3SC4Uc+QD1QgL0gPuF89NmTPV1BEDSnL690Yz5KrBeRA2vnNjFAub
lpP0ii+axbctIkgjtx3D3N69NexGGV3V9ImDekO8HSsPQcJtb4A5ANOaInA3ivW+dEtQDp6mJkvC
8aK9Ms92/MMA98BOYnDSPPB6pNIvJ40J9U90rNbQ/6Zd7jlH1EjI8dolM+jNBqQnFxLAYt5GOFfn
FDF1MKlEVZlCUBSpLAecCSvbCpUO68OcDVLE+nbGgX6YRlW1VNd3vvjMwz/3MTOWHt5nn3lHKXGf
fHXGT0HvNaQ5yxfHHhVX3hEXJsHPCTqp4z8y3I/yzzg6tCmqyoEn7R/ajxHfY+/80tG49NzrM6Ot
uC8rapPAMawS1DqtyNY9H0WPn4P5qpR939JSQp1rFXRmYej0CBPTQY/ZC7AVkRXKILd9hPdrlsXV
K+J75D85fxKflqqAr41TGFpDWXNO1wGG5uLv8bHvljPyboRbTg85wn8h6H+nbWYIf6rHX242X1sJ
GitkvU8vy7uVgVq7+8uUyI2ZBjkM5G0i/SNvNRfVy6hzM6pE7Sa9UYbfG466yf367ghyZUFlNVyk
pEK66NJwrXoigwjz9tgCJ18QdZSQKwU8jr1B8nG1RySDXNziXM6qUgypYPL1bfj5K2geRYN053JG
1TcHtLC7YMsjyL146vHP4xFpPHtZmlkQUaYeM0qFeOUDwstIZsIISMvsoAx/3KJo62xFaD8GF0dD
BUdBJLtFq2tIWlofTv4OBc4mEh9qUM2zanGl9mCm282G0mM6NDdlD1rWVbZzCeaJJEBIYwwf7Cth
GiGQWwHFhE3+MNiVdploO2lPgNh2pheSoJ1a7cbWKuo8sWrYYxH9LxKjFMq/vYCou+CvkJt8PlTN
2Rzi/HqSvamib4sY5sPXZQBVWPPJcCBNMkG+64EXBetWlJszCMzI6bVyxMA9blIaJYHEL0ro9m4A
dRXwmDbtXkN84Pcxc+Y9KSGmafzJwk0OJJqBE7Vbt3Xm0rvIQ4eedsyLdGkT4wMLNjnOSfeV55J8
82tFp1ZJ4p1B7MdKiJBWnWmd7Ibce9A4ZnyfceHW7tR1tzJhwPdCfBEEWeM/PYEkXenLuidhx2qc
a9hLzWLVGFbkpyf5YZVsA0IYkhZ2KGD1sNSWVZTZx9QVq9XZrH+yDOx7uP3HmQ03RamhhcIgamh1
KIC97kQ9ow/jOJYXVD4MjnLGlV4MH8Afc+QIsURIoY//53Qr9+/cR9EaIZbiS3O5LjAG2mPkpytb
RNwkf7JL+LuIjbkeoaKG2Am8Z+/qdd/DKMjznNS42yxU6EV0IRGlQbmCKJ6ivRzLSOsJqZplhXDF
gBt7eG7jMdSDN3Dvbf+6nSseQxiVi6/+pR0hEY2DBVuYeDXoGzUDsVyMIHHZ/CHH91YBx9JYUvq4
4HT6LJ4GhNlscF+JnUmznt+cepyq1eWrBfjJC1jJf9S9E9f39r+5s41ma7YAaoDcnyiOst3OCyhG
QR12Mg8bxB1uijqePWBDb+/CNAkJ4IbDm0eGwTzWWRBYHJNN1g6atTkDCHrt3b6kNwQM4GogxeRl
yEHErfx275EmEs8RlZmMon7Sa5gQzGlJwIBzNJ97H2XgvI6b/XPqCE6Gzpg6jfVziFJ001fqBQIE
TJxJ9cQfNOK7kHvRgxJiqO35gwpbbSDccRlois5nfkd03Lh8AROliVz7bbWoUbtdi4pKXvVkCIno
iLMT6mupF618DtwZkuarWVwVyA41+lFrxHDyWWvfVKJowRlyw9aN4BOwWXzqufjV3W6uPaveywEY
tGL7RTlN8mqXMtE0w2dBnkJtsrFBCk6g/G7qjyvuYEWiqlimz2eybZzjSiEnwDD9b0X5fHB5Oxqq
tSq/+wmJcVRetahjrVm1RN7ybHmSAPgd8uRwcek+BULPlf0R37auRTYRwpsdl1sqldhQ7d6ZspaX
ZkRyDKUiR6NQ8rlFEWJWITe1RR7q0NXT1Xm2tmR6UEUPVpOQZkJZaqbPgbT2+m79iJFVcklV/hkt
Yq05rkwM1oV3EsHNec/xdWvjwW4fIjPfQfpjtWEHj0wYAwsqBySMXZ6rdOMTG6NivtOdLWt0fy6x
DU/YAJjArbaRsQxlpzo+uQWqGzj+7XaBidfOneBvB0X6YbVhi+JIhW3QPc2foXlo1JIdayalz9X6
pLiYc9w/F0xqglrqH2uK5lzuXlRyP+9WxfsfFhGi1EgiWPiXcYVu5Gj9i1Alh9EqYul8U0uOETim
liaoEaWWwxlmFRbYiVzWwrUL7CFAQaDXmomiY512iBRyw0xrOUKdxM73wMOhqMxQXyE3FOp9h5UK
1nukegqCJN6OJqjda5kNQFHM3gcVyP6I16Kh+eZVi2Kp1dDxmxjsQPBdrrydfrM6o1+oIO5dme4z
/ubDZxG5UDZArlCxSVdhrlrQ7ozkmXitkmZxccxnRUWwL4q08hPr0u5vXHT3ashwyPmXB+N00mQ0
5KuQCnKo4+ZkTuma36jX49Ull4ldiqemJdXQDz63CqUFAS9CkV3mf6DkXS6FRapRkFmOnHvONOtx
KHxIak6glaYVOAeS3fTz6EMcr4MqkwDElNi8sKWz0I5R/f1CcVw7vFSXjtmBLzZu1rgSkD2Vgub4
Ow8ij3zZKUd/wx3PUUe3KbIy1aboKmW4OSE3/MYhRBfihPcIyLD8qxE97QGVvRHUypmPNXiBbs7G
6gj/4WI9r+4S56Jo9EsLPatsm+10RsIAw0OqW9l0Dh4d0yrt5Z937fZAbPVt8eN7VpTG25UF/5uK
bYq7wZ54rwvS3gTSYY8jNWyRDkbYaJY0PPRLjByQlevCzHn9f1blpHPENf5DP/+gVVDbkMwNbpCK
dd1DepdiXMHxCG6ugcLOAiklMf3QCadWT09z1tDAMOdzf6J7fP/ZE735yGQ6HK6KoxCv+iHukv7p
l0bzL8/IW1Qjp2puefAngF/xAeGAA7REzcycYA4/8lyskT7aEf94ZtcFyiOU14upRxOUGfZB1hWj
PC0EjM3vCovuXHKmnX0+UFaWMgE/qFovH2CfWq4DnDdPsJUyxnG8/7Uz2UoWGLGJIomWwzRNif/s
fCmN6O61Hj8vfbU/MX59Aa0oX+OvmPpADrf5FcbRp+V5cYJJFuL6I9icp2x6Rth4P8xHKLbP9iVs
rYf+wKv2C7mOQxl4smijxBMrGLY0zK/IlYj/rqHD3NwJB0ruWOc3zjM9u8ytYhsD7FV7wGl6xsH2
T/L1A0sI5Cr2Jx/k20u43E6xiszKhPMPGtbpqUdW/WO+sSbQDsLjzewhOUwivAFaiOpgetv/uyJW
4Iy10Ntp76D3NqXgquno+ig/Vq65vu9tlqK4vZ0nI3G41VO/BjWl2wePA8A5V3H0Oq2eqLZGmRKT
qsDSlB4dhh5sfanc8XIzaOusinYiqihxBgPpYicQ4SfHE309Smqbr7MH84rHmhwOhQj3DvE94pot
/U5+7e174MU9Du4vDLh22S+2Mxn3jrR2A9H+V37A/IuMe7XkkT/02BEvEUlMIb17+PEWS7GTyheY
0elV9CCfWtaP9RY9Y4nTt+w4qoMN6+XIAKSflYE+N2S/MRgR/yEmmUurkmIOLQkr+Jsk8d00xH81
AVbJqaEdhpzWsnF6lKxWlOvdft6Q44kYubyIBkSHzA7LGZSwouehTLTKHnE4OOdoVBMjFBha/oOz
eraIetlQPobG2seQ7sDdzFrC+zJGlCyUMAx8WoRFljF3DboHgayoG+WJ8fqKWKzBr8GRMAB/+0Ge
q16LZFoVsqaCBQQG/rYi8Ydn1WMB/QS8ZNtT3Cd8TX3M+ObZyN1ZH4AO7/TjGU0KSyXdpZgBEzV9
L7Zc2ypK5V0Hq9JLuXKTPWHVr/eaJydbOWriVJiyw8wfWe7UIiuQfhe+flHlSP+uEpg414vIG9tf
AHQ0q2+ZlcFcmfaQv7Oh4llc5CO7IpogbthDub+Y9aJgLCbwFC2w3eoTFlVlspsfWhHWNj01e6DT
5Hh3wkmRGIw3SQwtcMaIMaOlEqzymNzVhCfMkPPkwYNQ+GyO3LXc68XlIJ9r1dMzK8l5jLBYSx75
1kZ0C8VmvIZdR9N0k/cvuy/YFhowlMpQg6FsMzx2Jz0Y1Lhd+f2zE/+toUW4kxwoXzfm0CjQakx6
huTY5njnleNxeKFt6WD+bH7UHdRRnKDhJSh5IIbWSAyaZ7Ugh7OgH+VaeK+S+qYmLA3Y9iDUsrHu
6XMOAwhZMabBQ6Uu46P37js6H/ndRjhB3SlWYUhr9IQgIbhAN+OECtHViOMfEMcQh0vKeqa1VKAO
hmmvsj9fE6I6/Vf5i9ZapyVX9T7GF/kI52oBeaNmU00vGfk9jTsFsFULRCQPymsbEZv3A2Dc5VMr
QJ7p8DK9G2mK4V2biaMl8Aj6lcMprfUIRWwmZd3kgxdqCIbJPdLZte3sje7OGAZfOBEddN57NydK
janlkZ/xYTXkGxi4i19KQG7mKHJRdJL4tvCY4H28z74K2Lu++/rbzLJ/zW7fhPoBx58VlXd/mGn0
MciH5H8Ifsd51RmtsaPjdmHZxr4kuNWPGSVST9ozLgod+OVqYSs8V7DF6Zd8CyWvyya5uX5yQWEx
jpSrPaThBO5pLJcLAyzUcQY9fWZ7IvNhUVtZQfQp/2On6Ob2bmuA9YNWzPMpJToiinkytXzsJAx3
ULP4csp2IrAnEaOWdYBiOiSlp7ZC7FDdEibYwNUfkPJWPwoKn8G3s/z7pQWmrN9PzFm5SZNy/jZJ
UrgKrYxJfcSxKn4cVEmlyAEyr5U+ZZCxA2akMe7VXerr2yC4znkk18bJ4h2Mb/2iwmXESvUY6nLY
UWzraRBJoa0JRam5RyCz/N6AjOzGEHNlyZDGadYQfwEN5Ne1fbcc5XEGvc0/pO408J556eYH3Di5
c9wgo74WClp+Tdz+mxJTnxlF0k3GwcK0SHQR2FXIJAO2P0VS8aujSG9yYju6mrkxEACIa1BKdCc9
oG6YB5PtY1zvAlzqqH+Ve7lpdk7fnpQOtdnJ91TvhSRkdQg2DGEH6oEEPkV3Fy7GDSAT77CQ+x5J
MbqSa0bSNeaRT5h1kHie/6i27aUXkXa/MDe5lTKF5wnDHxQU/KZ3QX6h0M5obauhantFYZCLXvHv
9g6/Lu5rMtLE5o5vLk5HfpjEj5VGJ3NcmKHFdQLdE+gwmPiLzj1bq8A4Du5OxIcQqPavE4JidOuN
McVm9dDs1IdsD/YuB0UGQG4hsINnkkOVFy+djkbwq5cUNNCumcZUWdzjXaRr8b5x5FMym3wmh6zg
4/rh90u0pq1UT0h2BLCKu5qi1jNMsMCrwmvGnrbRaf3pSdnBzVn1ePjDmHOagJuWGdBInU9LBUzB
dGVORQ951dsCSRPfrqiEIcMNyhJMcng0HDrWgNI0YY986wlk7/4J/Supz/LgwwjEJqY/Ddmroxl3
Wl0MjbJNeDWkk4o+i/ua0ryoCNSs0JGuKczPEuHwEwQaG3ufjaTb4m4zZ70z8QKPP3t8GLpvRle2
89viic/ohcw/rOycwgp0DuJoZf8bOmkbPY53WX/VqWoEOilw+G6q1MRqviSueOaTTzzBZzMoqbwb
mETZTD0tcOBC3kLO8UxsiHszRHHo8dQwKvj2nw1g1F8TAaeCqJmqhrh3iWE/nyKAD5OEWA8XQ5e5
6EgQLPOSYBFkRhekn9P07++Tm7E3ecfc0x9m9vZl+rBlQj9lFRFnZKK50RTPqqQDTasiYYmwdvh2
DAFxTuXU/1AmAutvCw4GIB6dPlfBqpc+x8vKeun3r+dE8unwqMgjnxwRuxqdhEfZi3q+CtX4LwVo
+QRSqO/QXCbmFO0ruc88mKyz0qvjOxzKdsmajKa5W9X8s5ROwaPQNyxSpfSwt2zWeqPfY5b+t05V
TSWaUSr9gsG/2RHN3YnR+bocO/4F5h5f4BumLB6J6qlYy6nzU70Mh8vfRhFcEFD365PWlA2iI9Jr
PqY7MiEb3D1Lqd+EXayYsvNuJwjpZocBqmbhEAnYqokKTFv0A7s+E63lkqf/pcf1UaMJZIED280o
WQECA+ytEWOhvyjDSlR+818EjX7DrrQggkF3wfo5G/buFQG9dCez5/84nmoBztmpveNlSG+dnzDB
RxwNU+r5F9q1aS+zX8yU+Y4AdYtloKocBJ7XXePpYtzGprnK6G8l1e0/NqjnawjhapOiuyWWn8i+
sBub8P7XYVplaT2+t15cV+p14LUvydfrGnmyBz5W1TUvnswipIJPm3SafV/udezTFV5B3AJ0gj0E
vsxJkrdfUxyn09/oOti8R1qHVDHKW3mOZm267yO0TyqNI5cSx3qN6itln0CvcJJpRTq9kGpbP1Dz
wvQyxOmkmfcnqbMR4pO5pAlrqZOhHXkGNhzurDlPazK4j6EXy7R+jMG4GhcbjUtDmMSMA1U4DfEC
m1mghtk9NDg6yPIxMqfr+RaHLsOH7BI24QHOmkZ55tt/Na4aImex0ahKpwK/4ysW9/65xL+q5Ayp
r24xGNlbGGaYDqgwdUOVcx/l2mL04VQIs0T1cGK4vOB401uJHX2H61Ni/z+SwZPVQ4XmJFaqrNE5
/j9eUNk4COsSM5ootLsrDN+DVmcJSvHJezb3wWAWETK5ExXa/a+Y5cP6mKvyK1CMWEPtsExE4WF1
Tu/qTSnG6aFsPMA61SjrAViDtpnDkHTQCl4Dn0roFEXA2jWTD6mcuVK6gv6B8DezqC7OPGD3k/Z1
sbxURaWenxJyWRHFhxjcWRK5dR0ymfF+R5XveCul8gc1vX7/FTQJNhNLqkgj6rK0aQd//WsYVv+q
9TZqy5BhwxsXWdUEx5sgJS4Qblw0hqeZUxw7PxVS+2FZWhi9dOmItA7Cjw0cajTpV1XHJXg17sGL
Bpa95zWgqbofbKGXcbPM0vk3z3sZcNbHys3wfcr1X/h3GMb3GSMNNQtVmJ2XxwkPCzJjROARz4I2
iz20ZMr0+4Rh5UmR4nh2kmS5cJpZ2lYJARVT0TOE4c2PAULkqQmiKAcNbiax6FjcEgdJFhA58OGB
us2wwL1GRJOAtxPfUO/BHt3oS1gevXED4DAqvMUDtdHorQCjP+wWLNYDkbQFKDbF+gwlKNkw5ZwB
+WnuimtPqNt3dzPARSPQploKsX6h3OuH6AjBayhK4poLjWsr04OS+eSECBT/Q0ezlpjr+7qg4HLf
HITyZwlDeFDv4fHYaCp0vZQPb2a1S0OxLKYEU2gGsLXRkDlQLI5DKeTbtuOmiIkY7fSr4sOU3nYw
bHqNoiAvQNzjWcATDomDRRqTy37B4YDD9le+NI6lLcP67EobauEQddDcemI+NtZdwuVAGp1Vwmqc
Kqy0Q12ciR1VtpNeOEJBpkDbGBJX6P4jWzrx+DueexZioTcGsEfzcRFJecHMFTbmSHvmNl2C/4Zm
RYPijyFqATtB9Uoy2+JpfESDQWtFDzpe156TklCqcxXNLVHJ9Ev6XRf+sY2n6IqhlmF82Wjlq87Y
qnNjjCzD93PCoxcIy+0FnyTrKed8ArAJOqyVcaUrLSQ3/x5/UvmzOFxg+Vw14O7fhWtI6k64KncP
JNIQ3URG/O7D53A//XzxiWysScLR5Uz+euZ875kg99NrJyPUNw3DpRGBIQgb+oOcuFFyWteqjD6m
Suh1euvKQiE5ujK4nqiBncu+Ip4kWzcxKceCeHEh+1OE0ne90xaROoIS7j9X9+9BltYgZzVymqcc
/zJOIVu79dDzIfQxA6x4+YAf6bdHZwGPzR/C96ucJrDPE+UuLAq0YVfRJkmtdlbFCBWMBm2A6aBh
HuEjb/Br7QfM/nCnSDyvuM8tQqfkT9Xso5vvEgmzB781W2slPgN9ULI+ibFdRBcI1uUzpJmGSGh5
KcqVTzh7kgy5GkMw5PfJzluaI/JunUZW2fB4e7Iz3Ke5PS0JG5I69T90AP8iKx6W0SZjuZA/20Jd
e130e/CNU8sRG1NfuE7epo1zG/pEQuRmcXvvyP6PT71/ahseMbCNI9+ph+U7BvzkeAGcyWRRlHyl
qJGxIznbX7bT3FGJyRH032GZ4AwlBiscAzhuVb976HF7u4j3MD+++JZTQvaAtdKm/BM7+P2A7Bwd
+txFTsv5EH68zYvOM1IixluU11Y/oj3pSetaDgXlF+kRG4QQvMkXLo+elf3pLxUz4PUL3gDocSHg
vhuO3DejfFa0EnIv5VnEG0fpGCMqjkHeI5E2aqIpqRuZ0W7CGMfbybUhuCo+PDZ3JFV/dAUmYSf8
WukqGTgxHhMTkGLYVlu3Z5/3Hs+D/Afwa7YXEuOcfn0hlIiwHZJ995aRIXDkgaKsyztqywt4KR23
xq/REioc3RH1rp7ygCn/3X3FpEPmIskow76llo2/kgWxVgEMjJe0RiJIubfgsC7XqhCi/nbueSU0
JanP0gvI7TB2xisxaDE977gvZuGFNMIm3gbJWpv/i7R1BApdCPueHKcleftbNTAocMO1gLgKWmHt
6uSw9LH9IqqsMdaQWOYUjxe/kxwxJST+rFRqUeMUS7MckW5bcnhM2XgN2DtCfXuZyGVvndGKRJgO
pewuj6EmExNDhb3b4jNw9mxJEdJr9i1rj2Co/b0abxiF1KlgYb6Odu2B6sjoVUa5T8cvCOSVHEIe
lNaCvmhbbQP/N/T7IJl/6blX5ozB8be2ML2AzZEPmzrMbsDr1/52d8GyMd2zNZTEOxPKC5B5icza
vgN1juGTqtxQ0JjFDYp7igf4n+nBE0rU8FrDF5IfYV0wyHE0crK66yuUK9ODpA5t5jkfElE69L4a
xIillaXS/FrC8BPSHCkEm7WsZdmUJZKhOmgH7Sz4N6Y4nV/NaghXUIpD6RIEVUjZzt9tpJHX8oJh
DXd5p2ov8QFevhYhur9QLZx/s7w284b6HN1vdmEG0RLAEqMJF9scVTA8+iuOz3wA2InYIAZT61kg
AsBIf9vqT+zdgLNu0ok9Am7RRKqdPsTB3IfqJazlkHAC46lHRCqUtzaUf3jGCjroPHFDi8vciYgv
pWgAl3LAHYcoco8JFSTgZTouw6o+b9Idp2uvHuGg2Ra8Q5i/x3n7sBsCyR7RLrjo3D7NuKII5cpp
v3IYNa3H9Ao8tTbnGec1BtxfRdNb/qIXfZpuPHPmelVg6XPRj9v6fx00yFqgyMBr/s7tKiQyZnmk
I1afKvD3kx7Onda2qyMljvqDDkeQJHVHFuAxCqWiLGh5cvUND3ltbScUHZd0JgnSsyJCv9qLlNu/
I+n76SA1G5uD+MnsPaoNbFu5d1MXK0zM8bQ2mllTEKURLoSvYY0/c0vqvmRZHNqE64SBNduvLZpc
PWVeTwD5vmIMPCOrxQr99/TOek+1jTbMiG6nmzAnm0VNCy6E+yFim8cY7UojpxopAyYCVJZ5Tj3R
xaETfrpl8bWOzjNU8VSLM2q+XtIKafFOgzDyn/cLf0Zgfp72ZRiM7sDJeNNu2Vk6ndNRm1QuJ6O+
fSW47U3rlox3MBV8HLHX+dLesUV5xYJTuGWEW+s2varmQGMR5ZaHv2SzIEKpo5Y7AJBFSk38fxp3
0CDEqR8I+x0wquYv7ZOse6+6zwV4IYEaj7i7Xxv1UPK4GdpDucvECwrxP4YdjiQlXysOfeMAOsOy
YfM7CeOKYphLHBRmG3Rn5PB7qNP/VMEpNpa1OpGthdo8YwIncx9VQHh3IaMep/zMXK0WqdM410On
wkuGjPunBSBG1gL9D5wZdgIO9M+TIVpOXPdR0bCUOLpIEaHpp7EHM89gRxSvFY6kNkZDFzu3IKUP
doYFDefU1dtJPEIUXvazug+L3A+T9so6Axx23l2YsA78tjWRfkyt1z9JJZGaeygc3OIUYAEYfYac
iu4hNJI1Z/6iFsYg/YDEIEl8pPo4W746egqxddE2c73eGij4YLgPRlLhKB7SBIEK3ROppZk9780F
/l1v73eS6eQ9ZRfMswN18ddTG3xMHufPvHWAzbwlXThXBXk/U4gYk2ZkVSWy5D8UcvzcxHm81IKK
D11K0e/Xx2djuoWs9ooMBS60Rwk8A241S/CmAFs/yJKvJXkXbRQGIAZpY1Sg8LqCkVtp69y7UoqV
Oa6NTmRnSi2V4biBLcBnRo0HKnjheV9m5Y5dGYcX0qjc/jYnbNJWQVxipkVHh/v1ch0WcJ2SyNNf
JynbgRsdc9hZ5xUygf7FMu8BuOKBwZYnMG5ypRznAGzHfyqnDq7xtnSVpZvfH6x7GU0msCoe20+o
PLi6BcJ4f9/sTwKRJZMxUeLfVFSsOdiW0ZSozLAv+XbprGmmXS1Mv+8KvwYgg4YVh764LzOs5z4q
ZnrL93tDwiXfO/vPdSx4CBVCPALvKENBj9a2AEkHIQ/SHPUzUhnKNHM5q5FY2AreBYYdipQgQbbN
wj+RNUYQ6X/tJSojGBlRO+snvzEyH8y66hAzPuEduZKHtU6gD0t/To3YvcyF3uhU40wKx0AO45NM
efm7/hN9jH5t4hzxAM3Kd7q003w6banAdciJMcGvLg/72qMXreE++uJGeyq932GTBTjGyrw8sI0S
jZbEjb4Tk+xBfRVVfOcx6ECclqffbY2UuBBSG4DMRd4jcb1oC857+X2yRRPu15kvJXFlmvWFnq3d
IIgAZdAzgdglFTkP/bFv5xObOI0Dpo+L1ZeT3MdiKO4HPVSe4yHOX8wsQ/1HYFZHjjVHjQwokhna
8cf0uXwwWa3KQGUeSm6IuYZuy+p0E9bSBrhbP1VFzc7WRkk1Y/ZCzn6yOz65zO2mCE6GDxPCevnI
baDy8Lz+YTxN2SmAMe4H7eGUsh2RbYoJexXhUHnxdp6qwcI3gFVOsR2nMaB+lhmhCReFCc+Rc4gM
hsNKUPy6jTUuoN8xIaWDM57as7Y3uLypwAz85O4UQ+IgUfNNMNRRIF36zZum8dhnqbP+l0xY5Q9u
dehKzKv5oB25T/iY1JiQ/IVJ9yfTKjohuvBtSIgNeTHN6waofpQjBg4Wv8WUw95FEZVRNCmMpEkD
KsNogc6TD80gAaXeJxM+qC0URd0IyK/DGozKxqaolGiRulemqb4Eh9wNI6nSb5Fja8nLcsVSDdtw
PHZMk+qs5X3JIU24IA3mtyRtheUUrry7j1vcXsaANcF/ZJD1OpPsHrGhhJ3d4k6LegmM4EZDH+aO
ycfPoK/4/jg1RJZJ3P4tKLOYfHQOYUpDgD8TLrVkUp58wBAGD7CMWY72NYMclLhNnMRDvtfRZ9g/
88PeQY5JbXUisSHrjV+judD5muOsdOAuZOEj9CzYOoqiZRBpcpifr5edrc0mRG0t+zMZqixW3hq1
5DYHj02qrdsc3z371kJKLtztbsiDWrJ3P0qvSIC7gRJdNg1kmdt8fW6DNzTPiZiOpOYFDKmT2i/m
+9iPTupTCzc1V9kejXaOxKGyza3WG5m8/BoYu7kKcPUhdInm1iGq6vvibEDOwPaS2MUp79agKVy/
KByKwbs9xBZ6DJcT1aLyOVbStNUBBwYOCjfRlkNiUJS+Yr1Zhr+uWFkDaMQo7zBu5gJk3dxTj9M8
m4krMo7HzfRBJHGjPj5iW9tj48C4fjYrWvfPDBew7Bz7/OQyW2cmSledFDOHld5KUYcN/reR+BCd
lqf4WVtGnYLYUz6QuDGeDH0rMymNLM/QkTudkKS89CRLXg7HDkfNzNv9pMRgC2hxf7Zu486Sn/Q0
RKFDsNK83fJK74w3NC9CjwY9CXk4cLK3/je0jrouvFGp+luu5OML0wzx7dVFp6ctuO26yoIbW8Ul
wt8QW4PrJPZ+RPVsgox0t9TbOiadnr/7xCf7GRjCTx5YdcjRO7EqrS2hhcodA+tvjIDsTaBsnYHj
h14nc/YeY9kvE8SGM4C/iq6Ny82CYLOUJbdTXcYwQFQ1xgihgxgdkJ8v98uNRmGvie84YjwVRqJr
cWlG4R6DMuUzwVLz/lNDU/Yo6YNwxu1gCQNaLSdslzWgD9+E1ZEnwG0HwaFZO98OFwtZlo/2C++f
ZDp/bXCkSZp97+DWtDcvLa5oZPRES1cwUXpu5gjhxWlI+FeYNN3KXYk1amTfiBz/o7YnE4VsHYD9
Dq939Ec6BTlkcdmyXJpYscq5sgrXyHS/36aIMgGL1gUg135Ka8cyER5mYfWZn8FALjtszJ7GgHdn
WaY7QhYfpXgLDNmWZtCGWF3ZKJNADjyyxxNfIkvF9QQ0JGuhLNIdk5oqfv6rv1UolyuLfVK6gG8Y
QuE8MKSJ+6AgCt1vO0lFJJE1pdOgzuEz5/0dFN4P7R+ohmV8BOb+z7VTZVC3m2Z9xOlIetODa4/u
72l05gKfg5czZU013T78+qK++ofGyHjChqe44DYDD1YT+J8Paj3Oi42iQlamH9wrD0fCM6zL6zfB
mF+h0Em/E2OKhgyTdPeR/NWm/5OD6EEXs0gPDwakKutdZJqQzu0t8I5P9sT1bNE3UZZzOJYoPhGs
HSoeLkzjl2C9V6v3mk3iKnvZbE5+6oIHE6aTbqqgb81D5a/L8fOdVUPxItx6g6ZEJwz4A9PzNbDw
l/5PrbgJgA9n+4j8ciuFCGgy/BZX289rxKgjLMYgi8qEyW4IiPFOCPBHUiKH9p5IRjncRz5uUU/E
hQjKIYiWNadsixheUDWZPjE+EniOoLxuqv07Y7ultkakxFkl1bDqTJzxKJMpCRcXc3+c8h0eZK7v
Pl1qshIdAByTBaK0osRv6UaXx4tXb0erT0MWRsbQ4tHgHW33nr8IgxBZ+nlaFy0C20NX5QiWVDO2
ToqZc2EFqLyUvFyGJEG9lmiGitNcz1ZjsZVZG7kDE4V4PSYu0BmlBkenS8hqWUJPsVEZZJxeulU5
BmEtrKNmL/HUts4o62Uvto/+9qveRLA/B8RrUsN6IveU26uyMX4eldW0JjmeYihiSd0ngDzSJHrD
lV1q0aYwjo+yef0iAVizHm6ToF5dKOa/hZ7IfbEyYrCWmeG0TxDDRa0zVWzrBt9+haYrIJsVlukx
paLKp6PHjfQpxh0gK6u1+kacFfDv6GOUZ9M+KNYiaaoy1kBWJ3uPV7QjM6RFZ452cGvWidnkJDE6
4PN7TsAyi/3SY8xybJ03zGd/XDNjEtMSFS8yDRpHqONQew7Q/yvan4ttex+iTUyAuYllGwBltQM2
YSTB0SX1rAF81gYKTiZlQNwnf8D925GgR9nGjsK+oNhbiD7+LFws8QSOazCL2xe7tiHxmvJGW6Pq
WaJsVPj4ksjoGVS4AlSecs+VoNE/0GOK14sdwJmMAaAdl1ZQahI3BjJvFPOBbW7aAAMLIMePFkOL
oZ1ddTiUmmduFIZWgsa+h1QlJQnAEPibbkNWlSXGooOoskDjQ7rQoMaF7cDtnVnxWVof5VmQfUxn
Dc3fdFtjeQUHrU/IaRoMkZmvPiv1n3eQvreGdmZ6JYl7PRK06ZcSVfa+JXh153xIEivhMgrE5aYX
+2lvA9cH0hkSBH6sAJEhAL/B+q5ApyLk859cYvmHeu9gBiEiRYr6u2lEIL+/hvJ+XyjQw+nIQRr9
J9YjH8/+lc2u5yS30da8SwMpQYgNAsIw7yVCvJUWBWkYuK1Vg5fW9tnz2LvcfKV2l7Rc/7bQIYzl
BHAP4cRn/KDEfrfdZdPZQemqQN4DEAjjkpuJ/JnK9lv3rteJboG0VZf3SMYNPZWOfDdBW/g7I8Rk
MgKMAEpjOtUdGDcFWd/wGD/aGX6yY35kxO/zguPEV/U+sC8XD7NX45jaNbKOHxUBqdNS61Lmcq3w
2HVVYr68krzTWn1eJfpGnkkd6a8lXmos/cY7nBNBuqGGfmcuPT81Y7lgr4lN9tWVBu5T9xMLXsTh
SdbKnVQIhdmkwm0AalpQ4BGX67WsWDPe9ynVRng3bhDgLs+n922+qnpuj+jNmvu+Diaz8wFSJD72
Rz8SWssowMPcRoEikHkj5sWG2DSBhYsEvULo2aZafdg76hS2fNZXWjONLiswAo4mEbznUPUPc79Z
jdQqpqZeSdirEfobC6rkR9gYlGRMzfiqCICfw/EjDr1W8lN2lOdeb5J+FN5pOV4qXIdyovIiEYQB
fh3T4Q7wSadIw++vfDXiTQybMAZTLglWPrPkiMBedKshigqVmBJAQGoyONPQQMExmtGUcJnExIUF
qzfqCPAuY3aOu1jsd0fXkjM9o9LCKLnh7kMcZuPwqBGayyNur22cRgnyydRiBcBOq2dc8VJ4FVpJ
gqFCKq/7apTRLeANfTaWBlN430WheoWGpYbX2x/L7mlUu5JQ05Qhvt2htiMHfwlys61nN/gG9W4k
MgOrpTjsEMgc6nLeQ0ZaL7Xk7zf6lHGMtFsVRNH6wOA1G8/uxVZ/znSOblDuFXSQ8yOfV7q1tRmq
wvyB7tIwnU2HVLHiLiZ2gGGxKNP/GgqW5TsqMIJpRoiZBY8jkz65QLRq17wVZ1uQ8ogXYbQk+icq
3dEkfM5eY0i6n44H0YbgpshI1MTpP1M8VyDa111tFBXCwfNoLujy/CxOpEkJSrShnH+8CFeVfB5O
ZQ5CqQ+bguzftZLkme6DF1uFcFqpNe/yd2Yz207vT8qgVdvMeteV1zCjQU2+zYr4fdoCU+q3yEeh
gO4J1/stikPqpx8hJgbKTu03gnDtqjmaR0PIf3d2ar048unjHOKnKERLOV5iC62zHdS7NyZJF8Qq
vkaKrRaKlgarzQocw9jPBHouTy8qkkmzoinF8fm9H2L5PnD7pu9IyGGp/53a5qalIxmTR96FLjfn
VV10aAYPY18/bwON/S1BO8stclLDPGcaJVU5Kwff6zgZJn1trQh1h+ABeBwpU37wQ6qLvU99wIl5
nbOYgcSjw6pgCC6dtfrM41F1698PfmyrA4dX5o6PmoDVdvq9LB5WqQ4Wufy1gfH5GAzhnTWdxbvV
eiZD1km88n0HHTjcrPJacH7itJnh0ALd0Z8JmJH2eX86e72D1mT7GOpQHStAHYfEjwUWYOl9m+wQ
vXTZJwuIxXaPS5T/oTy7kgTnZFk4isUJjgdX9m6NlYapTQT74SbD1YRXCxvXMnyyCvOapwDzjxU8
C40V/BPfOAZ53t8AM9rXNFwt4fUFc+PCIZQ+UP7ollCSwYip05DIEzegHXEFmYBrj0FPMHOYO8xy
gI0wqhAPO/TAC5h69wTBqPmB0SB3eUKxA83no26fWCTAQ3AIxvXIyCZmxiZorFDose7pgaLeHDiA
ce2bG200xN/69Z7RgXwsZi2OWRqKSJwyj9hiYmHfBnaZaUBDyKitkQBgsZbmjpNgp3D/mUgnmOdQ
8kssgcjHFwhlln1xNs77fZGumS7vLzxWnHD5EGS7Cl66JkRg9uYmvFHVNUxOs1e5OFrNj2f2VzNn
vWDftua+2V2cOS8q0L8yqBvMfIbvdLFZ4Tb1RWV16E41/dgruNF66OtdDbhzB1YE4r8twD/syihq
6h1bFeYR+KCfXa0330XlZ9twGdVc/n6KMP1QimAXAAz8FSaB7kRuhdeqBVtpFjXy740Z6YLFf1KS
H4eqJ2As62+6TS85xVZoOr/R+Qrr7j31Pnib5GuFGgQqfBOO9HVInYZlEagqSYujHpzzDStni0wh
i0DQOcczMRjACQL8U+zeLE5BvYahn59su4IDCMkeSVpdJSFP4GKpC0w5KSri3Dsx1xQyXroozXaW
0bno6bFCyqkHjLl07/dZFaUKNUZJMilxCIKauH1KmksgLEKnOQ8NVO1kPS19vCCNfRVBSpAVY0kW
9KcqiWgEyjAT9b1FnaZpHNcN7et3H++Q9+ctPVkraioZwnBliVI+7/NXSvcQ/saNbK5NbW8sYb0g
xhXXHZ8Y9EWApfYkXRDHF3/4hTF+vGal+gGPKQFx3PBXzXeA4pHRVV+sZhfn/snnw5BMd/Vnv9qC
RgSw20d0c3fQC4IaJBV6cAiBokwKuFmk+X4rREvhXhvRJ9TMjbzW4uXrt18T+FiYQ0oRRnCz0OhB
Gqij7uxg0N50Bv5ZNrtXd3tL+/aOVw5UUUTeW5Ky0P/QTcoxBL6ldY/34PRIjPAYpyMM6WQgeWpq
UJWu79prqiMGiIrUd16ntnZDep8z5EwOg3Z3RZjh2+XeUN5NGbDuyGHJFvF81d55hGuuIuopuQj+
Ma5WEq5CAj+Hrun+XcVQ7DBK8bwh92DQ1i67huDHVrHtRofwZt6WGALDbXPWFbwUPWKS+l0HrRVR
5RwUIfI9iaAgdQJ0qysjEtpghA0WDf5WytLuFaaXnjYpooseLBXGr98sTL1DHvyDbI56ZU75e4rZ
+OS/pdWLn+wbH4oeVuHiAlwBD4fDEjhKOZhxLiZf5lD+MzWCWOSTEWaJ/EmlIcd2ydRpa01oiiuB
g47kd5S8/TBf4vJsm2GHBqIyePo+9CSuKo+tSasu75U46hDjHKC3BF+xvmOa9b+wi5KKMXCN4re/
xykqoUp3HFKdBEMjAh3OkcXXD9C44D7vJ2GYl1+FxifRsJ4oFzJDzaVV1WA20YauA8sWwzLs0oSJ
jCLepJMAZlxLX2O/k8ZbgpKGRT7DD6ykP5HG/P6Sfuq2Ydgd2PqmubanHaEbzc2qbHkhkenRa/f7
D0DaaZ11+RuoydsYmzYTZBGZ20QMt2dYUuYRBrrbfVg1jogQ/hAmzCOAkx7Kc8MRJq5IPTEn2fJ1
j/L8MQWW4/fDxZU8KXtrtMmt4zawT/NrXRFkDkYdWIuG++bAl7VCP7uRVlYrP3tFXDSCL71mcBjd
YcOgsio1rYLN0KjfszjFkFq8wdKVpWDrIviszgrt00nOz6lyYDvjcOJEyuWNmuL7CzXoln8odk57
pL08I0oMZ6brb9TpSJyd/0m5FakmaR7TCXX6SiFgN4rr4m/MZVnVAqVnHzQrUjm7R9q1Z3DHH0xz
V7y0Ow33HFGGN2VvUd0Prn9jmKT8KN2zQA1eOWBloJLholmpZCcIyNWmIJpm5M6tzG6u8p04n6mA
eFFTCtd6M24ZHLOZzjA60k2ETXEemPo+HvVFRR/0RYMAWpIrJXtOVWn9iprq56P6D7rXewTQs0CY
P+ah926txnE+6YxuKUDeMrsF00HFqxemrbQ/9J5zfcBhBp1+PiGufbR0mOfXs8qIwixl+l2Pr+rg
M8zy29gqkpUzQNZC73QJVXlwrVje8AijaC/2Cm95K8W8jFvtP3NE5NwJ1vDnGN3w66O1xJnNbCXe
MLy1owsHGj0EZQgdU90k6HbyR0TzndkP/y51MC7dpTDPjStFxRPDY0lQmLDUSKb1CjRRsyi8nhhg
vJKp6QG7n8pBh3FMQ/NqmFjBG9U6evVdPNt8aVXuJRULbdQpINOvy1Yg0BzSyiEU3ByHS9LYSrIN
ULwm8lOxTpx4QleCNC0yS5IIu2UoQ81e9tmtz9HV/y+k2x2A5TcLlTjQcj0ENg/h4Di7EzKwBDzD
714uITuXULKhhDqbMGFiVV8oXSg/jDkKqD2veTSwsZBR+e7+cjB9qPDO/xP3tl99uyv2K999JRhb
NBwzY4Gw/AWEIJCuX/N3tK69IAKSmC+z7QUidQS9raSRnev146SI5mb3cW9IozHuHsfrNrLgtEah
EXhBkRsEiplG7+zorB1Qw6RSADzK1D5D7xNaqc/vMODnnsibDuBLQHvIcGpdyWCyE2W2UdVcaD1s
mSj835PoEUYnq9t8RgJ049F+T/oh3DXaJGuG2kNc0baKN5Cff9ZHX1SS7v+jN3joqEI6lEYuBI81
wmIqFd9tYbyB5qjr9LTtIzVjTKG4bAfGjf0nwkjrpOxuxHlrxoyNPBpUWToPSCZoHv8wXJ3oAjLV
trlfAIpAmDSIzWCQEbUbOdy380nCM/jBC2lrYpLi0zFeKsEAG8PEceoKTfJDvldETMtSkwSTVHJm
QPfKml9KVO8BoK8mb1CtVNohVo8PsP6m5kMTX3H/DK273q+KDacHRNh/wEqTm78xHf4iArwHzAN8
ruE37geKAO6Mmjr7TzQW2sIIstVTGwKLqBonhI49Wd+ExphBsmMgiu3zWU3Lduz0uDnWLOBBcBbX
iSbjRm1+OoQNreoURmOnLESHwDCAZr9isfKBga5131edg0aCjROdsztPycZmE6dcZU45Q4T0TYFr
Gl/OwBiOiQdU+OFDV+D3zEQm6GikvFBTlYxCtvrPHsTnv3fRvsSQ/3FPuSOaXNrUOz6GN1PJzGe4
m8HSg61d54dNcTP5hmUDsbTeiIyrBFn1deKN7B6kvGQtCbVV7wiaxzsJbIj6oJ0Tw+pGTE27o1By
pose8rbVB14jNpRcf/VFq1NZwVR5Va7IkFFjCO6fQnB82xlrWaJGLLvun6Hq+Jcveq1jZzGZgS3r
t3RoJC239I/eArOO3u3ppq9BtT38XGb64bF0VlO20qlZyt1kFmZIp3HiY1YupZNe0PofROGGRTNw
KN40rbVNGzssE9Nk7YDjqACc/WZ2ItEvUg8dVUbRMRRERoedN6z7lu3xP8TZEzJFKHDhDgkiGkht
7uEVBqjPU2wNTOBgObCHqHKwVCaVczTkdu6hv1PqPRD/BxW2dASbXZlic3vvfWg6zpMgjk4LOYDw
JaT87ggLZC/wS0/r6QhslV27ZMxzCBITKa6ptJMZ9opwaXCSz/TjcAP3AOVFf42ej009qTDHvgtF
m41TbM6d/cO4KayxDh6OJ7RkGrhQipQlS0Zbl6b/O7uBr/8rzXlsvEUUoldf013NlUIDwLEtIa3q
JszyateqXbAMVpwuYf2LAeZjCPbamgBrBiaOuzYtk6z5n1KYhXWXycCc2LV0VRoABl5uhMTSGwLx
LR3uO64GFrHaRjVlEDasAqigx6xjUJzeaxzVXKp41F1tJndKVLaD/t9wdQCfrpzqG7TVfoks6N4Z
UCXJsjh4X6qJJfx0EE9bKH6+7/5UAE8cmFGZFvoBHFkievm4ILt6O+qwWjkE+BSp1RVBkYUO6TZ0
Tx0rCALuvRvX9A3L+f/7K/10tLuPufkcCbX0BTKgWYvFBw4cZzdISH5QHqHtulPvaZYPMNHqQekk
FLdrQR17GyzyHc2Leyj5JnbcU/axMXrNz3THDKkqoljxR7YbFcP90i4lyJGd4TT63Ihejp7rbveI
MBEgkgFsLEf6NE1UA2p+e++H5oFEf/XUG11fAE/kiHzZwLNB7MEMbk5yI5veB+CHKc/ZvlRYUAtF
JCAyC6OxKrHfVD8RLFPwQfjUSqnJNLOXY9hWFUTXNypCTnVnxxlhGiJMV7Zimm9sxI1hee+BPR7C
jq6H5Q3+q4rf/WVpcVrps4a3koT29i/TW96YfXyUasAqfcVIEhsZt5cP5366eG7NurFwaH4BngG+
MxaojhglHC7FH8D9U1NJRyQQjtkAik5KqkbtOAOiHFX3KMuJTw1ptxOVY3Ge09wARVMspaHgU4d1
4UGP/Kf/X4eiFKOpCrQwGGIdQjkLL2R4XWOXOQQWCIfn+nAweRE6vJx8AUkGZVxRVjoE1V1sOP9P
50O32A7PlGnKVR7qeDGlMVkm+fsUhnL8ql+JJCPn9IyLq2aYgWHvKFIwRKW9s4uzWlVcf0XirirC
Nzi/A8XUA7bJ98s8XJ0TCNZxx3rBZwqJQpX4Ip1WvY2pFPRnD4FQVfsjCG0wpxUKo8luhPuWYyrh
jkUESuVenzLM9w93rzM9+VB7Y527tqFVXjPOpDLjGg3cifvisITPmyRNj4dKbk92sEKDiiaS/Qc6
Rgbc3SbdhBc/lDV1LA1qgfR5T4xOzYDKhtMvVmk5FHqurbKgS+XEzFkTvCxhWvMD76cf3pAAptoK
Uqj+K7/TEFnfYBxSTFQm122+SL12Bs1b7cu3S7GTYaBxh6jXgKwUiggrkwByhvP995QcVKeFiaOr
6IP+CDCj1cFZAXVzitHAlK7YbIfKoz1Hiw9KiGRsyhijThCCUSX5O07S94kCcC7SreRegERIF0KF
pSW3O3rDEoAlBHPfAlSePG8R8RGZzi7e5m3vcmZE+qzOP0K6GL3uu14XgIkRy63kmRVFA7gK//CA
8whOENSFftkLqNSMLsaz0NitIG2DMbUa0QRtvcmaeiZMcG6z12+ePEkIjj6D7GiJ9/zx59ZWM2RQ
npXAsK0hzR8PYVT4TZCdPIUo9qdNqIQ3DK4owK+/SBdGgaXfcCWzk0tSDcsHC6q+L2C9qJCAUlCM
x6gZkb6ntvwJ6vJAKzdVg2uX4JRZDmimnTIWXsRyGbR2eS1oRQ/aFZnI0CGgvt73oHtON/XGFrV5
f2UR8AdMa2C0nC1U3ctjc5EKKi864jDTOpTmzE9EM1FstE9LOkXHbSxiTz8qGQ3yDrcuNF6svHZT
XkSGo3RjRhZbyMDU8btE0cHmqz/OZhA3qZ/vXjkxHXeA4rW2U5WnGK8KjJnKNrw1zFtDje2GxSyJ
VKE2ycHhCHHHNSKmNI/Daf5VduujpvdKZNBBiXUK4RpGZRcaP32kG4J5nH/lXCKXvoLOW2bTgii1
V6GuVP0oN0kymTuKnH7Jo/Vgj06uOoIFR5Do730nhs6uSJLiwfnXhp3FHpQFkvn7Rq96SbtYn7Fc
YUylh2Ioxdc3S/6AHSEBq7n42XfaEiwdEU+7DhVPxzguVovQoU7SKyz0Fq0Q2DlQTtBZVGG9oU7l
DVVninlH3DW8PLSJByj0XIMxeX0QiMKQvhYxbIJtJT7Ij33kuGFOiTYb74eC6HGQvxQkBXk5y/Yd
IurFDy60TnTWFZvJ8PW6SGqIa6rIlyzR6WLQRgulWKAgswbPm1j8cw++qxvKniNAdY7tfQTAhORA
E2vucpj/edpWQnhTgK9R/HtQXtYZsWsbgaQQqSpJWYyOJ3MgoZkWDz7+3wMR7N+jYtScw8dzyEiE
6470kxpPC55y9j4cmS7AVC9mjRs9blgteqowEpWonwerydJAs+wSeDZ11ZfkSqhU+ZWAHkmrGBSv
HdXyNAuQ/CbAj8YtAr8Kr1olxShMjSAH50/RMqEsNWFDDI5pcT8bnLaMCkIxNGYzFyJSYgCv9DKI
UmHM7WdSkhlriEQENyuHHWGQw0skuw5EOOTbO4tgp09y5Qq/iEuPDRUspDzZQHs2reqcIcfrBJkP
aJ0IG10W8QSCb34zs6k/WFZ12bnQBK+Hf6V1pXsDMqOFFXfZATPGQ8jeXxYpzbA6Qrnmcvt/mhDX
iAtZhVJqza7fawpXi7mXCi0zyMHx9aY3i1wxSkhM3OCRPEk3pVQysQ+Tu+CnuaiAma59Rh8leMHV
3zd/X/27EU+q9ct2DSl8E2rBMN3/BY3XStak1KImCBfcG/En6Xpa/kom2jCBTUz/Q4C9eUvIJQ8R
vUUBAwNiMClsJbeyAs7J+0FOLFOJLQ7EIKO33w5SigKMkqgFVhXGsbimj8uzQoEE4gX4Jt1se7jL
xb7PlF6BC30K27xcjAj6/4wGy7fKIIspFeXFijMSFpIjBmwxYMoTu6Yhik37NQp24MmadBHp9p6D
y78wt1tDVKFRek/Nl5qvFgaOEpZaPCBAkJnahvKas8viyZQYgnTAJ8J1G5rJhEd/VO5S1el1t0Mx
fEB7a94wA0yAzpUMSNb19G8UVZm7O3qR3vrCVYD75pS/VAPbpBZEndMPcKY75RFswvXofGM1X5lD
5ikJSVyegxL9cA1F7ZIoGOCfPGdRWdQb15ZRBtYJvs6eyIzxH5wyDYrlTC8q2VP4hsgcc0iAIYA3
bznbjBaI5jUrnBaUI3mUliqhqqYHgeSsxzC2a4cgoBtpkOrUw1tA3/cxWBupzbbco9I1i1m0X57S
NknGzhYH0FnWP128F+sW+n9c0CVxVO/wGGsJTFyR2Q0vVYwqA2BYSpvUfO6VdE1cR0TnSOKi3mLZ
WS74Q1uq72bAR1fHzuTEkgqVz3ZYxrgvxx/Ep1wjY9gs2i5B3hyhbHDjMf7KXOn6m4btHGmoiF9P
Mj3xIxpL5EyD4Phad/jcl+1uoFqf7TPzwkULtGf/zx65rqc9fOyBfyHxVFCkpBZqQolOyS9Jpo5l
8YKnCjDOL39vOW7oVSCMTZqyf3eRttkMP7WPDxHttHOs+7dK/fQafezQn3Ati5wbfWMP8pgT77yG
XEVxOR9ipDwL5FAaMoVxH34aa5ksavijIas6nVYCo8FJ/f9HWXyylGTpsq7V8BT2rXHqA2YWY/oQ
CvY9PPPDD6la5NtVcgEtafSEWaAuszOVsMmkZ7u8q9P9XY6bUPdQ2QZvU0c/iiZOQeqc2XMOLtoU
HcjsTMpMiYr0ApQ1UOBcyvmAGgj7fF6RlWzPzRoa1KvPDSMjugyrvg5Kc+LpevXKyIlAMzktO7D7
bcxre66C6Cbi4QqzS6AWk2heyOgEPCiCNvuPL1vtaLY5FpepHgI9xhC35W2Pp9Q1cyUe4r38NMrz
NNVYPuBi59p0aymaw+MPRgDmtXJ07nAEcA2hKekXeK5h8CLWMCvBA+maOVbqovUraYKQKD6CFZK/
9r7NT5iG7+ynHd31Fke1B3FVdDz9Jp3WDXl2y3v3pryCQmUOc2npdQ0D3kqXHX4b176tj3LiWrS1
hBYBBED7xEDgKBEzk22oZG9jtf/lYTTL+g6GMb61PMPYv7kuCDTRKERzTuCRZnWw+bmxUqs5KwjA
7cEWxYnUSt7EUnfV8acArn0ssk5kkaZ9LGszg8ZiCjVZnmi6ppvobJV2QVg+2HtmcRlArnFDlGjg
sCjYVlfmtoyljI9nZ6OeI1Dj2paGeOMRNhGuinWGlz0ysg7d7zf/yunsmJIujl4ydwtk0Z6vu/TM
A+7FW8G+/GwXxofu4EVBV42uQz3wEoA5z2xgyVYT7/kRw8Hs0BanxXPZDmxgIb++vl2Rql/jkXGk
JaFOSTv6koniWlLi8QEXfwq0bshzNXLLHc9VIULwnQZ99K9zYb1TX6TLXkODsNW1rzBdyAlGb9E7
i0/vOg0s7yxkX6/QWn9P2fKtIIb30Iyrx491icSU3aHjGiFFc+LpRLvKRo9WR5Ex8ePZDvJ3CB27
4g9cdKEA8FMjr6XCXi30xD6fs0rr1MbQZ/57rOPQkYx10oRqKsHUz8TRqhddwdoBj70CLDADF6Fq
+/y/rnLM60CPMs4X0OUk2mmQ/Ax0WBHmt/21vpifFKXcg0w4FonTWNnM0TsgU5jc9VxeUMgh1cid
edQg2a36T9d6JRydZZitK2a9nB2AqD3HFCqnG3Iyx05dFDGjP55lP/b4fbouT3x8+smN55YSR+Io
+cOYhIkSqdt6s20sWhbGNPx2bZqyKwtP5PyLMvFoDwgJFDhOZ6oc4c+6QBsvHTxj9xWoVTviqVcR
pudvxIY4R0U/ElbNDsh92NcW3XH4ikvzQEXI92nPlFxz/fF5mkKKjhGK1moNK8Nlmb8qVgIG4/S4
wX98l5Y+nRHo0UmXWFTfjolPqL4I3Nair9JUMDyPW6OojXeJWgH2kUclVZYYtfWsrgdNCo+utvQu
WCBre7CkOXAax0L7V+j8qQ+9/nSiFlLuzMRSYjF+DZgMg3MduftOogSdlV1CfszZUZDhVdmax9Oj
1uM8TpuLPCL1QISRtNtjwimmYcVok+2oKrTvwC23U9tKQSCoHJQQQV8U2sgaCEYMgxd7HxSnqzbz
CNjlktZ+7Gdm70xmemr77MD/45SIR+yt1dMCYGBaC1hWO7T6/06njS/6/HQAMQ+tEZ+RaA++noYV
YwJhnFKsBzy7C3ZGQUSbFe7S1EamNeIY0mrcKy9UOZ0KvLPFezO7tdqnBLLDn9XsIDtofJR7eWcp
z+Hkxl5YByLmzGadY8EWqxbOXvZwHkI9W25Hyp17bpoCzzVPl/tUplYyRHEw5TA/XhKY0zSiyXM0
GZdez5jXDDva8hpRUH2md3NxAyqLYKuM8cAAOPo8nOu64NbIRO4MgoQ1dZktjVfDA8hXatZ/katk
eEzN38cvF9Bihap3ml8y3lt//zMStw/Q2GhktbWLmyYxALG2/a8BSpw+4Q3exF2SAfHTIkVbcxKM
sh/si6qbEYCu+7qrF8URQz1E4603mstJphzcmF47i0uI7UBqH9QsJLc41ySD52kUgbbib+JiM3n0
wZ65Zlaf5ThNpkHDuC69mEIs3OoY2Y4obb9yTjSC+W8t41qstSW6o7ph7JzBl6i0F3XXKxJnSMf7
YjhG2nOMT4NgPZdsqC3mogkAg0TYV+b86qNlxKUoX8e8/X8kqbYq8X7TDhTWYNoiUreJAGt2ntqL
pE+6974uRZELSOkreZF5GAMU74ZdPK8jN1wKISkg5nzgi+s3seDf5fjbDtVXe20RV+QxOPASGeV0
vJUcDZkXXIn7aXAN+QXLvWYwEve93QtkmuMtPx/fycwIDVLZZn0Y2OWJaaq6PmbMLtaN6yfzjYZ0
fEw0xqGps8bRkglLjLqYKDDrLnfrIV3eN8GPXdh1KnEYq6WXJUNTCCxTB2nT4Sj5+GS9bSv7Vn5D
+tPwCi67OHbJHjxrfZCGM3TmUqfWIhd0/Vt6AevGQoCEBdvoY0KODn26yhQWwBhBLzKpBEdoRBgY
s0AjYaMf9WcHtL+//0o00KZBuf0KONi0eoc1fXBm0UNsJ6dFsbimWMhhdgXdOdnDRjlKAfkXPFk4
ALK58E3nbj9mfOFLYk9VQrEQZVTkw583X/aLnp0WWkS6bDWr7o595633110HlJjd1ohevyTpwZ5Z
lyrY9dEJEWKBu7yfkXUw1QuLNM+Nv+JETr9a06sKPcpC/f6a0X/oPZd0r1E3ByRzGmOHrL5+N5jX
5AxE6gXcf1lv8Kc4Hpo9QtXXfXQktSXW8BkjFHU7bD2/vbNEkEM21yo2/NrPmYO5xfJSM6LNTBp2
/nQ9xSUc7C2bpOrFvSGJo8hsjysWl5AT5oZesQ4R4N5n3D/hkVJO+W86z2Syk7MTJzU0ku0oCqWW
c2kfttl0dgI3ZqPUQR6V3hNszOYLATIf5d6GHM4SGnUWz0fvnqVmGaTffO8D+CYgxHNnpiv5oBPN
nvaa26fhQcdS15V7//RXUUjcRslu1P/+kYiah/ae0LfwEh1pnMuAVZg4eT5ftB+HITstto57dYsQ
ufKCyBRWS1nI68PfTmG93LsAcaXzCq9/YAdpubFlERfz1JCXw8ftfq9D2WpzompmuERR3yKYB/r/
AfEVyHAfX+OHoYa04HAQIjGp/X3Vva/80eGMhICS5zCN+dcjG9Xb5zA7rbYmlI9+jCAFWF0AksCU
OodEntr2ZtcQQSsDco2bIkG4c4Oc4PslkEWx16ScvL9+EWfqrquSVYaHmwKYGUACDzm3j78JIn37
A2nTwE0pwaA1bJ6T7HgLye57EV73m69VCnnfYLk5MIhuZ/fLaxDBUZy7ShOF9uyGUwd1qOSWPK0U
j1ng7fYpX75OrgD4cTEk7TX+tuF6GS3vQ1IwD5fJ7fEfB6TA1tRVxHNxYf8gFSChk2ecWS3hI0Jt
VW9RhaJz+oPS94R5XbqJQMmZlfCpOUTqDE0rMmz6iLUlzxKmls7TjPPD1x0OLuzvZCOEFmM/2gzC
SfuctkIB8qWu6lyOmXsqLePe+on8iuNIcDY+9X4QDqbQPuS+TwmIZ5vCXJHoRmax7h2h3v1dEI5d
sICfsd053zIAuLz01UXoitcJ1AfCL6uBBBJ3lg5PFHFa+zVs8VnH5arNk9ESw+JPQ6s7WeRNl1TA
aN1CBCtmb2JJ+5cM2MMcxJEZCUVYLViedP+bU39TajooAaYmRNbjMs2kNL3w1hOZP3npR9tGsdWX
4D7g4kSSaD7Gp39lOj7/TgxwLlY7Wdp9/vK15zmYWeIWcS9QRjiBr+odV+yZYUYtw/2A7X8S3WKv
ElvaxNFG3Qo1fKNpOaU2HGGW0ETEtHHJ/eeQJXmdjFzrfp1EtgMscrPqIKdLaEhKF04N7wF14eDS
jb5vFY2Qgb1rTuzz4zcEP/LYjHIbJUB8qL8eVGz8LwEeURzD8AMTXjxsSK1k1plsB91zLl85HlQ1
WLYdsueUHNkFWQwnfqxLwcnryWkZBEbWDjqVRTXIPDnb7NdBc2Ky3FZsRJQu7z+tIRC9K5tjf8JT
fnVq9KI5IuBQ/1LI/3Gv2SnzDmpfDolVRv8N/VKqqPh1hg5pb+yQWoSP94ErannbcFjy6s4o2H+c
cJATjvVB/svPNaPN8f3vwfnTgA7NZeTS8czFKJ0aA/ds0IRvIsKoKkZt3dsatj2dTQWq0++Lo0C+
rK7IHfgcoZuyKz/OHLrV65NBTC8OB4/AyHVrQu0H30sSzVuaLpwvDXATidX99ELMLmaEnTQD6wFI
0JOS7KVkQ+IGNOzKogrm5/d+xUDTWqLIB6dSxeZ0m0LrEiWpNdkWXfSqn2+g6b6Ilfyma2rF3HSt
Cy9tpWpbo971IADlXjKuNuF8kSd20MALJwofYokuiQGwKzJukBpFyMqh5YwNv3d/NbnWLo7MnNWT
Yx1jfYtFfwzd/PRKW0xAAZUtxQ+lhNq81OITFvAXrNGWlCnmanOEdCbAE97GCJXQwRXAjIIzJGNI
U4k3PA1zi8rjt+g5andscQcrgTYwFgWYgoNES4RYVPL9KaRJS65lZCN671kH9z2nEQ29dQKFs62p
zY8ybxewIMfoK7Bd8UyleZJ1z/OO2jG+jCbGs/KUdCae68wlr8ZPRkjg51Rd9/73EKNuw4qbV0at
zWKqWeF1WJUJD4yQIkL0NDK1a5ekVSVmjUz6ZHAPYbHuM4cpjUi2SxXVzVDOTH/h7K561ISzx0Kp
FtBIVlfIQOUF2X+5FlvBmSxA7X9/Inl0HqOPtD9XsjrP0vva2VZHG/gq32blo+vB4rFN/qMF0a31
DpDmF8iTxpQBCZo3baCXbC0NlTr5v6d8OW6dIg87oxvxkAbKHRfDfvEXQHpm3LAU350dIPAYpiOv
NTBQgrCf6G+4uBYL214mhqJAqOc+sV0ruNtmkbiwusIb6NarGwY1zH0omYAzg+pRA2O5W01Y6rEi
AcCVIfGUzMMztprsMy+PN19h2MdlsEefKnYEm0bit8rB8C60fWbUIjwvXU+Y/lTB4CoBfIy+kL9Z
N6pq8x7PpJnDcS6c7A1/iGf9h+RmakQY9XxLoegMkEdyDw9Cb3IIhUc52OgwAxDZl921lr+clxl0
olHgM9Hib3N5gStMIRdiN7j9MQk/0Dma4rBKELtkVEYDIVkR/VHzyapjer6YuiAlQrgO5P4A9rV8
3G5jFlymJSZjwi7wXfXtM7O0ylyFwPRXZUcZybq9Fs9boo8236TEAruR50yAzXx6rVGy8kA5BF7o
RUZWl+0OuWiSOG8G3D0YSASkehaj5U5atCiC/9tr/riFErkFwCtniJKaRpJ1wAe/HjsecL18NBAt
ttrMd/fUKDHk7/AmQ8UthkSPRCDmuXHU+5NdvmzGh8Tel+jDyYkwO9Eb6y2/4ZsL2Gfvcv+5112b
Xsgjc2+Uai7wzo79hDH36w7u5xVCPHEUK7keuvFbCo8ETY5QhJ1S2YbSeysLo4ypyV6H2EMrR8AQ
aRzxRAkx7O8K4O/s6ZY6oITFmvn4N+S+c//DkM3rIs8isiZkyWYilVBi+qxffUBBWA/bMpB+M4nY
J+6swq/12ClA42ZIabzncpo7Zim0KjMUWSQFViOIGN9D/WRJi8SaEoIdBc/ws70cw9lefLyrbYtz
rRV5Hk2G32Y4Ur4mZOeZ4vMrC8OFNDi8Io3jCwI////6eAGbdqJrtQlLjMC3sog4mTUbs8DtTH0O
GiywYB6LAASD5W6UpxOt/V7KNTJjJ6rt6r6WjmJ9YC+KJ9hYGxeT57tNnTh+LDy87t5Gx330OjhT
sFYxJnsGpW2RYoUZ5cC7yEc3Tk0PXkwMKB9l4yDM1lLpQhLdxGnXMWMtI0W2a8R1STBJze0ArXd4
ajosQ7OctVorKcxar8jlOerNwjQ0IFtukTJJ7MqWAAUH6Z57xSKWGYlJ1+lCUt7fNAo0zm1HUmAx
l5rRQCao6lU+vpQFJcoJQ/LE9IYJAkWqu6SPNvRtjKzbMlWFCD0Co1pYGhmERDpUD025o5hyXcEf
pBqaOnD4Tai6cE6Tsrlm1UDWOIbS54RcLf9YEZVDIKrVuLFBRR6ccnySeYmAf7JGa5X3zImdjhK3
+bwVzPaOATEdFf3Hcl/mJeU6dKHwOzETAgK5aXUsATdNd4ADIoqau9axx85I/yhigjRc7GAXYqyo
Jr+tc10yTWbflBJuPYTDaogAdBpNZVahqbDxPV4mnpIR7kWUuv4SGDFpOc4TlxGUV+BOFpLMXruK
gnx8CRWlLjVbjW/mZb/28Xq7RC6lk64/GWp/iYgsY+n5ajeLh6agp/JCrIH8/F2phdQIhTUR4O65
/e0FH3mV9IBTf3y08EAJlz2A4JYQYBwGLx1kfms1LQJYe7nwZ7JedQhksQofRE7RP7dLbcyQhQ15
L1FiRyAXe1CY48toCVft78/bk+R4vI4zcmzY09+SgdIt7r/sPi6I5HWKODo7xteJJ6Gc6pTUzSUO
kjIeu23ITaopQRPI05WyMR7G20R4zyC5NfFIh4RkDQ04qK6N/rXAlBFB8+uWXk2+olpOmP2AYo8z
KeyajPRlgduaC1uxZoBHVjkVutUQrxuQALpVxAh5ckCAG6LFzIIz2iLDxe3+7WKyXqmFD9z62N+I
MiKFthuKpf2Q5WM8KWKRbo0X8gDMo5rI/g4Y1n3/0wi5zBW+MAnyMovy4rj3KbLhgzdthNJnJKTX
W5nFWSHIlLlV/9LZPDG/J2t2kMP2J4n9GIU2ixdRUpyRVtRWg7a34XEcfpQGSB7Z71t4s29fHpAx
1oFQKDwoNNCospPi2W7ljfTi6x4l8z71cu9bJzJ5HkQq+CKQ6JXH7dyLUx/svQk2SJP/mCWhSUHS
vM5GdqrA/g6CyeG0x/6t3OCQIFoRhuP+ZGxRZOZ8piwU0jH8iB3q9kWptd2A9VzEzVPEQN/OEDG7
LQ1gUCo/qnwNePodWVGKsSUU3XMejFxaMc5txqOz5JDWDDSMwenhp3m2TPumcJ0Fhgilxc8Jaxk7
kiJbplnr6PVtzVWbmtHbNuozR+f6YMryJ9FmQUaRp/BtQFQJWnfq6fpYM1mltlLnVPxjPWRBKvWP
TRGt0uh7D0dpQcrKcQ79OhybCO39hs0je0lf2o5Hc5M9nqwM7cspQOhrNJgOEtf4wRVdegqAsWvk
A77XE3j3EuPoQOf9gvNE1Lnz0Iq43fy5IgFLJTSkGtgtfUs0sruW3GLc5w2B+1mbOE7dsAHJI671
sw4L+godmLBTm7KSpxw90A8ooTaHDiquIuNjPUfk+3Hy4f9resgRLi3/owTicEl0K09FIzdvOfke
QQZ+N7JVzdT0TrErwxXIvbJc0XD8Y4rWCbrwC4KJcxErjogQmJZyqIwoG1bWJ+V6xW2JfTTeGZu5
cvGZz8fvnPuZsXvt7G9iwEBra+robvtWLPEAaxEXFfbCWfSKk3mr5VypiMX3B/dmDm7rYc18bDry
xDWucUfCK6Pil7RwyXwoYr8OCIxJUSGQSjmMFn7gy/dGYhd2egfBUA0cFJ6dwjO5g8kr2CjXQK2R
vb+0WVcTIEfgMJdSGKNz1wZrJl9VW0DCf7I7lpIwka/Cc62CF7Hm4OZUN4xcL2GIso2rTj6/G+wS
lA7wUmSoOvJXruLbF3UUKk3a16tSG5ZbfywsQuYbvJSH3chof+3pXHLNgZ9nMvXT4RAW18bHZyOJ
i5BokEfid2Q5hxSWnJO/XJOVYsFTPAq9w+BCvoUKHkvlLdmD7cW923jaxoEcRef+PuR9t2dWYoUb
8OlRn+zIdWwKJtaxxE5iy4pF31+nNmpnQb/n/GlyOGLOl/Zj8eN3ICNu/qAFwh14GujlTWnb4XmZ
t/UFBxMC2M2YlQ+VctbyyHbY9AV0KRaQW+wKS1n3PYaDycbfpMaQq3qRExTCXjJbUmTW1yUev8RF
cjw/TUS9GOsQGNQmZqon4tAN8TndBdmD1Ytc5L5SoHU2rv4jyIfKa0lVtyZC7h2ABodD4deDsKhw
VZNOQZ8QegEqM04IdBnvB2onRocffIZVqRSI8n0nDoSuSgfuOW8e4aAwEtsCE8P3/uO794p9NMtO
o9RCY68GERSJBerbtaUmG8dnehQrm4YFrlOA39OrBpiisr5Fl3FQSZNM9ttqa8pvgPX0eR4tpN/O
KjdynUCKl17M8YgUrluICc9cEuFH8O2TtCU30z6TXxL533ozZUJxDIZ5XgjWaO7UDAdSuBDf5lx6
lbfaGk2ea7iMKvbJ/p2HeMzHN0tBMpcxaojlL85IB+pgHDAvz0k45IzTWvz8fjtNq5tvLVqPYPs+
TAkb3mjsXbCT3zYzDHUOl4k2A9tC2jxeqey4hrSa0EWg3YyKN9EPykHSvPmfI5u2YkbYE0Ql06DT
mwyeZT1qDcP+0z4PwA9lqQk37EumRDPAG5GlnOJNQ27blyq2xhiZjyzJsxz8BZs07zB2tVmeXqI5
7BXrnU0edcsjcKJui+RpUFhJ4C3lb26qDYv+rXUlEReLFkKrV021Hexrg3ROiYLh6c2Mink6tnnb
ZqmOEjTFHhUeC3Epgqn0Aq4+SX3AkN30gElVX6B5AcRmnzz9onbQ/13/RfDeo/04Dr31FhMmY1Ca
r+yB84N2AC905M68+0icj34i316V8DaoJdG8Q556gg/zHDTHN524I4Okx/OhY2u4lmZB3+dk3Lon
1mkHUtpTrAPlrpOYiSa8UeZhJLAt/7CthMCv9N/JwQ9AX/v+COs0lAKm+Rs5IK/KCQfOa8dnHheX
QfluzbG8WkIhrgReOPjuThMNpBxnhOxozydRwNpdbXrID3QVJ4CQcPhImVJ13mjZLdH2eVrIiy4z
sdat9x1mZe2ZbqUv+S1GmWvEt4H5vrA2Ov/vyEDqJjXZ0+V9CeyCaZUsFe6saQhb4cTvdmahn7ua
s+J03TrKENmB8FeCSOy8v1IL+lTSM1uJGn5CB9Rr15pIgEKT3fvNYRY+V1ZmXydajYRT8M5qtJxu
eYFghgJnjrSSmhJ8D07rzCXVLmJsanI2koEP7hCuLByWAo9b/TmOBNLL+WUHWuIJCOhZ/Z4T643Z
I209h2DAHsmk3RUVLXSJV7/nIEfG3hyFKLCOb3EzkLl8zi9QXqUB/CIWY6fZsTFAw8CBlUh0ykUy
g6arb33ZLrc6Yb2TUzIj5sNI7sE2i1oKxoRpK2Z14CBe737NlQXb4E7F4sLk/uJyZLcAia8L946X
6V+zSv7aF5ZAoy0q7rc2Gmk4LVjtCI2FWDEEujreXuzSdz50S9pBe9Ed9jnd88zoMQy1Go7yqZfe
Fh6p0niIPnBQRI6pwgCz1IVM3OYXOAo4Sidh3OSRg122RaxzxVMfmYtJp4SSkzLXFkiMYEROYgEg
bCVkBRBGrJavQlS4oi4oLqqrL2Gm/+VZHP1+WQKTcKUuUYOLFhzpv1r7b6OAT3pj8gnyDp1H8cA6
VyV+i5CN6a2IGREfrclCBNU9YxAK+mSUp3oM4Io7eoPRpblOv7Wuf7GhHxZtFMGLt83T17tZoPrl
bYTJ/0Xov3zmiEakEeMwNiJh/Um84cJiN+jHxxJmvSs/1wwWSN9HvvWGjGA5JFJvfywkhXhPfAXz
NOmj5IA8BgCBJwoQHXEUkgcnD1qNX/ig6LQ3zuZ7jLAKlL4vCyLHm/x9l2uLFCn9XwGjJn9rq75a
cGsD0D2huIfBT+j/aLjoW9aaUGin24reU5G4auPstqeNNqncCVdSi+GxBJ+7N4croPAFqhY5hXj0
u1P7Smi6NNnk2tobwqtU4uZcL2uU7p4bZ6PPontYHyCFGFL4GItDEcSrTrVDyuhPhvzTDGhkQcwb
GS/MRLMJ1ebyIUogvRF4xbQfBY/umVfTe6IsMburvgV51avOgR9DRUcJc3eo7kORVztEe0tCha50
ldEKcL9BV1KM/AVymihYuFuXOJGJiJpuE8oX9zzt+wue+mDWz0ITHhZSO1Pqlr+RsgNxt2tB4Jh5
s71tfwveekEuxThr5vv9tpUPJ3R4KslkGZzL73WfVYXcRozlXwu2I3cOfryvgJG71IcBP7en4Ji+
ZnOGV/ksYtDV4FNjsYxR7w7YhyU/gzKAh7gUV8aRo7CyE/Q2yaoNS8FbJTIPSBdhB6tq6Ju3GWmj
s6fh2uxZ8HPmZnwk22YLXXqw3wSKi/EqNdRTQXtSDG21njlWkGuA+XB/57a+F+imkPYCw9JGfxk4
80Ru3BxuMhjXV9Z/UBAm4oCU76O38nxX4Jh5LLTs+Rh5Yt30fNyCzhVi5du+XNhIOs+M/VQ+ST2J
oOqmkviOz0ah/9nlXfjsRvAtsCT84qfeWQSHhIkHUatzpfVlPi6o0Jnf8xHY2zEPmtBdgM0zwPoh
I6Y0sD7ENLDDgQB20kV4oXnCMloRD2ctdlWujnc6ImXv/Ko8YfdZI1zp0rgcDYUcDjSCus+nylt0
lnfgAV2eNWdCL+KySUsingErxmK8fkkKPwylU6b0X6WLCnmeokM00AKZdOmmuJtKJ+FCpniuMGZ/
RYEgl9V+by8xRxk3NIKqyKzlpPD3HZY5OlRxvt80sIpSCq5QIqwH0M7IQNbJbpqIDa71OhepKBxN
pS73y2gF62Ovv2/wKqrOYhuQn4fC/DRmh5iTuzywXfDFUz6yQZQDYepMPt6JhJNfsiG5NS/j/zDx
0g4R/pD6auJefiSVS4pvnIuQyYCNRD4ZSQvTaUdqIWMJEpGqT0BuCvO/Y739it0BTFcDUqpBED/D
ReHkoxjEPIHN9aPgnvlenMnTxjR7y2gRBfsqMZwdvXrOo6+s3i80EBvwmgbHFjRppKWl9/FIpwpa
L53Lt7POFt9md/fJ0jbGC9/JB0w4GLRc/6FRfI81omyTVPHuNWzsTGI1UqfOT4YjgKwlwse80qkD
kPj9FhNuIEI+uB0nJeQWpFzsDrXPvO5p3UsbgL0XxLGOqyJ2cGWZyQa2tDYYf4qJAHYvWIVGx4sx
QfYFH4QF/t7kVHCLj9ML26AMM9b0wsq6Lzds55RITH+bW68ahV2vUIqZ7f6atNugGEd3zOQpDK99
EaipgMJ0skCr7OEXlhgSxEilSxDQRogNDyxo7lv0u9yu0ANwF/1cXlREVK7Px9aBiwNICzomPXZT
xiZIAsmPAjE4H6WOGz4KM+1EdbcnS/NgDBGez50C6p7GWMq3gLjvyIIEPlp+CibXPqFST21lqEPd
iCYrY0crrRTKMWHYBNEMk4BO1ISU6O6yhoMqf7r9TSCogTs0ceOQ7OyNEYHvX0RpI3kjR1Jkkjd4
s8NE1DapXipAhgjsWfneErrDcYMYvWPLsnjqqkJE77isGZuI4XsiGgQnwBC9eeiA2btmEIViX/3u
0YFcyOTOyRq+mODRL0Fr+xwB+TTaRGRLzKiUoqsS1bmKDrehf96p1FsDIcN9LvMvC29OiXL4ALMv
U1euVwnwddKOXhSLJ5ChHB2yKaxXLaBvcVyh2jr+Zo5syVW7Lwc71LO1xNfKVUsQ+n63Iqal2Hl5
2mq378zP3C/++ty4jgov5Xga1X9LKnsyMeqAxkfagv5OUz1E4ejYjqP5cm0LpPSNTVcGOJ+dNtiL
tPC4s3KLo3czxut9IiVYENi+128es6PqTgBiVREOwhjBhJznA1nPOKR4WAx/osKDgNErHEggc3GE
3u4I9gXKedPi4CDcm8ZJbh7sxc01JYgGp3PwR/CiFFCAv6ojBKrvb074McxObRu9iI/DVs3qD38s
sTg20J7SqqXkR54PsnbWr53t549UmCKVeMlKD828cht9brinikQD4xXv3wnIeVdSF8zTg4xGJO1e
h4pi2XX1hTvy5Xa4qOO+VGkrWjkPQVL5hQF/t4Nd9TnEziHi/rGWRMjasqGPEMmHnSIh0fDvVpkw
oRLdYIlJSSQJ6EHiVU+qEN/9pPeqHcMfsm43RNsMeXJVoeplvTwiLXz/7e3XRxbO4GA5LmLwv/Zk
VAtcO3zdOjqOXN5yWs0SqOWlzrVWEqSRAXTVgWc21tvmPjMuHEySH4UeyDwDmvUUeY33EI6PUYq6
A0CmiEgXXkTxlLK7pPXGQJN6LEf1FIv9AYpQNQj2YcrcEyPvvHyR6qQ8wBvHlgRGQ3HGIdeKOUtM
N6jXtWW/obsl5tLKN3dqhCPkyhk5eRWTJDe2QYeFn8Ts2Yg9lBttYZUMb+jyOaVtjym2hgCFA3cG
aO1N0bPW0axg652dkaZaGc6EE4PpIKwTkWjd6eE/u96kIU10yUG2DBB73G/Bateh02v0S8ca0Coi
9oFASXYCrMUu6UC5NYFOxOL18bOmnxKtJioZJ/r+2ttUJD0auDAHP+mlzuIms/su6QRVNNu51f31
gaKBZV1i56+LJzgVLkbn3qvMCg5yr3K707YQ/8op7SSWZN2/bPtVSP37hOD3InvYWc/uH/222XBk
EuWQcD1GYTUtSqxPNlnFMGnGi8KZSvMLP7gXYEXSCWw+ZDcoFKM6KoUpdx98AJCsLV8m2kvzZRzj
ED8cEsDG1/raTdzLp0lBmJjR66m/chwsbQ/gGIJTgN2zyGHj6CPGyJVeVVyvSF/zlyrRier4i69e
epvvn8CYdOQS4vHBOwlRxEBChH0Q2RC/odD92VqFIdUT/m8HqaR4abqce3lEO3Rnt9lECvsEollY
Li8pa6fxZ2l1nJM0RNcDJRmN5pzgjTIZtlzUpmG3ThHOV047t5+iFkXn33HwWW1jLuZXtsTl5uhu
pWmV8LAORbWppZQYoDLpef40ZUwy1bvGVWiWgPr0h4cchn41OzYo177efd+cQrNB7NZdifNExdfC
Ac9ntl17xGhwmnhxzTn1Ejaqi531CxghF7RRJ582/xfTMGUER4qvZ/p954MXlHhbIaMnxapqK32c
TR/2pc9uPTz/0+St2t7Milr+1QcTocLrECaDDd+6wun6E9hi5ibLUkfjX8oatU5moxD0zfAEW5h9
OYaVmXXRjq2WX+mNNUjrTh4QL43LxrFvbUC4tZ80UN5Ntd07HOiOa1pyM3CYwwxaCn/+vXsmJ5Sp
TDyM1BICwl4dwVuufAvhSBeeI45HDAw4wX+43lnU1egaspF7RfUj23P5hVaFFYBuU4scUIRMjZzi
27elL+/yO+h9XnEPvb32eqS2RgyQpUhglrLEWwP/z1yo7rWznXLESsU34xgXpA7+QDvEQl5hmckD
d/u4cXiVp09TgRhkDL/vHFnW6KWhmWKFIU3ZjsS8+oDwz2Mj2+LYZqFFDWv2c7vrsFMMJKQTfFNX
xrrnL0kt98udyrl5fbOm1zse1/b0b/ntGKqpbsha4XjQt65Aubr3rgSI046Lu8l5RgLbEXsbxeM1
9P++fPwUhisDzyMpIjvGcWBYJwtzDrkEfQBtV0Ey/9zGi/gsqWWBx1L3t4vifu0BUO2qRY9ZMLgo
AQlI8Ro4AtoWJKXvV4vUxREOvJ3sq+TxMZ+BAFvD7/yFhAccWuMBKqEBd/nnIFQ4vOcqXEhFAdMc
9nOZEPDRaz+BHPmT8GRI2bOZf3MROxlVevzngXkR27V5YWqZy2hkXS2xN6UVCKZA63DGDx94EjjZ
wgjtRMBhS9zXXpvW/BnJMZFMNe7kUZa9ULk8kok9C4IqXaWVtPVSXatrF8c7wBuWpaKMoRHNyMRI
vgQ0muXBCQ66KEqKk/Lr9FbEH+lenajn0bNT0tvaGAegC2VB3ZMYF60Os1F68NlEOSfSfQc7Athv
HJqJK0Hqme/Z9NQgiwk+vU1fbI9srLavYsiBm6KU4eTAlrFT5itUA6Dp848bLaDRbUo51h2A1Rlb
zmjViRN0A+PI5/INLLSnuHksOQs7+0OBF/pFF5ezC+nUmo6Gmv8j7afO2E+/VwaBb++gorvw3z5H
voAJz6IkYyzqmpnJArCyB/Qv/0NQapptJy9MWOjA8HwPDavFVG0jm3qfh7OI2ZfAwaEmLSND4GoZ
5Qm7gVA/RB5k8hgX265c2RX1z+LDDrcdjLlhPgKj3IxBe5OLHeYmo2HtN/f8Vc+4q83n80Hlf1/5
FqnvCiY++ORKT/H1a9A9gZfvyyGyYwFiRa3ZLCoSFopYST+npceUS7GwTDcnjTN3RLqbx3eLWgfQ
Fp3Tu4FXQxeAtahkfniWtqYsHyCv/eC+85z3MClYtbd15U4LSXc/zwV5cS3XiYW/KO6LZTjof9LW
c8U1ZYoYQqloRUMhMeVse0XZkDGqLaQOQnv4A9qnT16SyLdk8+d+qcVWlWbhRKKmE5gxYTErTZSF
jRNMwykvEn5H5sR74JU8VKMHiockpWnvhsOhQG/97KWjOhiISYueOIRMbA06QYFw0do/n/He9uXE
CVrqu9MU4Xmrn0/4aY7G2WfywmsVTrhAj0SvrYdaeXQ380pQmIDVnL6i3NqoFf3qirwksvNQS2ch
Oo8GyuZ88hRvKU6OoRR/eJNAH2oC6NXVej9Myes2dUH0MWGqWQ8or+JtFpH66AeHYvbz8RdsDMdV
T/WLmhCQLWcyOt9NQxCLfqbdqyfHGo5KLHsT/RycqjOHy0ju2Q6prj0h61ZZ9/vMUuH6d/b9XbIb
meb2OH8Tp9I8traqpAqZ2cTMrahBxswa7W5AWXNPEzyP22wqJZDCmmeSVx0Qp6T1kIUOs6Iy2V4D
uHuV+nDTrYnZiIkqevuK3BNK10g/A9KbQR2pDuB7XosQD86eIFNxngDnnRxjaec1JsMpmbbG6OyB
As5lMPaMxu7uUC9YWADCo3VXtab58vAyI7iQt0T7c2ov80azEuzYEszssDxXqnl5hdeYxTsgF14c
Z+TcSB7q7E2Bedd5x8o/SeZEqCV8Vs/Fh1wLXm768CxihrapRFmbXfyFVA/cPrJ75FmC4OVXRMMc
xPyIcR9QZYI6Kf6BUwHC2v4syeuNTEunirYvmZrlAvMFlsPzIPfKcYznRriG0TEDq58oE5j00urs
bBO42+2R+bLr1HxniWuc7Ur+Q23z+qN5VHdGwM0WC0rjKuudxpQ+jqaJQOdF/xpQKWvhuK0BL7AV
LqRtQJZMWYyZPEt3KAYaReJGZCYo5O5eUnNhRsfaKJWENSZ9JBCds01sxkPJ7qB1ZOdDxA3VMuGs
pzhrF5o/A25iTJO//faMoW8mo8LtpQzkUzBw6DmsVWpx/4l2hYaKTM9ChlrFRN4pjBwjyYLnDEVP
ejybRka340F3oo+l58YqtzKe9dPrNdEUCK+z0bVOYZNf/Ms9pTziaG0hYlzw4SflgOC/rXBPobFd
qCx4GkOJv0qnpT6qcXHT/LMncn3Ojk1icvt+WBhTLxNijts4+Uu/rdnqvlf+6UuYFz3hjWa700yj
wHTYTAEk3Z0KmoWx1H40Fn8RSYE6hPGhC2j5DgaM/2Xy78sg168AyO7HkALBFdqbAVaBnbeNt2qE
sLr633tOJ1qh6NSh21mgcsmaxKC8oaJW2eo21A1pp+h4ERjf2ixc+JfkEdxF4DLGEnfQYrUhVyLZ
xyZS8y4OQcgM2LpoEeWihHuAqMcPdvlBTgwSLCt5yTwuzg2kBZbBNxtXeMQic/1jqICDx4fZn0Zw
bThfO3dYhWbHuVrcpeeALY4yZLmEaa/+Tql3R4veIuDF32aKIkV+0A3cGoPdbNpO9E1iC8kfM0Qv
/pyOChW3uiT2dhhFS6h/Cm1c5nB2x35xV0JdH4ZiYTfuWtDD2YXFUBKL06MOgNIpsxYJWUMwTWL9
1bYDjchMQuNwFVnnViDmszmgV1Jxp8TUvTbENqQq+sfV/GnUAGuaGlp33WAnTjTY+uC1LB+PatZo
Bs/zLT8MxnkwIEtb2dOnTnw2bKbc4Yvb/s85+3DbUjPYi/I0JW5QjVV1X2ObN85mKaPE4jQHEEx4
NIDW7iBz3jV1DNJJqv9XwRL00AOEyDt21mdtSYSWHOiuAWa/ihnfSOnc4aLiZnqtLi2d5rl7FOKS
xMymzq2JvIQIUPD06t2y6mrFZQYk/WyoTLbbWbyL1wOR08rcEcVUFf3WHckf03689mnqh3AQG82z
gnF/OVthbedPE9xxH+NAZj2znqHrMlFeqYwRhB2k+kwXDwwVv86rzVVJcG3sheu/NHfCJAKd1xM6
Dltqhm9Qfv2AR310ammmGrYh42bOyt8g9HmMLun1oeSz2363rmjbEsirsPwCfwUoDnzD3rkv9uFq
o4OBEFTCLa79OFo/i2blpfmfmykGRZkxBQPfX01w4/e5RyBI0vvoUsaYDkIeQ7EhO/LMdiE4GwTQ
XSix10h6hW4XUqj/ZtfvJZlCDJCNUdlYIaYH2LnwHJJdT4N8yjbmbGR0PaNrv3/6aIHNJbxSFCt6
BBl1vsp0uILKXild6yFmL7dyR2lkV13JVvj4hvWN+8Rle/jvch3rgrjPtfseGuZ4dIs5UVeZztss
qW4G/SRHyAiDjRAn07CrXQNg641JDm97CceW6m+ZzmrWjZ7SmodyIGdf/TCsunu0uHqUTsTEsPl6
Q0DDzyuXpgr9lYLvc7gleOR4IuqJ+7p9yVasmwJQ2JjxUNKGTqM2DoHw8RoTkt0smAfjlizmTn4c
EehRAz1T3PUmdCsZtzaRZm6YhpPaVe3iz3+0pOk5QR7WwP/3/htmWvVTz1WBIBoAYme8dxgJhedS
ab7fMHKk8ugByXlEMM3h342+Z17c24yc3KdtlFug2VSg+PGaMp8B6NMIGeUdNIkNl24qycM9NBd7
l5vZGnh0G++aX4yqziiu4RDDOD9+Y9uvsJo/L3EdBkqZiUUc3sOyjXOEZ/le9d4aRxTqB6frzYxR
X//1+gxG1vWIbHUPFD08Cv82JjKCZfDWSNceCe4TUsu1je90ku08Mzt1qo9jHe2d8TKHV5Q9eMz6
YgtZH0Wz1s1Zw9uPs5z0dEedR1Gq1jOuY3CWmJNq03i3RzYlI28OGjTCCT6nXmp58f9rJbYFVy6E
6QHzF8bkEdfTKqtZqBdvEOt06HOne2JMGRHfkt8QcCQI0w8/NhORuCb64xtNmPyjZapJO0+xXLUI
J0cFLRP0QzFwkQbb2xy8yB3uvNDzqflIGYYCVmomOOOr/MyaYur6ehh9qRRXPKs+0n4dglJhECbF
ReTNjWIFFHDHO3ScmsHYia/7GVSUzv1SOBWa1lzxtkiwhTjJ7cLql9vQcyO5mbSBznrrWhUtMmHg
I6zk1DY75f8ytiWgQM64eQxCEjzRrusyLu6mqBREt+2Jq/Q5xvEja1VmTNP97Klp4gIwuE3GFUwd
42Nz2iFMvpqMHvXctyZ/5XXmxGEzJOyFP1whfwnmxplGW7ST1HBmXxVfYzFnFpzP32t3TY3uDiV/
p5+TlRJZW/lZGpZXjVo4KwOZJhoiHdOg6+nLmZ8Ook1dyJpkJbR8iWjrRjGXfefmO3tk9h9FTpL2
MAEr5MPgpG1PjSrPGlbK1sNjxBJfOJL0haw3q4P1FYqHUQmaOtEnDGO7MEcJuvP9JuhVHMk+3lwk
Tu2XFuCbn5j6iKjElBbnlrOCxNViGVwV39FfjPD4DaHyldkOl0N2WEtTL8qQRItj5lFkY4E75kp5
h4lfmL4G35b5XtX21gZPa8lonVH5OZc9DmKoc7nlE9eyOkM7nzfxefeBa9QtJ50D5CsOJkQlVowi
ZXxtU0VHCGQ5PJCu8HaUPZylhaASWRLG3NvWPBUtvkP9Igzgfrk5dW9PvYddgDZcAXCW96NV0OF9
klNljB45lpqYnf4TUQhxbP3CXh2MzlLu3mhKNCJ/ySzkrPYN0+JzjC57ftNHD60B9oymj/+cQvIV
LPjSMqFJiCkexJATEiNC02Aypr+ul2COEXNUM1XBgQsETvmCCLMjd6dRf4KaA68oJ6slMxyBBNTw
oZMw4V363qPVxUSKpgpMVYKcA7VhDR4/skGbemWGD/gM8BgcklyXCGE/7Bt2nkig4nJ1lVUoaBjS
pGrKiaStX/0kTCbmej0tUYX9RwllwvQK8oO82fnH++1hn0+h3LY5BTZY5Vsvs2Roh0DTb0g1+pKf
LuoSANV34C8GyElk5JLhAZltS2SL/MTOtNNXI7wDN+RrOG3orPBnTMffDV57OgG7yAABmUBZgOUY
R7kIzzSiDwmeNpGnHoxnyFcLB3i3aAz3Le8/WF1Ao9aTbXpALY+/QPl8e4tP7OJNL6epyKvshBC+
kdQbm+N7Jok08dW8Pr3mtPJd7calw+/oqx4vdWJjiykNLfIj3nolyatX8GjSX5btvZDXAiAJYqJx
RKe5ddCixkr30EYtDYCbDmANJxtLZ+7ryU+ASKPX6KrY+9glDrppMTyZaHAS7fEp4bJcmMR7YHaU
2pq4FyGoL0Pe8h/gZgGt9h0mpBDTq9KurT1gU7NC+9Hb8PYVU1yCkzWVZVGBoD0wOlfjHdgQGS3h
vxy4ZfkBgc24HTce/XFHKNdJPyDwJ5nwkO/RISHdd9be3LLU8YWRdHEZ6NfHZT0Qiyihu6eT3gVE
16FhBa3J8HcTNjkO3eHmxN7mvEY3nJha55MGEG/I/s41HQIKpA9V9Ad3d2IHblC+oxnHZLhalZhs
+y+j4lKee4R4icCk4Ke1YP2CuHoZnmUGDI8hgpBRhM6dUk9k974kId8v0ukoF3Ks6/xGlFHETdds
6q3fZz3RHkWw1nvSHTMFozdxMPhByrcBRW+kOTfALixzgMYm6EQTlrtvMv0s3hpeZmsU91P/ylxg
7KzpjZR/aTiEA6tpYrNjqbenKCHVMfv5sO/Yvtd455ofTtURRxHbM5Qfj1LorvZEfLYFX3bCvMt3
J5rxvJeG0nVe2O2Q6tqtrpEjuqlnCowWnKy5wxtePFcUYdR7SIE4v+HyHjYSsfm/xehxA3rc7Yjj
pH/MtUhlZW/WnQuv+a+mJ6vvTkeSOGj1u5MMK/pk8Gtf3GXub0NUB5axtEGcS0OAkD2+JnykxbcC
Qxjat0eYTDz4BTzQuvNWvyGQMIWlEEbdzV/Co5c87cu+rIwypzIwZGR1SFLSI+/rgxSq+BYLJ+pj
xMgQRuPVPC7oyQbBkNPw3r0FSqDU7kS0yxHyE0hBrav6UUmWawrYgcIJDthzPZTYz1skAq1tqmwH
iBWSy4187t8Y4MQi5cabf8kyxZ/WAYKkGrtkf5MUhs8S8oaBPg9YVLdMfSdJn/6ickfLelDRnJeQ
unRAXmGNArRcfGl4eMwpm/T0E7jutA3uWH0wmw95PDtIYLeiYuXID1o22zz2MjCR/qezxIM4JFed
fCpjAXn4Jegxejf+IDMMMRPY4iT/DVdc30/QklIHVWPoPngrH/wLzHbNRTb9nx70oImf0r7xVuY2
hQQ0WHVFtAKa1ZeK52Ewt4VgU4+3Y9SYLIW/uAHBziFPaK7NIYmN0Lv7BrWUdtxqslWWPbsOjIs+
mzvr9Cy1DCewbvkPWCN7txQhS1CPlDbWmvZnZNcc2t1jVTSpdaFMPHA3DBb18ZDqyffSeIxSjmNB
z5NYebZJRwLRPTSLeyNGmKfQ6R23W8PGoSm8F30GEJjJHtRxxZhI9cL04hGm+Enx2B/j7j8YZoM3
kWiGaNaAmQYNom10fXgaLfdeMCTe6OevrnHZBilwqp6u/iFW6bIsNOyIUIebO3VQc2EZo2x/21fr
G1/IUUT325knsdxp6s9rPClqU1YZOSVtr29D+rOoy9i6GkUN/zhE3l63FHTGT49XkTKwtoAGI1KB
iKslW0+8Qm5T4oSiEYfjHV/hWlq202dBhODxjaWYASr3jbHG+MDugPib7mn6RjSt8WRp5qVTSMaf
+5F3aCrL1bbGumrdteGB7zPcAClk+ZoAuoyx9OL6ztDzSXhUqpxyLHzrhC/dKq9qH1GEHMQSF4EL
89eEmCO0bXagMneky/iRE/+4wMKHMen0fj9f1i3p93Elnmwjn5d6Sinv3qIGMEzvPDCExJEDCuPx
PbgWToI03SYDNRK40VCJf0GQTn29dbFh9EKwivXd/T06EvcgkvCKg1TLU0dswVbvm7zTuKYmZN2o
6YMKJAdYcYjHswrhrXPui0U9l9lsUMEmKZGmJ3ZvSs6BxReRzXt0w7HB/cyCsCODswiN3DzXRK1c
rCI+W63iy0+Mr67R66B0GZfo/42qihyZUOpPpIhZb8qPPsmV+Dng7YZLKyUscLyrZ+0YgcpsFfL5
z6DGSS1PO2+bER7IZgqlp8/4jfSs0XOvZ9owa2S0A7g4RKLWBAoBEegNC3sk3zy6/K0pmK7rDKo8
+8BfZbJ970Gl3SOEF+n+AJSKBjoyPS3k6mKnjeX6Fo82OK9VWm2E/tYkqyZBQmY/FMUZ54zMNQsK
iWLs/DYx9vTVJ/bCFoQnuv4zLbQHozzcA/0gZUyzEtf9kfJ8wHWlUvHAbvNkJJhrq8YqDT5UJAO4
wcLrP+t3Fl86OiFRBmwK1RQhYlV4XKnHSsnEqaquUt+YCdvBfHtnVxcXYOFgZaEvzuxGrgVIyfyR
xFEEmQkJJj8TLjG9a6fb8YixQPwSBXCce7P6PVMHaWu7o/s0ZQfNqHuliv3bLV0roXQD6qVNupaV
VomAKtkJagR5e9IdsGhlSt8x+i5HPyK6S9dUQV297SRBuUXhm8ut/67U82ecWtlZtWyJSy1rEnDT
xDazv1Gux6GB0aUQ+7d3kepP3TjTlJnXyj6ABtBexoHWlYHqdlcqLZb6RpAgZINg8in1HdtLnHEn
JjbEZ7sL9etArXANPd4UIRegJjTuzelaCc1UVDvhtyhrAg7NKtaPAhK7icUCB1XGj8KhJInihlp3
rljcrboE1oi2jRoydJpIukYNkfEkZajO74AQeJO1MnwLxcjFFYTr4oLIazWkpXDc2MbfghiYs0UJ
zxs6PmEaRH0Wi/3h6OCh/uuzEiNSPxYuMuA+rcHE/Wsy77p7kPQDREccALe+hC4uC9RbXEvThopS
ttgdI7fUuVAZHuP0IhCwfUtpdzanmp2sIU1p1TB9vCYkdUzRgIDpJY/0EUKFozxFb0nLAu0jZjf6
08LnAiE1zKv8pli0n6YsXMVkvYs6lmyf9DpOGntGEQXrZ+ra2Vctc04dppmAPFXwljRCJIo11ZF5
FMdM8VHMEzGjXdH8g6GW4C5qvXx3eRVTtSBimbXwz5ugQ6ua3wSlOk46jUXKg9iWp6mYSd/fbRP/
hRwiA+KwizienVjVKRTyyjNWIvjS0+TkFZCfHRgoE6C6NjJQOO9jPO5CjtNjv+pzfwceffQSdqaZ
jAtquafNp5GZ/966PEhv81vApzBRixmPHR658nvv/SgGtoLhYfH+pdb4SWMrD/+PLf3ljRYePcn5
z+rF2x4TKMfY5Ber6bbvTNh+Ah1gSMPOa6GHj67MaaZ7IMNyAeowl1hywP/3YXFGKeSnyqOq4lLh
g//UAeqFxOtssAEkzVxAiq83JL3oSKvkNrZ6r5pCfhEDTIBBfAMx8revGX6b9N0UFieIOFGND+nJ
uV4V3XnhLtOoslnHQbo4SC0VS3bahwWO+tW/+iqMFX1WIKSYav7olOnvrR1OQPD3CwSb/DhBMJ9c
XFcaZbyovMB9koZxcqu1IsTKIf61iWBu8rAkWc84qSQ4Qm5YbDNOcTPUzjdo9Wce7RFd2DiMO5Q2
wlifhhDdItyzANUiECqpnyZT9JMaJsNVBCweY15jsXVFXk7zohlaQUjbILHnBJMSfCjbHzgDTtfZ
+LkjD1GUBC/CaFAkDgqeMdCga3c9NcSI4hwCGWHey5yVeLt4zSAhDTy642dcMvw7cA/vzo3Gujwa
c7IYrx3tMMQTPXxnbdBmYxUuTea5vBGb/SaRTXUbElp9BQMUkx4Z25yocII17nVRgHKIMzBc+ujS
/nyeEDvD9S0rYQi9abfrOPnZz7y9RIV20op9pfVgoPNcey/yPChdOT3dYO8QOowN4roMzyg+2+uB
ROd+VceHiw/lANyBqjk6/y1m6AKuPCBuOSdJ1lwxhSIUxtkA6mvqGgSLJf4IELQPE6P7A51t0Agm
IVA/PwJ4Vt9I3UtsDdU/2aV9+8Gb8I50lSpcUjBFerLr+R68IuKNZQbN0pG6RhcNpc5vHWlA0w+T
0qX907UptFJ6EciGXwrULXhlPNFvPlVLpe6Ib5GHLBbRzFgsxVpD7QxYkWaw8ewey6bhl5a5+tKX
cUE1MVFdtrx7eXERlqeXwkZk7963rAYhYS37aTL9thWObV2jXAFrhVoKE5z4TC/4HUUSdun8WkNA
wACL5MnF/U+I9LTniyTEc8pweCNKsvMpI53H8MX+UsGby/CB5+lDcOHmFXLC2oSr2ZGzdBXUeu2O
ftMfThWG6m02LODDYe+zzUTs3qWCdbHnhyxk8GoUNvndrx7Gs6TuCwVVOlWuWEnNMRvh5883n+Dn
e8CltRa0db0uy5yw4bCszLManOKDda3HpUn/iD0f61+zyPKdlgEmHBJBHxY55q0jcrSQ3sZ1D9R2
g6sE+x1ZUICp99ciYX53TMz5x2fztxqulmc3JyctOjDiA9A8UdI6LxO6YKTV2Rb3iESSS/J2phOU
lLlSN6uKZm9iWbOT7wC65cTejxkxvqi6NuYcsinD2TCawV1WLKIfWPKmlLG2tuS9MbtGTcaEmHX6
eXbcZdYjZ47d4T78AuafCs1Vjk2nkKNrNYNtEdkavGYcExq/LM5F1CjpRtXSkJOgFVUG6jQoY05V
iqUQvkJnvgACjTbhPoJWyio121u2midV4d5aUQ1lswrll19JV5zHNVs/XFg44M8vLy/r7wFrXfX9
jwrWEG6W8mo1foxn9csTRxD/hTNDVgNyt7gwOU2D4ytT8fa+JzplZ2sB4xrkE907Lfyd/vXwdDIx
4EfMpwZexlOzERzi5TsW3shqZh8/i11g2M7k0uSxroLUQbuGKsS5GUBU/njGJ28EAR+A8l15gIdH
GjfJCPyOtwSgL9PgzYX25EBOGyrAwPOFdBg5nMKzIzZyqLr12H1xBnXf74uHt5fZnKOXCmq3IGTE
rd9VwRAM4e9YTOdIbJewLbg073tg1XYGEfDkUBhn7fGuJ3eUPTuoTCdcY2dp629PPX1LcddlvAp8
0sQKKScYTsvprtQEKT8aNRN6JhTY5EQQS8KaAwY3DbMcwZkp8oT9e4hd4ZsrDR/VaXfhez3Yw5x5
uuzAg+4hdYy2QBm1yuG7DiZiwpcZrH2qCJlzHYox9ajT3mUWp95EEBsVOb5N4iVanXZ7YB9F49Rd
YNVV9WjDXFezvak1VVkttTHEc2dMq4mMfNOhJ+o14M/Y4UkWcJCSYPqzWWj8A5NYlU8mp8ChsLZq
51n9R3hPI9gSuzm5aC3n4w4h5oyd4CQXopO7zGB4j3TfwbrGcP3ssN7osh0lZTURGw9cLcMdUAig
QvRiiPgLaflnkd2ruDwcrts+J7oy4uMOw6iYEJzOSIwOqGRy5efA2nVo9qqxD2zvfbHQGZyTzADP
iATnJ3VbI2ZPHMaW+uas7cUJWUOzMzOeE8dOiGXYz6M9Q9HO2fRIChaAjk5U+1PxjyPbp16DHxOx
A+q44ABt/Y2n3KqH2Sba3NW8EVsLkHMVIG6yi0YuSqoT26I+zxlPAdDNlMxVD1RL9/LJU0AUfufY
SJRXG6XvgN+XU6dD2iLlIVmV2xW/qE8q8e3/CzYUilQZh9uwXeoKIrsTkwPlgJYP1KFsRIWqKF83
9uJy19PuxHXtewYQxt77TMau+5KJBAW454P6GPRAFn93AcwwHbxlym4cA/emcqNM5HaqRCVSFQO0
w4M10tp1NLrzugQChXsHEVjkfIMU+fpi/+jfAKfp7gQJWJ9zZKTydiNOJm7MpAZ3WxNk2/JXrf8w
13WZ1zS6XM9U0VcfoD3OXxlQ7ONlhGm4CtqMMMLvbo1Qq3Q9YP64dtLOejNMZWb8dE3M47W/G/9+
VizR/El754TR6PEZAWV9aL9Ax82VTv5yBdbZqY6KtcRxQ2bj/5rQZ3Y0iUlFIj3yr0rAjx8P31A/
/gb5QjDms/a5ipq4Smh98LvrSKUe/KjHQP+zFruz5cF9t54XlEQqzKQybneVle/vbhdYS/NDpwoM
B5H6lmWlyAeTd8E43jlRJLi5EpB4IKVVvfmcqFqXZNYS90RJ0clsJYxQ/UcLarnQSzP37NQjrJpD
75x574w8j2BnYZywf/9om1i857kZLJ4l1IhwisD9DDOlPL9j+8vm10v3sIv2CW/qphTHqWgQcsmF
ukOi6pDCbxTSXc9vFI9sbAq0qi70VO/zCENlaaVxaDEmRetMEPaf6ayJVirVAMs4f4egUaEwAguv
KwmVC/pYojzlyGQxShx0sNbdEQh5UZS4gUolc72d5gzvTrE4rhxUiO7g/GR1QpfhcE7CDEr13fWV
SxY5/KRNO8L2D74n5JItoVYXum2YKOeZ5E50EsdUqvmUNpSkl0kS/MxIVG3fW649n7e9HVrhp8OZ
Oa0OZoBy0MHEn9aA54DWwbBR/iKdNU6eKnyFU1XiLL9+BByeB3XeuFoMQTQk0+bGnb5QJn7xVLoF
7f5sXpBcDAm9Qy/ppdX8+fJolABiu/OYXL7Ibi5BFOtvLkQLC1KgWbGMH7axxvcV7ulIXYW+CRSI
J6Rc61yc5EZaEl2wDXDButb0b3Dn7gmML+5PlU3P73+JHsv6ATWJFIJnz+TWWJeIwiH1l45kb8U0
nZ5lZc3j9jnwkyGXK0yBOV+LD+KqBtFsVjofZl6Xt+FfwItH9GZJEQr637NsLp28fGXBw1dVS2G1
/DIEUX8uljDx2fOWeQ1QVZLHgQnp+uiIjC68WD5LfO7e8RxUHnSZGc5oIArbKpnVSMNZwhyUzoGV
ePdcwdmG7+h1tyAxWMdv+8dxpQcGKerA++z9JdH4EmHedymWqfWHbB15iPSL5WHjRB66IjF07Vqd
DithLzBhjxGu5A9WREJrBCvOSi/HRK+3FF3heeuKgXsEc4PBoul2JIlU46PkmHLPArEJy2f7xpE3
iFyA/eG7B8vZsuuoUIEMvw6CI+M/4h22C7ktQn7CUuEBcZP+SMeIzA6Xf9JKB6sN+zNgV585b3mm
Wl0rQQGgX2saJDDRAYsRsfuWVxCQO699lqipvWqwQIILY0RVD1jAliS9E0CFfVi6/ikTDccpr72+
k3S+VfQbZJFvCJ7kM25F8Zp8ZX9hARy3T+z4LR/+YIm9vrRtikOkOZ29bnNOuaFNarBF8OIKj4jS
O5x+Ds9wtAwGEVFRTB2yRQdZ/b6/N2sN0zdTJBw0p4suq30R58M+C6UdVO4AAYR9UVNmZq2HeLco
6q5xRwZdHFX9jVaHIjKxkwaMI9EK4dW669rWNL3Mh0cBlKCnbbvcaruuA2VyMTvbPrgj5z2Yew+r
LFjTTBxPAUvTmNTldCG0uGhczkCcg5Q5M1ysaj6+750SoQEjEor0B64aBR4g5vz0se4cluxH5xXr
pGBSXlXP63b8eO02cSdo7rN6eprEkIKL7XvWZAaEcNVgFJXon9ZTa67sqeDA0wbrDr4wqWHE1qC1
89IClBUOOVJUFckdZli3AmSgCGOac+MnNTa67JurcxJ36zunzf9MAgPZTcAhVWnqPDmhmS/DODLQ
OjSYYnVLaXCZPcMKBai+R0XOeLRpukD3qP7O+4DciYxM5PkN+CgseHaV6a5c+bBqabb7rj0j4tK8
6zsTWrBWNXXSg4/ygKgtYk1T/C9f3owokn3Z6ON3kpJ8PwsQACYpUJLu2hyWpXq/cks6be7Jpzeb
Rorf56JC9YESmWPGT7WyaRpDnLAf6U5r7VevZKnMpmdwHk3zO9C19p1Ec69Av4exO4RAlj3YRE+F
EDLY0Fj5xpbfjgs+0sfyie1PteuiYa2hiEQHeQ7HUMDs8Li7uB7/5jIhp6C8ZmEucDUSgz1wvL8y
tQzy93on7AnHIAg3jTA811ulqgfdA/SYuUcdOz+V595QawMcOu/Tk9hVZY15GKhiXJuYNs0j47Ir
t5liJqnGY43nQCDVlDMUKQiOnkRWti0oomI8MF3CVZCLtKwlrZ31jzc153aVzv3VUwvb5WrXpMdM
57J3vKAgzXS+LQaor3cI3l74jeXCFLn++6HcGRHZbD7/TPmCUohUNx5jTamYZ/rVELR80QkspJRB
JaNViBYtUcjf3qY2Vabk1pIL2PAUYEzl4ZVm66GqUY8/x5dPLHyqfk6sIfTtVggiGVwBtQHvUOWO
eMZGLT8ka9Doof6NTkwUyRPWDO3ZJC23xkZ4F+xNyDWjsgR9XjvV3mrThQDTHSgdRl6N4gk9bobL
gU3fP5Eo7xMVd7RZEPN1jZwFnCARaJlJ4tixFo0BKoxF4+/3iNkrrXa8MGlYUrszKgWVcDikza1e
bBbc4Zt6gkWi7zMGhzhyF3xDFQeSGDxg9GU+H33gyK8wIplSIGtyQNFbfjNYlOmR9HDMYaTWdhdf
F+7INiSG6jQl85PQy4c1YQd+2Z4OijJs59kEkyPk6yxvKSJXUKBKkiTO/d/77IEz/x0+4riepXq/
fMR5JwTERTcFYxm7oOeKSHLrXZzuh0kxdhqc0syVBtdfJdavKh4Rx+D1inC0kPO7HrnaT9STcUy1
QShsseRVVpsVtMjkIlQHamkTiy6bOIX3qwd42CKamPXdXn16jBZj0GYnlRhzjUwTcj2SOdB9vQ0+
g0Gdg2z2UTGhX0OjWWlYUY3zs8dcLsYaDq1o15QmZrNbUie9EXSg/k4+Ws7UqMaFmEXU+T25lt5z
Zp4QZ99cidCHhEEiuFUchx4w+CC5yHkspr/ZF2kOE2teyn+pZzH5azaWHvi92L/taIYCaD4x2HDK
CfJGwizJRHmkbkoWX4ccRvFQrXFgnL9Y2zXXc6t7B8qsK+NtZZ3dxnKRrqADUgh1fAbiErZPgJe+
CE3JXS+q4uhk9EOJHZgc0qahFnn6JShj8eL8uXKLnXElHQgstKFfBgilm3zgibu6KSvdtRmOMpzp
m9j6TJe0UbTjjFBrEG7NOMlm8jjPSXnZhLeV/IM172NovnNjJ9gjDpauOY02Oz0j2mOpSwEHfwHC
B0vfnKwfOSTXhRdqukKI6guqZtjpzJfwmCBWuP2ZmkKqaKs+4IXBb/u/rrThze1xLVaGtAuppK1A
cXyo47/qptcOvZrugx/vW+kF4XguuXhc5rAzcozTN387BvvkYygZuiebEp/E8PsGP6ByajCp8xTj
+OX8kBqZh48wy9/r1vcAmkCFd+xmyrAfelEFcgkkp3ZKUckOQOlBCaQSlV1yRDZdFiF7vKCs5yL9
AjDtfZMQgM0+lvPdZYOIbD3COvGZpMDn7q8Z9oweZxpKtnvBI94X9sfu0N2wCmnciQ0mSDEitDej
AU749R7s31AHCdoEE7obhHvRHc57UiBQua5EOqLShkh7RDNWvAX0Ew9BazAi4x5c0Nbw0du7qU1F
LD83/v1Jo44D8zcWAok5mdbiaMh0i4MD1I5RZJXJYIFPpQO0jRiPSsFZ6D24rWnBCn1+3ukJI8kL
B44jp63iNcRaidR/saI8BA2yEsdd66TGQL5puvH0FfRnMmoMOIkwJdU+WoAq5fTuNTKoeaelJ+i1
j4PMclmhQ8FxzEc871IH33i7YGPzJESO1Tv7enxulAbGC3jycfh7/tRSCQOn/1UDAIjawXUYGlhy
WZHwjniQeQ/DVt8pnupxIFk1JvKPo1PDXe5lDueOxYoQacgQAxPshB7aM9hkQPNSQ0NJ/TKmG9U2
AdLV+nGka2K2saH0830GCEGlErSSfKhIZjhW8ved9h6QbFcnaXh/6495ImB1nRXAgEtNYaIJCLxa
bRN1qs3k0y+qNCp6LcnJst2n+z1plw0K8kzldXRrgRgspW+5JgzVT/tT1AA9jRBajblxZHKfQuSZ
ymsODM7oLgIKpiQQ6qLpBBYGBjLMPndPGz3fUI4SvlaVtaSKfNhJ6hvo2ZddlK8Hplv2AlGame3P
/6AxULKhooyj2ma+o5fJtCZTLuH3IljPy4H8fvPHPS2/7uR1BgmAlaWdVZZUYIkrLD2VKSMMD2ME
vYUKy/RMkzsar4idRQSNJl8BpASLozwW3AVHtCExRHWYySdMzncOEfIevYszHRuyliWoceL4dX9X
s3qVEfhBYsmTW7BziJEnpJHyIeJbPY39UbEE26WuEwwG9r9kB5spPYIsMKu131gAzH0uYXOj/XUk
GldWKcmV25KAZ5GQC7Mf9l2anKLg+hzHAYW9gcNuCy1af1579hFWnZ8kecECRLKJqWwEw4qxXDoK
ru/3BH7Dr5rhJ9qNjr0UrgqljcxBtOr/bmpdaAdoj2qgIM98ot1L5BVakRgpRn2qChopN0VSJioN
vZdWSdq72t/JZG/+dWmm15B4jInIsWeB5vQ4VAMcO3U1mtBrbbDtufYjF42/GLNJrSfP/TGXs6IV
LfXapeCupV9Dize9+nsKTHNfEBGTuHfcjLG3/xaGs/1sAaMoEr0J/4QK77GLlHH/k9rNqSjBVctZ
m/PH316mq+q5vahQeDMPReFX0p27k5L3f1QRPCI9Ai4yr+Kgfh95KimfFX23FF4jWa3iVlM4Lz7Z
OPI0IEoSF+6HzTQdXuY86MzHJOcMCifOPDkm64nKbhRGxgRF24IxrDYDujtg8/3fA3lOBH/xRgNo
jcvhlK3FU9dxtLdgB/upRoQUduppDpcffBu1nZ1ve7uSWhftA5FFlz7W2dodQVr6af2vFcPWbqNh
MZ1lgiGvW6DHUmVjeWBcP8JiOiKKi/hhH7NGWvKMm+0RazNvBZ8XAAAXZMND5LSygiGo2xYxvMvG
oD7tOD/W+bz/SvvIHS6hkcjecRRdaFrtxXvOmIQxHHY0XjULs9TTQRbDzwsGnLUFY/b53dn1IOZ2
HamUPkJ0hSiSq1CivjkOfzhHwme5fsYZpKg1t/jvSHhsuqLJ3025PFxBNdDrrYJVSzWZjnMFsoH5
GhwuToI5toIGK+8WparanqTB8tJS9yRqUFTBzyG8GU66Wv98oGOjTpmQyb/to3hMR5rAeV8zJokY
y8Y69LMugbsda5XX8FMtX0KnarOPDXPWmeKwit6nUKVvIq1YaN3jDgatdMFSsnUNPfr0/ol4uZ/Z
8ymbNNqtHSoLW/5ihTLY2J8e8QYfKtPlHdAaMQC5QWrbHkHdUYDHPqI0o8xXXTjJuVOBcxKOXbnW
dRrBoj7D7Tzi7BKQg3e+pICNqc/wNaE+hU08qyJ+1GAIUQQ3sHhVJUInrF285dDN6phcIFAhQAq8
TvfB9WOyTLqWnWAbAINVRE0GTI8z1vYqRwIQZFViMxwtp3d792eO4EV7xOxrJ5rApiFMGiXQlhvm
nxYX7jJAEeyyOHIbVNRyfqzTJ0J2yZo3E/ImbYnNyjmmfovuSKBUtWKdlouQxs6Wxhdk5gVkw8iu
dyDHj5dALGBt7Eltr5XefSw5uQ5Uo4BF+x53CGD1W+fQPKdynDd3hiTGPMG967677sGWE5s8hDdI
WsMJKneYP3PVoH/801pzHtEtOX2yXjwlSiA177KZufW19PGEdmIPhoEKxaUEcCZ7bwbEuibxM1DN
Ggm10/imTW69pN8DJYpjQaT6Dh+WdAA9+ouQZwo1PYMjMP74kFQXEbX04sTjkAtRBlrZU39piCvS
OxLkZw7x+2LM6oUbsNzGVyY+auQjvRBC1vEPzw0cpTx1hM7m2CznzZag/lbX7xcJAJ26QvuH3Xlv
Ok1DmDjvkkx9VGvA0XGWdLq7KL0QSA3mQJVQ2fOkDKKW16o340A3Ja6AZDh0tIbp+wOH3lLoCp7o
W6mv/r157cSwc81glz1mYZoBngFmM+02/ojMc4R0mjsWyL3zrKOtv7FV3ENZfl7y4u+7ZVgezwAh
5ih5y24yCS50GgdYoTaa98kthG8an9AG/YrLBdcSPGCIlq0iYdkjR4J/ng7Y7Qzq55+z9TuriP0S
jw+mFxuyZUQhmxkH1ZFsvjhiID+ZiK4IuZxWyz+XkPwHoroG3gtoUp5xu5wMts0tv1OCgnnmvsTp
C3mgPINQ7UbOipgzQpA0YfPrdgwOyfw7jGKCA15dtginG5w3AXfLSI6lh/cd9dtzFfjR/WQpOoN2
Cxi70zptPX0B8XzVu/6eOIoqO/Jc+wu2FnZqhDfxQz/UVcmgVUx9SHn6eQ8GIVoZWXgGNhipqPo5
2zEoy8p2hooqr/OBJ6PaI0LgIqAafJOAJlG5SxD22LoO1RwjRVMqmDBIRcXRSm5dbiIXx/QWszZu
Frnt00+HPZj0OUiyQ7uccdrMgOXcKgDQGpNaDkzQjHHS8+cSY0KejAROblJwJhn4gwx3uxwwQvrN
sXxAtc7o12e0o3tiahb8nk7Ac+gpXE92FxdZZ85CdUv0WyIrdyzTxrBMEySIMXjT7kb6K8+GeTYc
bJg6YckUx9zrg5fvmG4CqLlmcUusJB8lNJ/r6asJoAhSEbnc+qHF3B1Tlz57HJ4/5THwv7Jb7cuF
8THIotOqIjIK/UtmkpPrzYzsmZNUeHIys8tn7CulF/fR+KpUapA15K6ZiQqvIFewiL0ps2kf/b4k
hrXGxt9aIEju0o6ZZ2BIT/5uKS5X2OmbN2fvzwOrZ4vijAMqq+6hE2SPEvKxpQYI6RMbjOOatWWR
d7H/Okedrk3BAHnynU3PdeN3D7cDGdZHfRuGWez8CQPUc665MkXeFIeU3SWstDZJj7fJ7HkX4sFm
SkFNknXH0Xotw/Y8NCv16kwhGEqrle4HSV5dp8V7Y5seWrCXtuRNxkIlgc1hm/wyoy+rYKsSf3ut
mmqSlnaFw+AspjGKILVIKzSgpFYkAV07gu/UCNFz7kS/fNWmyMsW0VeZB8ZxnPeLGaTcvOujpPmO
3cImYO7Tnkw91yb4JkYBA7yYRsHeqAa3yRtEEz6xhaTesiZB2ih6sbEG0jCy3/OEQ+QRg59lrwI7
Or39MviWFQFWtgo0lDhrZaCbWAD+GMyPdA4KM1By6SMA4HQHbj8huKasYzXQM5kdXaKy3p1PQ4aL
xtZjld+eL2KFhxOMDMLID3T9IUtDi7h25PbMJTaD6ongdVJqkQxE+KvRWdSFcjP5R//KafTxUWem
4xlWrMNtuMxaF+YUDfzq4BXO4CQnHsNM+Gxvhrk9ZZrzW30nqRqCMHmcNfHvJEcZbE6Bxvt5BDHv
kAJdlFMw5P2w5vFcpSefN1DjGznnj70/WAX1qXgbKGlPwSsmhwmsW31f3it9sCI5FPOFFHvvnHtZ
ow3U56f7MztgKiF5sscH5v+p6RfyBGVO5ReJlhi3rHbuXzzrBZI7nQjErdJUze0NPQqy9bZgYKx3
0JO+kPA37LWttZ9Vjwdq7/6EHtwGm69kN8mWYlkC2WISTVe+6aVBU1lQvZR2sQX+vxCopHTPEJTb
mMkSngGOoDupH8bvpiZNy92W3ST4JjkL7MZ1a6CZm+DbwLmCyuwXdV/kbtm43cncivF4z/YbMtph
RZwYomKe+BEXBWCwcBBYcJYeX9JMbLGzg4RCXZbpiMmKT+hVyiufyfwxcMxPWDzhUfJXTqddf6Z+
OOlZabwwoiyx3g4Ija6m7UZI0lHkgXZBKZrWRT0F7TEFisSR1D83YtARMlh3S23ZnOmDRwFxToZs
UImxHpPxpTTNZDBf/Mo3D5pucaU1fUW7SbBT6yF577Zh81B9OIerYk9iB5huZauoRv61zOcAs70K
7BXxIPlxZ798nuZ/5UjwDSgJZkN7W8NNg6rGGM6djbVt3eY6bF09eEAdxXPBr1mErh2KOAmMWU5t
8BOp5zE/I3bzNsrIDKIDk8Ffr6/KVp43TnkcBQFscgCC1XraBmi69czEgVwp62lLz+I3wWreuuOe
fNFx1AFEyHd7F0T4x5kV2h9NJ6IcVKrZNuPnhrS9zQ+U+1kbPux56YliOdKdZONtBB21CHcJ5RZK
B+4JBrM9vTUyv+T9UaSEZJAd3lr39tvJuKKzZ9roZj/6PhjovCqNB/FlkKXHvXzQWE1ARzce7yCv
u0uPQGZfiI6so6TUlU0W+x0q4klKqVpDnWb0MrnhQc3hgTrqpnBKmXbxPLJRMRt4iY0KUHkYc8XR
w6GsiACrqALgTXMOkQ9D5I5bim6XKeiSZFV5UHxO7fPLenItzHVoXLoJPuG+tkJnwFrcmxPiNxvf
4LsrvG4zSfo90FZQVNDoSJDWxMGm7k3lWt02yoGZeep5nqXgJI8T2usU0GvoWMVU5mTAmHJe1HmC
kTWvWFrY4yPdUiO3527r3ktD2/qkbJ8k71GSfVt/AkvmyMbBDoVmYMeXupN75OqGdM82wLBxO0r0
buVn1N60UBiKY2ML7C7ei6TaicoRK3DyS+qFZ8ED2PnGIHWieURee1v54OMMB4Taq1qpX9WP0XCx
m5Lr4ETXzqWwDNRwoLctJugi0sUtwUOJZEyBR7+o7zOneek6VOuNwhfQo+kONK68FDazR+4jjfGL
T22x94qIMCIkq6EawgjgZT1uvvYi1SAyK0BzxTzWXh8TZCZ7cljsMZSCRlcXErdO3LDLYE3QfUFA
9GEO2nhUHH8LAzDkXxlb6k/LjvQHcky2W9TTxsi3Ksb6P55CT+gs7tfUhHnbXAQ1PeRiAqqcdwiJ
6ksgs8KcnULghHL/o8waaHJEcx9+3KfZ86fWlxgmQWTCZaqy3dTO8C1+QGT7RjbLDuZKYGiesBrU
8ZfkLed2UVGzW6W3RnAox4EKcxNr4C04/s0SHooUQMOGyMo//VhnU44K6HO269toYKDc/RXtDZ/1
7D92thEoa0+Cx7RXwGWL7CrcdOlI/4sOzHbHjSOdhPxJaBZfu3+Q8e2BFtzsZIbRcsnW/xKH6qn7
GH3Lhm/7Bemyd+JH/uVcKYMWWccYG+gqLe40OIJZlDsnrdx5cxMsP3nojCw2Mmw+EKN069uIIFdM
ntEEkaZivDSVw4G0erZA1U1ThUbzFHU+FS6njxatWueQzTxqexuOazUV/ql6eKvbyX9mb3tNFoXY
6/tdajqXhzHKQqFYvKW7vDqFxysRHTSwhfpjtOHwE69ps+hyKj6YU4pa6fXlERwCiEHRogtyT0CP
BD5tf9N09Me/R/G3/7YCKNJvHmlWQPvGJEWWjQFngtz56eozGNj0kvx9cBnB5r2LfA6yugkIsyYb
3wunPSLzLd3vZnGi+4/mKD9e4yvKwcCCr8hKVCmiq+S9DfPIzXOdCwzwA8UfBFfdP3Fn069AkV37
xQnV/BzAJSkNebvRBtXE+eeTh6fpZSFEAhdtgFexfWWRnheAO6DYy5ukmbJ28PCTMX39fl+OP1VN
4J6RIFNUaixQiL6Vw20TLT7FSYp4061IKUjuVsyeU3MOe0PUlRgAAjvb8gZH5vAPWzZZukMSQ7dX
bjGFbH/b/KUP+Uh/vtriFMAF+uf+ZvB6YgN6M8JDikxc7wDP0/7VIuom9Z8ui+u8aPUhY3VtoCUs
1+qzUCVuiANHYLWYjdDFaw/ZAZnCVglQ/xJoBHi/1zv1xErNzNLDFUs4/VkrCjRNPMvhPQmrl3WD
bFYwZnLUXiw27y9a/IF11WJOrgDi5VfGbEfnXokRiCrxp9cc62nlv3KAziQ2kFTqPQJa1ObzPPpu
VC4Q9pDjg1oHuThSR/ft2l0Ecc2Upwpxk9VWuP/qY1h3ayrCKbqdZQpaejfpbbw41LryZ++kXJdk
d1ShON7lyjlaO8xICf5qKraFam/rMy+KXHIVHP9W+AFNB2EwfPmz1QBsKvCGO4TKNYmrWhzsx7df
f55c3yk9DrcMBThhPG16SVmwn1INd/tjWpu0eDSfWOPK8yCLentoT6sB0ZGMVee1pZWRkvyub4kT
X5AhSRFgzhnUzNVPTDP2wpQA5RDE73BaJStQwGkLeQOH6gQ6GZcPDWB6pFKTTL8iCN3M4scbfEwP
c2CwKh/EC8hg6DPWzfZNMzWSP74zT06/G6lzJHBFDyBVM9wIBl6OLUWQBM5eczaFpRxujNM/hfaW
fij+Aa4R8yxI9FIHEx0JOzvNml78fRDVV9i7UqVzAD/vuiM5t2Qkr533Nxmf09D1XLC/NT8qDeb4
/vsenTcby/6B3q4sd4J5r72/8lgFs0bw8tvynAkWfcf93Mzo1yem5vr3azmJ5jF4Jbso+wrpmkP8
qaPIb8rx8uVl7+b9j9u9LwGp79adf1kleUPQ6srbakDzbjceeHNYlU+RmRQWKpF7YoTlbG1iLlTK
JjkAaYJ5d9+VQ7biyZSIp96UQFgFPeB7b8JAYlcmXjr2ZOnC0Q4Vw0nUrPdjmCnEmwPY/yKsx9bc
uEt0wcmP422p3NBtf1SXU4TsFHFq5pmL4Nva7wyqI12jJn0VdJlj4sT/0ukzKPhS1SgW3s7Wi7gQ
nMwNyrZbd/lUhDcp+1I53Nij+WXTqylD0ddJ5+Qh0US6KHoDqJc7JCpublcaouMj3YzOvhtOdwIR
2KDf38RA5Tf0u1Zgyb3BsDEKazlmqLE+5vZRtiINMsKH64nEsbbFN0HRJo5K/L6WPLcHlzIAugWB
i7xISyDmbVRl4/AC4GwKgBW9yU1zHbpYEn0xu1BNWqS/JMI2DhWcE84+5UEGBEkQsDv8981ZFdiu
gn3bIUl61R9nBJ56A0PYT1C8D6LR9ec7T1Y4gJuzgOpQN2WR6xOM7mdCG5fZb5OpSlWr7K5DPaKy
Pov0vFmc81qiN+ZzCRg4L7qYxSqr5TsSwupe0SKNPlmApG+kxNVPNGenEF4+AFVudJ6McntFrL3Y
TdgxENWPjFR0QMrlplkt7XIU58aTvDCNyEIyeUQl6LQEWfWIjx4SiXN7UlYHXB5wi9+/qzPc2lDM
7lGvHTcj74alAm/QeZt8k2Q70E34Xle8tR3+0UaRkUNt1J5ll/Kk2FOzWXiXGihEG5tsgeeAtgf9
cLRKgfEvDsOVqdacUs+biW0hPieaPtrdfZXmRg5nFtpUDOEKWMJ51BvBDw5N19XygLmNjNVVH/Vp
9C7ySPz9Vk0rcoa6pSecgVqthYazEZ6ocLgHRx8leGXjsXmyvdQ8d919gk5Bv0GXa7A26CDlDeBn
djlkvd7Vh2cNcuXJvZVEpOqNL3F6SJpuEZG53Om51A7ZmXm9VOwj8zZw+TKLz99AgJpioALRP+un
IKe3GnrCzNXZCGAe22h800+WALhTpuX5aZ52i5IqvX5HCO3f3bmsmEqTgfiSjr9A2LQZX3qMc9TZ
Ncnk7Fzbil6L5eT7PbEh0ACoIcVK1RgkPVll29p1ghKhNeAUYB7QE51g9C8LbuXmZHVtozyI0AiP
wTSGE8G1YO81meU11aYGo7aqD4h5RUp6JXobgb+zFM17FhbSmrS8nOfOs/9BAJtTDIW8AEEL7czZ
8pOM/BD4L6UrOH2p517OUJD6xN+xb+wKS+AsQSU41T6NEKU1pMT9wZ4DXUrwFUyftnLugJkepfbL
npRSNSKld1zIEIITj6Y8KBZngJelgi0/6ksBLopDWv5yv/DfrcjQYFFmJScOxWRaJpRy6EA9fUge
gUdj28GpapN1zKVagx2ET1hiUNl3YqdF50bwckhSwzod6iD1HMAQr3Xjmtlbxl79JZFgmggzUj3V
hS7ma3ieBcgLwqAdaGf0/qhoKwPfV1u86Z5CI1U8UXkG1M1DWV1R/MkB1cRN+TtxdCuIGzPuAg/S
KAoAbF7sbKKyPr2n75GF66zjHx0+Iad5WFN3F+aUCKQ6yyBBfV+JWOows/ya6ZiK9xSKC6E95RER
g3dlqN3Wa/gD6Fx994OcjH7usal5/N0CgL3SSWJRmLNDpCjbX74zNpz4nScgAS7trZgOP6beJcQ6
iDTQVmukQaFYXhTh4Xb+gmmm8GLSxWWmyvfb/WxaJacejsGOC79aRPnTviuu70m/y3FWiS0j1T5k
ddPlGkbTspEUhnrYuX7HcxP3GCAV1CWnQzvLJtbQyRDR5I3Qj7vYNEKV2pXjA9QUrJAVRi6MeCgi
c9+dJ7WjyGgRUkQA4Y8PtqLoI9La5QUJSaDRIjwe864Tixf4IbKo/pugmPok+rt3Dzdbl0rTt8fK
bUGAibl4ujOcFO/LPTm+nhXpcwLGPfWQCa0G8NMnp0F9x9DsMVDAnR9w5Z66l81GYLqpufZWEY7z
zUVLZqKFwTJlUhj6A86nw5GfskW2AJsWsA2QgkSqvjS8JILhC44APzExIWV41kCvoPFOIIjjxDW/
cbuPSG4nFb3SyB/9IC9APp0UGlcusMVVVnR26LzPnTJ/jOmYK5tt06AGM7BHqLZwenhHfBouPXJt
fRqVf7TYpNEwtnUxommGLnCYPoyDvmHO28c87zMjrYvlD0ZZSPG8wII+qSMfZKMBcCTVeHjairOP
/vMl3QsgClz6njwa2G0Wc/8QtIkdJ1Luaz3UdwxaEsp97Y8YLfOJ5jE4Nlw0p8gNbN7fFublvA3O
d7JTTpN6UbTFUXsTYIgPV59CNQ57kinI5bZ3UQgCl34gXbWPtfUz/K7wrSC+YQNNtq/Hu1i/i+U2
X11godzlBz4hILGigbPzREOUvIHBWDFPc1PhUUjTZe7sKPoHO9/PdF5/rA31tLpbAmx+2FDwT/dM
Icxr/9PyE/rDkFfirf1bP3tyzW7Yna722Bfub+s4fPoHPfYq5psM4cuXGcvJnuqc+Aep58NR2mPO
IYrnWv+1d1O2Gpip14QXgY1Qpva4pogNfXX2RN0FavXbzTtWQUzXAShXYCNXK0Sxw4MwVZ4U+v10
wAS0PgQj13s1XP3Tbjb+qL48NJhnC8wARpGU3UFKhmjT6T8FWY58T+AI0nTR4l4hlqELQziaeMJh
2Bj0UthCsuaXl30jA70lEVDkkt+rK7uzAOnsykraLpE5d/iZdLvFAonYS16n/GiMgKeGtTbg8DmX
keLZlEOHu651EztXypUCnt/vIKwGA2Gbp1b8Xft1qprvRvN5B6HVCDlN4MnamtoYQTouiDSqAFiu
alIiDnOYT9utkRMSFRXSWJ7JMXQo6FWvuSDo16IKhJyDGPMHFKLz1eU4JOJKTtyr7Cx5ktUcyWzW
gk8zlwvvbQCsGEZUJzRHuE+4mK+RnG9WjW+Odz+khsF0OUsZxZcUbsOgIe/rc9QiqCJSTcKJEEZy
pnLsNWTX5AR5S59L9BhGMwgdzt09YDar3jRukLlNad4QZFq0IbjjPzQF0AK0ux7rU8mUVavTYtim
aIwGvxlTH6FUDIVrXe5KsswSkKojsQ93fnmp/aE2kTQ5OaEMOPhnZFoL+y0BI8vgzleu5sUwwrtZ
AIVruB/I3zoJtebVXDdqyAj7UAiFd1cknP/jCp/bIAL4uPROqPQCIfD+Gz2vCj4IVeHGnLSgvrzM
fPePJeVoLooQwTQ4d5D1sZW/QQdVVgMlzU+Pdzi4h1Jgnvs98vL5UjBShzFjQpHhJ9t1lPbKG67X
3cL4QdyAsvbL+U3B/SdkDwBdmci3rUNyQF/yOHxjUUh8KGW4jK7yRSoCuzVquL6CcnlEkpkeanoD
7uIljDTw4bZR0g0inGop7Ottl/SdOxlT5VRadRVGnJWfTdZ4qIRvy8gSxCSHazpKZWHDB7r6QupK
kaetRQ76Xue80lc1oeeQlUwLAQrNPpNcJUlGMMVvhOJ5OTS2rAi3f3rxrKOvEhz7IOPckvDKklwG
6eGyStrl9pu/Vy3G6lCxS4DMc4BxL3/XSDAvZClVHWyd+YTHE3TsIPp9CDZJUhH8yuxaUwRP0bXE
CIZGQj6lckYrhUTF8iiSJT9CtFSy++0+UMv1rPIfq1Pc5dDbQoAwWldVtBjYk28f+uEM4d7fBw1w
7kf+1Ch12hjK0Lk7a3xvo5qy99xIyyRq5NwfAkEkwk5Nbg4T5kKa3Ix7N8C78a5O8x9W5GazQCjj
aXRAsR+pwKCQfQtAb/4L9v143gdlX+rzo01vqoOELDKcCy9XaEoHTq3coqb3ktF2MdGbu1liVZ4R
ery79XuBFE0S15LTLFBa4N6YOQzau6N7cv08gtJD8tpi13q7MxKNOuCb7AMDAKdXx+V0avCPYnhA
3R8CsItqjTdc3FyHVOtySdJvpgAzaZDO0UoO0lE/SWwGb6beGOg0v5asiWtCSm/0QtQIn4UhGOo8
JAXmLNCjpJ7XL3CDEwv6R0Om7UKYlDU7pcNyo8wGIN15Ij2wtwzQE0PGVbG2iGt4uUcsUB7pHe85
1K/hpf5jMzVKkG3c0nhQ5KZorytcz4S8nMlnQIbu1vLdlQE2FTwNOAwpjFRKyTW4s8fWLVph7Gbz
w4CrNPfuuDHJMM9TiXPj/BW82OaNMBoLf2iF4FC8qnZbdFvtqQadHZUEVl3f2eoSa58kH099xU5t
+IPoTF61zzffSarmLLAKP6Vn2+EzHhT+L/sOu8cjJDM7eS6YWHiobwhktjCroNuSkmjrmi3J+9kt
tET0wgSdSuSgv61sPPSmuQL0JcLCJz6yOIGiMZjb0pg2+dqtFu5cVtWAjVSfyVgSwgZ/Dytxjrqm
LqBmErbcqP+fqXQEBkr6cxrcLskc2oE8gKet4CffGEI91MevTsy7JaB61IuZwvbsBoxVzDRAXRgs
pI0ywKBSaCOxfqYsX1aQe0d1FhmvfF/EUnUew7gipNhMQ+MizZY5owqmC6Y6k83CBa5m8a+36xfr
K0DTZ9QTHH24322YVZK/oXK2j16m74zAYYFKMXsxskoPR1vJOlib9NFmLE94hUBnKA6n2Xn5sFuB
ZrNzfgKpiHZXhYHs9rv8k0/mqkEPK6BGvuGYeRAe8uSSe99yi5FdhwL1CDhVpLA37f+PYyHPJsZL
cCMMHo2tVtoHeQJZu4wuMCB0h/pQatjlvusQnKZKYh9j/ANdipTVPBKujjJK/olV+H+Ow+TQsstI
i2cKnM9i/f7OgJSKmEaKdo3nXY3BaRjDzOaiLd8DdEJ/fpqzUOP3GVop1p6xVRXRm1GUkDPoRt9J
9jQu7YyaMRLERIGoSsplE+xFtMYSvcCZshoCNlAtitrINJ5qnD8+2hiwhzBcO9nQUOFrhCyezdsi
tGebyzGQjNnst0ixa4nk5kQYBy8MujIbPaYrYR+BE0Ev6hEjjP+iSljpJI0j/f/L5OBVlTkJARYM
PQilc//hHFY9Vfn3NswqrR46yt09RMwqVSihnRbtuVjVRR5oQzltzG/5fiZtElSWrJ7jzlzy0XaQ
jUufZGHJLDl2OAY251mdJDndMmuO3TvaGNs0oyJYClt8ByEXjXw+j3f9PeE8qKUC9ekC3pPb/QFd
FOfDfke1ICxtFfGxNyRy3lD35wbTVSEDAaRgM5wosZJ08de1vGOiauwIUAU8k1Gr+v1MF+qj1460
146cm6Xsb/nDoHPIgzDaDBgO9J+Mp4Rc9y/vRhrgFzqMV2PNKMx0yUQJqLwMY6wiO8WOppisxfWB
u6yB9Kmkeve0MP616n+VgS/TTYGgIghI8h/YcVe26+ju7qS7UZnh+nMSnWrB03JReGGqpsTYgvun
rpcki9BP9ZZtNUYMVTz4c48PcShLNJylFRS8EghW0TqOWB7DDIwZ6ZWGpSbWXoF2xKInfgazpA2H
7VY9NtxUA1MWduBF4+RpaWuT1pEXY8tqHAglx3mOtc2xu6c1pZCCXl6A37NIAdmfr0hnVKvr+x1M
0qWz7JigVBsQfp67rew5s8oLq7Z/caT2yLgq1iEZkKS7w1fxdFLjBqu09jdWI9+EPHH5e9eO0g0L
jeM+IYmiA15oIWwAR82cELGdZCmhUU/mb7Iv1VbC0ZXXIgLUY5tGIfrw+y+w3w52LjV+ja0DUm41
AdmOZvaonXpvyWtPwbknVgwjaSG04Tbbu/TOKAr/l22VEXTex+AVEsmv0eoLnNV98yvNVdC9F49e
vprDum730Ac91GzwJM0t9+OKVQzyCRz1SlM4vnI5968WhLXSpQ5kVFksda++UNBM2Xa1qlLEF9XN
cHWK6YKPsSWQAMMfq1CJ3b0DdxocEFhdRymtnZADupPYMPTuO4iBr27jN1DMm1tZjrKi9VZQpSKX
3vql2EUSqbzY7k/VXZfKGxNRst9N0Kl9Y6LUqXT2P29GzXfElt6ZFSbtOdvA2rpt0NQZIdhIpwoq
Ci2bl4mjD0C03rMTUkpLBJknORrTNBdjnKWAIxTxSd1gC56/JNJVNrL+zAasa9vzjbbOzuP1Ks/d
OqWi0RRMmJpDkOia2vn/Jp6cEBz8Pa27gxaBsdtuodWkM7XvEWAmBw8s/jQMoSMfNOzkgEISsjcE
s+awkZMjyb9/V88ywR41FRtPidVx+151k8A+qsYDg0rgcNGgOrZu71tHDjb1TipiqVCbempFghNt
qWCKsFWgJUoFsJCBp3a0Qfv6Is6P1MeoveiyjMv2Qxj2UhUVIYoK/A4mOEuWuEYQ3bUaSjlXu2iA
nmeWlHl5xtPG1xqAHnVtYf3hN+9aPQrPEIx57bBgXc8hF42mRLds7grwxuEoVNtfPZyTyPTiMui0
ha/eL/mMVpapzLIYxNNvSXxL2Yk/p+Z8HCEMCSkSA/72DoMKQhAomlB8w1KEjOzDJNpLNT2DsLwe
UORocgCQ1y7CUieP4vrIJxHLGcHaF6Z93dCw0VxbcNPbQVj9kFlNp+3Qxo/KiPzW5Kz7VWqFWgjf
a7DHyTyzsXlw7OTwOPNY92N5lo6FeClOeBLKey0/WY3JnvlmaMDUF601ax0iV2XMlCxA48l1JO1T
4zcBxoYu3HRA2p9lEs6UCXpdguIH2bdRhEZxpcYUAWOqLG0HezcqbkxHwO4Fcaex7lzq9N2Z+t5v
mgLnwMMpBPem/YMaNIm59tUxfzvxPb/q+4wCLvVECJq8t5s6DKrIPEsUwQFzdlqEIWo6tdTmIDl/
iigmbP9UcZJBPgvX77hW5cPlzCD9XJzcwYwhtvWuw2xxozgYZ3VYK2w6zxQ0r3rasIe+heZAfpU5
i2qAgbgIl6A7lnUsP2c9OtXNk7lNLLmngLxvcXHsCAihp6FgwwHajlppztSGYLmoyOtAyAYiM/Pd
HngP6ndZig754yb5B/kCpZTv/5Gix5AFKlCi/cJScC6Fo58hkrDSh/8EoUhxuICm/Sja/4fchmHg
gaPc8+zF/3xlfu6WBoKmKQdWD5ykD438CkWZWlai9MNUqLBo7PVWtVcwo/bebk/snOeB9avkvxgh
JnOopFoJq2T5Vi7Qw5BNOTF360bGC0NdDK8B8pEOFYtE4tv2IZq32tWuzFZ8yj+9goicpCQM8rx6
ajtSAjrhd+R7v8mOUryDy5QusrMJb4q9x4xPB0+mgNIejWL+nm+gURbXhnOpsQRsS2Bu2wFw+Ndx
dBojSReX6biI54Fr1Y+2Xcjpyi2w9lSwQFnhr+M2zqYJWMh+zXzxofWLO2TN+UBZAc4v66TyFp0S
OonkaIXLXWrAYEpLco/smDxrGYNa3Jd2Y44mSTz+iSp92odjwhZ3dG9cg/eyAD8iIKlL6NHEI5UW
FQREf1PJp/c+VPDJ9ErQk+XM096EKO3tOxED7ijhmKgEbxLq0Biah+1rW0ABAdJltVJMvu9qc0zt
K0pyypmWc2St4KH7+vZ/5hu8LrRw+7vD358FJZ13Y5KUTj8v+DbXKc6foGRo3vezLsJ7oPPFw4hg
csA0NPzRWbZc/Q7h45Halj1GOZlVUZn8ns7DZrIZpzYrxFtVoiTm504dDn5MmALGceYBp0R7pYDg
/87PRo6PaunhlfhccfNP1PEEnLEHCpr6Pp7eqQauXdwpSS6qc3Hpbd9dcU2RtodstzQoXp+5gbfv
tW8Qjhh75fydjKYNjHzswL8BumWDE3SPWf9AEhrzIvfXXd+gmt3o3/3Ft4wutDkMtamjL7gSmY9b
E36Z6Yt6BjIz4cqlGRhnd0r7rwMzbLbRuvQzxWPYplrMIcBpNP8Mcfm783PaK1dQDACkQxJq78Be
/kg7fCuU8BeGX9i4xCBfqTBb3Q6b4LfGAOYvhDonHKplM8AUURP9Y6sZx7nGqsPtwvXlnyRV2iXU
/aOs0kUWHeN793DGpArZ2lFQPww+dUGrdH5iH3rZ59LAJJF0VDfnNJPyavb9gEaFg/Pr5kCdHXzb
kqoEHepqQNATaYMXidHg3c+bUaqpLJ23oY8V40PuR37jXo9MjoUhZIM09JMZglF9R5/Ffg+Bku6y
hDOwJF3bU9i1X8Ztferaq8gYNy1/09wF8wsyJq0+5znHNni6bTL0nwDtlBck+bawysEH7qZDvnd4
okKVg2ECq57csbtUiBz+ldlXLGUOLjKiQTGIRRwHL2qpcQjobfkDDGg/KtrzYhCLCCjks3JnOR0H
0r3UTl+mUS0W9UpszXT1bIVvtoDLSQDJ1i9r0KQvXlNZ2oQ3p2FVyE/sfRM4MplRlubZMChJe40r
vDcjaKow4nD2UHw+rI9J67+wBBiX6rZ2WCTd+DHJxjvZ77kT2BH3eeaDlEruYDhLJhGynqd7J2pp
7Q4oHpevr6kJupwh0IAateZuIvpr8LUdZ5MJF0uUWwAprRqWy/5B7kQ8y8HVDp75wmo1u1kuESqf
piY7vA954OTLVfmfRShfQ/NIFEV2dVttNwIPPx6lBhWRuFqgTlSu0EEMo9W2cEfj4KBRsJIp2Uxb
dAeLj/2k06GmSmobEbLQHmEcEpoMoWCAbpnvaC7tkzO1ZnA7dhvxiUoFaY8HtU4FEph+8l4gRQRG
XWVnpM2MS6GHABUYXy+SAP3eTU/pvSvHiMlDx1jHI1InawOh9gHByI70FDA/Zr7oL8qUaLwte5m6
p+WJa7YL9pjCZ5V/Qo+TFX6W8H8/NrQRvq3Saxo9NS95MOUw9QBNNTZFKRpmyyxqBQVJDbpUUK47
wUw2iWQrXMXAkxFC29ZQ1F9/qjm0GvcFUhHXqJ/T0w7CbER9pSZ0mDNAMGWClPDY9iNoFAlIylwL
6wfBHTOD8QE5BXzxIeQcDsMvAr3VClc4fCrc/lJLk+cE5groMplp1OQYnuKTJ+sW6KU6GpOHlpoR
cOOIpWi4YcNx8Xa1d0OgGFX0CXet+e8TZyZSvuv4CBiaQm2rErnP9+cE3+rYjQpB08PWS2uz2U+f
inTBLAxVhmTL5Kr84DK5Xe94sGf96q7ytNSONL8YBZdMMXLP8bC5QaIE6Vj1VzIrpIqV6LGUUUcL
Yq3m6XOpp2jP3cu6g10ZPRuAZoHtFs9j7hUBOsffYKAx5axG5HYXHHhSSFN0pO1Up8Eg6xbHTAqd
8vZ1o7DJIutIKWDeKVHZido7zXc+KDsxj+bUkFYPDlKpOg4/NiZTCQGaNc7CjgjxW0aW3f728mnK
+tCqzMSW65UJpFYwxe3YjwaUk9yRklU7FrZGlBV5F3OYHap42SrN6H3FGAGomz7Zgb2IxpjHQpS0
HayZG1zTniTL2n1+bxjR4qu5FL3647Oa939LYEwo6okgctWV579bblbP2QmBBYjAVS5mfbM4FKd7
IU6wvOuP7Ifa6UXxBG/VWZOOPm3wFP5bLHBSNfkq2wEe5ESHiT5vjiH1rEm7GfJYk9ORxnilEXsR
ABHL6C9k9VCBpwmg+2DB4WUT72H6HWW5JHxLYBuYi2FjhUpSx2Ihiyj8rd4V/KqyzMg/TCTvdy3i
RJk42rntoy418vxLS1H3MCzo+nRkoA5rEyR2rerQd/zT96BCLpLCw1KLHuVBufYuuWW86aRvQw0J
v6/tE/gJdECMm98kGl7fi9ckYEAxWhI3YUT+mYX+LZ0rXBRu3PLrPSReDf0q/cvrhXn0uWhPGqNt
QY1YiqOvzT93yDJHTMAx2L29ytHgZbtL1FTUQ7DB3LhwV9AFjKNhns7Ovancs2IKa+Ob3e/wdC7q
JolW55XM0yyeubD63lzOaLnjZZVQPzD14mwOwUw75PuFUDL+kkIcTjsOu1LHqp9N4lBSLkfb8VhJ
8mopZqcTigODpNOcc83ZY2e6LzSF24MaF89n69CNaGVdUkIqj1HUHvUG9lhjUlHvIznpd8x61R/f
gl1lJq8PFFSNk7dYKHyjLaRJRRiiBCxIH8Kk6qUD30SRMlOEG+4e5XJ01SfiqeGpsiLD5l2rYJ0H
YPsB2HMNKely7ATQ1krk+98qBaJDNtoCFtsaw52wQVhajZoeDt/q/VWBZW0dNS2d7VKwWX6WXx1V
WFVaE9AdJDak+B46lcum2v3dNA6OQvL6HEblY7QKZH7IP6t9Jd4QjesteZT5mrgdgvq1JjRk5/4L
qL0HFJQOVxUp39KozwB9HOchsM1brRf1OLRt3Q0LEdQWrfbkAfwDFDQHvO7UWa/sd75IZ0NAx6A4
OW6JPYdc0m9LwXvYv9T/U2SKzP6xQF2qjaKe8aX/J0Tx5iorF+riAj1R03B0BO3bIiC4wxTW7EQo
56Ptpm8EloV7qI+4yuyqJG1UYCu5Gk1cBhUVqZ9hFhkk4T9ZL89StcQk8foXV6qygXonzmnL9HEK
5ue0CB4twYAjpPohVoaYRlUU96OuVukzUQ3NzSDqJhRoyMR050FBK018YVD62VYtQNor4N7XtTeJ
ivM1PdMU1OTtNbHXBuH7PMkMVEOZpXP1ficJkUP1dtbZskKsXhae7N5WXcgqKan8khKPrPzjAwml
EcgtjgrWQEiMeww93qhg+mDlVofq4lGwW262hwZJpOFIDAY0vE5YQAeVWMorj9xuWLz+IyGvBPq/
2aV01RJSs1ZELHtCZKVz6jNtZBdsJEGNKe5QEOheoPY72pDwLdvB/7v3w1LrqD+qoR8bxub6vJBT
p+7ZU72PXGNICL7EZUS1j3VRaFG80TtpObGNChKEUegDalgNA7aOouWSm1MZP9iTmQNcGyyWd0EU
2mU0Ij4CldpIjtXuulhwUfT7pPaBjcTHiRn1n1HVcWPqFKnS1iRTexef83JWTWknnFLdCxUNJnSg
oLIm0H/WbmMPRzLnF3RETImVSFzgTe/OQkJs7LGmhCsKRwCbKRKsme8tK2+Y43wlUhAtA3rnNIcw
5Wdub/EklsP5kznUh/XUrxO5IxiD5ZZqRwWBFPe7qO2US6+J5UmQqO0UercT6y8/J9B0/0zJbbFJ
J9ywNEnZGdTiEKJAet7q8dJM1YNn6dfydBGTnDOIb8kvWd+5UNbwT/Vs3YA9tOUx/uixjH87vvPy
7tDxTo9vmtcdZwsYO9OvaR61ClIpMgmoCfTSUigKA8ZFVDCDvn66SbWTFrXeekNPiU0gftw+LQ/w
vkqM0aZgEkZReM0+YuF61KFAKloS6KRqK39bpEOabov66e2f9BffodHc5VXQ2797jEHwU0ylf9qP
9SEZ1qFgMEWhPNptvbz5QViDEuGP5SL0iOgNdUbJ+ngfSrXkvzmrBzi4BPnet5WmAzHzQfuIhjxG
+ZOUA0iYX0DauPgm08IMTgsmjCcADQzMScVAVJ0jBKgUns7h0CyBVWEsbwngBNpM83nhtUxM5Xbg
o1/Gz94VBYTHuz/EbNJqlhRen6KjBPa7+ffT5xFyivIK8NTOs/dKS4bXeZtmKtK95whk4fCcTCiZ
91jixvjgdl7EvE+hAN/qQ3QaCZRhuPnJpn87DCqr7uvpLF9rK8pqQffOX8z2j3DRC0Otl3U/+H78
4mFfbdaK7ALykyv6m+JCKIX7k+sy5tGJyzt0FmG3GGnyY6eNIJ8IzHTY1quPACoGC1j3AtUC+25j
yNY8QGpkOD5Qnz0Hdq+/y+1vohiI4+cFsxiJzEkuMikFoQrBZm8vsQre1nS0lQnGkMs4cEUPaZb8
8YacgtA83ZEuSnDZLSjJGYtMt9MOf0mPqvGoj+fJAafrORm8ngV3yJlXnq19/8KRgHxEofvMieVd
A/Kfg+79VLmMpt5KNSVGb9APMhR9zZcTpyEpvwtBKeNIhtYgGkdpD6l7oiPWKAdAm3+2uaTD61aA
rvMNLZUHwshGL5+dcnQP0ixtzJT84tNbYEW5Z6TUA0ClcFA8Z5hYkYCx+hmLmUMrJ+hQzikEb+ox
RKKdHwzrf17rvmm2OALUXNBa/y+iiiHKD8AiTvTZ5C1XXs2OSAXGfOhY40Prrv3rnbEoua+oUJ0Z
+uHaa/ayuF9P0vdtkDhYIQEx390ipuRhTaYb7XYn25n4Svq2us+XX6zqtCxPjYwOMCq8fe8Mmh9W
ng+xpca012pHyXARsYRHyRu67zlHfbegCpZzN1e1x85i8CUuDNbdBtO9y9xV/GhoJ0e44BQ+b9Qg
9j+JSdlgIdwY85s+Je+/kcM9Fk9yln70f17KMnbGfkIp2vW2SxUwe64UQp9Yx+6sMc2BTWpG8t9y
YvkyoCBZOPie9QUP3sFHy0fJ8e7u3+gBwloKCuNHj1V3CfixY3vEjwp31HFgyI5GLH/Ug70xNRwx
s6fx13XBN7halC8Q+94uEyewvgbuuqtV84Vk7YM+hXmh7GbaeqMboF4cKTcm5/xXDYcrJjzd2Z5S
T7jrmJKwMK/tl+xzbAnTwLeBclpXuhd6NAFBLrAOM5hthKx7gNq2UALjgfVSmLcMxKuBXeuPsEjc
UZHg2a3bDzohg4BXlx977Dcn64PP3Z4iuoPD8m1Uic0RnRItKxZ/tVVwZSedjCPJN05EziLHR73w
XwvGcn6oqGVu39eo75G8XBHqc3KaPivU1t/r7cKZdB6QPk772dPF2JVwSh1o7143u/M5WDGjettj
7JymDMDeFlnqCCrFKgrh7BxlTc4Jy4sOkarm6iXC0yTmBxHryLUB0t843n7BnkTMZq+ZLOfVz3Lm
Gwtx/UvUpruZ9zBBSIe/0d63TyixPWoO1ts/ogvj191Z3Vh/SamWqqNno6pEZbmZQaANNblpiF5A
fGxBMuZFo8xLpWqaj+AW7jo9658iAMgDWwThfB+w+DOSmCQXs3IV6XTEiF/55UDIomhW3hSD7irB
slWIwAZurzTVFofbHlIVExWA9CagXKacRwxafertF1cC8avT5EVBCvcGGcihkm0K6uf1M4uKnFEo
f7Jn6wM4wyt2Dj4HkBcGlNGqYSGdt5YubxxoU3//RAMZq+t+qQx8N8TWURw1pdYc8liK4Vyk+8E9
jb8QoP/WKLOoiGuDpFWbmykYQVis64cyCU3qQlN5aq+NC7bM0jsEPrQ3Qf65y84wVFEHLnz68OCR
ijuVXh3aQybu8FQMNBUAqqgr5V8btSzMyUmjUGeyz8l6JG4VRrLBqHJDvSR/7LJc0kFBvqtvWDb1
RAhIhTP4/Mzz8zsfsK1XB8EI4RyJiVZoFBN8he338PPTx743oiskVvBEwfDKkKABSKP9SNzXmqvr
cNWlY34LykB2aWtAXr7OJiQ1zTAW1+gGUOErY2KjRnm4oiJwSfA/2Ym76WEzXynthYx/e+PySCEU
a+xwYxNfzn5RkIo281GUSoddF9qVxWfK1xVunytUzQ0AF9aEuWZcGsiC4wboFpPHjA5KUQYQGoam
ZR6arfZf7sbE9cWQ02AwWyJjI/ZNxQkc80AtFRXsPBsgoCNzfr4+vENOpiN5KNo6ov8ybdWCuans
nOU4Evfez8dUXYEo8MIr6o4RuBAE0S2S5q46NHSgyFIOiWGwDLvgOrurRNbz+kcste12iDmLl9Cy
U1o+WSmjo4ha18i1zGmzWooqLrjkc2uB/7aHIDwl2L+AopQ/6IxvvJPkiDOqzgauENUdfs/MC9IB
qH0WWgV16vMJ1jPRZOfO528MTbTrTdZXNzXtaWCIRlKXNdtN380GiZcf8uswdukZFnHuWB0IN3e1
sCVyfUXv2BVIOQquQiYr0gtM48pNz2idlxruZq1U3jzTRh74EImvaqXVuZjdnYd3cCRamnRXu41a
8UB2gb7ZO2c4ybqSxkAYTyiVQabdBi8/ob18G6NfQJXJlSvOefmis5D9V0Vxm7TkSz+m/H7cQ0o1
7QP51sQYDlZbSH/wTaCWnB9bGIxMzzi8yCU5ZtdLL2A6xCNRG+p+085O3RVZSwsfzDNEPzrHlr9s
YoheL4o5ZD4hki/Sa+qnEkG9G2iZbua+ZULqjF8xnF9ljL+n45nwCWljMzm+Zg2Y4hGWYtOp3SIW
6zIcAO1YfqGO1QQ9vdknGtrKwG0GzHxAJ4FQ1x23j1qZdQHgl+PmpNPyfvGwmo08hiD81nhKAILH
ol8RXsLAmJ+uU1GVdLPgYQbLuON4eluDdLKcdC8NNK9tm76gSf3jOGp9XCo5udYou4sQq3k2yK39
WYYntkzs2pKrLgz+ywRNLLZW9joJspKEDUkJ77+q0b3cU+ouKFzcX+DvTtWptvygpTbH/Z6po/Qt
k6tuET2voG7zL4Q0jPC6VjCY4IbgCOBgy94jyh8Wb41vPjxNidB2HI/Ax3DvQ0v89u1cxwK5i6Sk
oFzoeUiD6jRsHaTfFpDCRgK2uicanf44rYx6gvCo4N/rULk79a2a7287aDWbID97JGz01czytHJU
Uq4m2W8xiZy65Wa6GB7Qfo5f7oktYqrCFB2ijLeU01paaYH7aT4sTCG6y48mKB7rA90uv+td7vgM
NH9tPaKfBj99wAn5SqJdDirLTUaVqe3McvL6+P8ysPUdVWxA8CaKGMfBKrHAYEVaTr0BMdHYQyqG
8T7SjqutF1vFZGZVz2DqetK75ETrFCYHyCpSnOnoUeCneyuBNbN9BTWnsdnL2wAFJAbCtTqiCYMd
vXabuqGDXVeBmQkjWZTPoI7AwfXvNBeFbaFHwxytpSK1p90jNmYt3FyKoRuovARqCLyOw4FaD0gb
OZ8C5+FiYjxlbvHFlsCaOCSaU4sZOHTTn0Goe8DowKrteAwyWGvf5cE1uCEKq3AxKn1jhCVDAdJF
CZCI9qfJNumpmZD6RN28Tzoy5QtsUp8gw8kVmCY9r9P1vZ+dUtde4M6+3AD7n+mdR2ie3vvhYRyb
L4h/KzjK0lNOOP2xBFCOJ7KaRibQ2wHSy5uOYjujJ2XoMKvpYwp0GuJgkTqb4PrBgNUAYynwLHfD
SW2fZiv/NoHO/J3vyh21oLD8iakoclAKh2qvrAmHGSMGuNZPptT2ptCYvx5LcqQv0As4OmhyqVed
/lZj3/eUcCl/V34Fg/XzgF4Us4WHJvpG8LlpPY3NqeQM6hh82HQ0b3JzHB2x29QhRAs+lyjWa4ZB
+ppA5UT52PPwzGfLVm28gbFJfjZ5W6vmcJrMfkwk7FbQwmp0IChbV2hJQGq3OBN+KCqGytICZ6IK
IRaercOXn0lnnR7czqkjQPUxlHER8GV46wjl9CHmKNO4dFLh6RiTvSYPUiFGHQYWnLYdOHt0nkqH
gKrc1+BGJwQGWvooaoO+JJH+iTIleYwRxSdOPoyWpKQ3ZPL4RNJjCTxZ+y4WMrorpl+OIierJfk9
QrMDBFOxULANkgX1hqTz0c9LriJtiiIihzZFQgqr421EXKjk+wE36+hHnho16XTgkzy+ftm2XSVX
GusIpC6UhAUwEa5BrfzBxJziuEr4DDp5S9aOUqMXkw+ZF1FlOn4aObFOk+97e2btmDDpeoKirXV/
jFmIzswFFiAeblPXx4GOnPgU6QhBHQtFqDoLM00QHpAVm7JPegv4NlNZRDFkUwNz07xTG6R7gSQR
kKWCxcg+MGsKM9BI3EC4tNZxHY5RZ29hz4y8H7X7vd2PnmiVQUu7D+mcdFMPY1KWjo1j3cPkT7Ul
RvXA76CU9rUKLBD4NwlrK/Hlsr6ppceagSdtuvULWd7aUqeUrUiPJyPARJAw4bQAFUIy70wwyG9s
tDwM3AX1u6C71QnI7qLXION7KpgHokXI9NYdO5aiXaHiYtAS6iQQsukm40DltrpMDoBHtC5qzRr8
4JgFcoTPldtTmMR249xNk3vufyWwsHCJWthWUrlMdw6J06znf5eVQeAKMzuOhvXQfNaLmMmCMGNN
Bb/qljae6YrCgiX//sAQIETZHtZrYVIRS7fhh6QEog1cXRofclv219AL7zADu450SWpXITb3YfZg
r8nffKJjIdf7E72GV6umnv8n/9b2yUj8JoNUb3l1g1td9+uDrGpC3kqau6e3fegNEX/N3CMIfyXJ
PbRqbwPSrb2YYvoG9y7epktQenyWuhLRJVDGc3lDsY7c17IEm7zdfmOicrdH4X8ZnmbVKpABpviU
MZAYIYcRANX8FuKcZz7R31Wo2Cck9qQJ1dw8U2VVwpPZttarKHypozaOcqj0dl6jltBH1FUkQBsi
CVJchfmvjb+1J1nYrUEpPbJQw28sKyVJ8O8xRL+Q26m8bpK1HaZqNzP3hKnSf/3D+Es0Url4/4Cj
X1MG1v55UrMNGmGU3YAhDJuWaosUnefoJWoeBdeFHFeACp9Rz0Xdl36IfCSBcAGD8sbV1/W3/sOo
H+F2RpZVLR5ICbos8WQOei3qJ5wFu7CQ+2CCyjPjzyLTQTF6UB/1tURf15DhhrnSN6Fg/0x/0tET
ZvRLvB+kyhuErOnpCCy8D9Hh6vsnKge0PikhK6eiNns8ogWG5erNWnnZru9ZGHJJZcP4cBikZRn/
WkuAvWeypGgiiQnZ1lmvuElSz3VsRC9TtK4jBQRXoqnqoi5CJhNuxRugHKc/Bgd0SyT30vaIRYAY
hkqRN0bdem6bHhTzkFMWJkR04KRjpY30V9X6Y7QMSc0JlJ8ArLBjn/bF7D6vYsK77GQlCkIpdfZZ
gUELEe7ad3C1rTCGpL0+3+q5sU6pOKL59XNdvgNSrzCzbVkfaLKm2coD8BC+mYW3VQR2/3zpsz35
W0CwlgqRkDYy37fPOmsLZBaCaBGM63V0nmt1LOF8AkD1Fs0080lA3ucwT1NJ7iK6QzhzV5VvEzd4
C/59f698O4UwwFiePEKbY78PCalFSjvj9G5cUlaPxR5DE+heIghly+QmUGSS8ZvpFDSnKsDGZynh
ldAK4MqPO8j8S67GPVliymYnhS0Kfy3XHaOUeiziAKAF6lBRZjk2oIl7ifaeYMVS6g9PXUJvVAZT
mxkogQUrrki4e9oppA3FBLdGccTRRcJvEHqfhmCEREbHk40uvVP6C/W6rGjbQ4+iJ/IDiMNlMpZ9
YnlQCBlWglWeaMkn94Xe9MbK2FPMWOSRTCEDUqSDhydQnWU0wZZ9QPj3kCxUgK9ianSrtt0GeGcN
+0G0Z6GJ9rw+V9F/cxHYK/oyUkAgKEFZXvC9Og5qBQ4V6M9D58qzpK6XfX6W1TYj1zUexfu2uC3M
nEjuZG70ZQIIDJWKpBN9x1JjPZyavMhmXjuedCFmW/uqc8mxceM8tVtHG2dExqRJePPHuk+fZ14f
Z7NK0YMEiNbexGYAjPHy7cdLO0q/ogziCZp347v+hn8tP37UNmQDrtDwskvqWfaMpQU6Kt02GTGl
vxhbYAIPN7MrWCVjwqSQYooPtupOB+irAUibsYlab2K6peempTSSV7xCk3wb041+bf+/OPJgbweR
wdya6ZHlE6woWI2+iEC4C3JYfZybjjs5biYOc042d2FwzXGwrBOOvWsUdRUU/QGzjI3Zv3Ql6oay
6ezwTYbVAuC6snD94qXXTgdrM3owk+nXDMscVDgpPsTynHhd7qUc1nOYaT3enW/ee51fWkL0swuZ
qMnbFgthm603xUM8L+Ly7dTHfoVXlJC/2q0UvDmpjaEwet2rJBDV+OkThNFKOhB3VVPtF/vQFVVR
EZz2tQ70klrdbG1yG1v1UJbhHOTnnsuc3rAlE+VeXayGYsevvZfDcWTqlsL8Z1yjWXnuFfgEK1hg
ATQKEnupRF87043X2NQh7bRFl5TjUe39VWoMJxUm6vGCGodrqtgfz79qz0UFjBCWWmASb8yFFxNC
tJRR6O23tvdgcZ0sYyQsE01D+CkGtlh+NoqOQRDBlEt8hB2XksQWckMM+QLA5dwM7k2lB0PKbGwt
pQHpCcXxMJ1/+ZIirtdv3lIgp6WuUOPr+Eb75I60SIZkDI+lCySehHxLnci9kP9pdzOjUfS3dLJh
Pnz7R1Dc/PDaHOXpww0fmC2TdFDEvza5PI1Zfm6l+mj2KLxLzJRMqBEGhSYpJbqntM5BXGY5Of8/
Ystg4/GUkAtI0apgzfT+LVWMWWA0HdX2S3cIS7AfwsZR6jBLkIx/XWzNohkDlbfMpafkgadRxJGs
Og+eB6eu3Dz9DREB2cWYu4uBqJF6KfaM4LaHNqf7hcxPEfEtFy7ix41utPDLH095BraJZgxAYSVb
RVkA7zsgQC6r+od56Bw4BAJ7aWyY864349WwImAhS9iqqNv+6RQTAIuTjXG5MD83FMelUuZWQ0ya
bRqso0PjpTa/RoDGzL+T5Ui7fDQiEXjTQNEyHXVRyjHS5XJxcgbAcdvBBb50E1uyHLxv+jQRAMGp
VpLN2j8f7eII0+NmQ8mEedv+kUSoo2Our81mDkcjht4VX+ptotMBBEMrOs1HX57yvTr2JTD6g1Lg
Zf84ez2iSMdKzljKl8Pej9SZxcxgqJSU9mZUmz6c4Id8WyWtDX6eO+0mZX5j1dHzcLCUb/vD9vIx
yBGiI4uj4txCobKWoLp19CZwElLulsebclltOXQw1rKpucfpOWfw+um6FUwUuvbcLn9EQEZBGzgt
SJylsZ5TwdmpIYaQqS4zi2D7w1i1ZC5Bc5CcAL59+HmA2nuBdP6XobqCIo3PCQVR1x1joRwGSKIa
E3eSFC7n/pnNU+0E26fRQgXvoRP2HOu5GHXoWuupSh5yUF5xpXVDrgrv7ugwIAHs0HFrydDASzMA
Piggb19kjrs5PNQ9BrAmRdHsh7yuV/y4FvzgUwFBB7sC8g51SILuiphcfBL4lgZ3gdpABBjeGia8
G7XgZy+HYnCmP+SYiFE/fsMiIbKVZbncHAqMP9IT8C1uOGDA7Rxby8cKmTNbUOw0+ggkYv2wqsI1
2FnPdRSOZKkgqHnbROazFOgUYFq3PpjgVYhKyLr8uPNzdwswaRyNhjw0X/yEv8LadxELGYsHjS+e
IFfO62kWT5GrbWTxkVoU8/lGBTJ+bEgVcxfwBZJbGlq4fXTryeJ6vxlMBfzh8XVsWXTs16Wug12s
qmHoaP1brvs5WfNG3sCiHNmFoUx/n/ZpmPPiLybWfJb2QsC8Mg1b/QNcO2ek5pJTb8YseiCoo/1O
jFa3yJ2ccUnXPRY3MNP8XApxqUVNwdUWbH6Y0mqjpkGoEGiS9mip/VzWcx9DQr+nn+tIc6AuCQer
xVKTqKe+FdIwjzDVzI7OIALgGxTv76mJik65GLqXeP2a5XpfyQiTlOs5jKDf8QbTJb7cYujKKobV
Lj/4EG5L0qvtuRUWhRFrkuLPbjp6aak3BVdimnwNbagnKV+QyPrSSEy2wTyHia5ahQIo362rlXi5
PaQd3ZKl76LLe7bZXH1YEF/JVBaF6mz48SRRd8LqO0DorbRivJ/BmIxS3aOCLvqPkDqR1AUZIuQD
fR3y9uEMRuRRimLPe6LY5BZrC5oMNybBhrk7bcyCkiSvp4GQlxgA+7sUw0uLF8ahc0zjYDHVUh5l
j7hgzycR3BW6/F8Y9tAr10WKkWGWNSqNBW+rLCsoBo7Xhhx8rDa6NRk0mE3xXAmxP6A0CjjxOyIA
Ngds5SE4/JLWeTWcVOIzs97E/pZ40g10wSw4OhLAAtTnyA+vbuGoDjd9dBPXEfPRBjmsb8PF3VP/
Hoog103TRsN+zKP3T4gp8FR0gphJdyaVQfiQnfYWfQB/uszaze17TLJvDmuEe0wQug0n5VQJ4rwI
fD+dflXxWHWbnHCCFOLXVBD2wRNweag/+FTH5Y58/CUjosnzdo0TT+A6IPJuAn6eHYBj3VvNOO+m
cuz0Ez7PAEV79+apKVMj4U/7bvqHyn40mAZZx6ht/F41LMiYv0EQMTVaRv/mDJPurLGRkh9KPRXZ
U9dnVN8HLvx7rQL6qZNpALtaukKCnu7vlanThFRYYpI5AyYKpEj3P7k0dTGiCV7mUrxjxtnkw/25
Y06pl/K7iLn6uX5rT+A+YAl9naB4I87nA+NrnbcdhWeGYef8STrlU7w17lxxgnQSMn4dbJ4F+UU8
+cWhQOG1iaQEYqf5ZQgLCOUJpqoDKMlqNuf/pOYUroXl3Y5uGFvKZNdx6xKwD4HRPO1Z9YvdZrj5
8Se3FWZqE/sdFpP/lGI4LywCzsHjOoHZ9nbrrMBlR7BE02ovXlMUaMrHGK7wZZ/aD6NZGUgkWppS
UgqBkAUYNyIRWuUFbzFKh2F9SPqK52Z4vGGyX/fg5J90VnXFsokOzNMbaK+w7qkyvRx39itpUXSE
vkscJSfbVV3gm70iV+0q6cbVDPBBgRMGgcMkfqVX69fHr1r4ccTQDLi5X3tTUIQFMVKgbOk7+qMy
qHu3IOuRPFTpZhnF+2p/yohaadE5OOBb0142BkrZq7FMWIo2rMw/xp+K58lYmYHXiVayF8cex4FO
PBOj06a4sqgNgBBfxQHtN06pvCxl6SBzn1PGzRbgLRP+MPG6BlihfRUqsr/xrPdZa4hMz6CsEnHn
zOw1Rv28k2B91bgSZb5vf98mSsACZRvoXMuJEnmATHVtzvNbtk177qm81Knbvy+vLgZqy5V5vGAD
fPsN8ZvjQ1LedBxvpMM4MIMDTUkH5q9hrXH95tMQazmwcZmzfx6FjAme6w+tPVrDuyJuyCgvzdOE
s4317wC24ZCP4G7zIaoQYG+UZ3Hfiv8VSRU6UOGMeKlRLF6Lf2HAEiBic6wuDfG98J3ZCmZJ/WtY
Ov+sk2SQRWR1I50UShkpKEogK4ov4lmJ9vPTv7jKYaMB8GSI1RmOYlMHzc1TtpWPL8zLItcXDYhs
EIgyZKvsy9WON4ybl5PzbwDYWQ7x5Gr6dEm5Gy0CgIRWC2zhQY2+DQ9yfX5apyTFOjw32XSIRxSZ
Nefo5PeTtAz2f4pCT0pyFoMpLE2xGHxbGzDDUlut0sGrZlvw1if/f7qZeYdgqA5xO4QWVIW4b3mI
y1zBluBsYQXO94pcQpGsuLsqkvmwFMb9GIfz99knR3uVcIVchPh/+PxXhjCzyEmSHexMGCcR8l3c
ugkehetCs8nrgV54VPThN1WJkgoMDr0z8dPKPaAzYcl711sDZxEo26+FYeIUHjDsYLet58I/OJ4b
QrS99Fd1YokjsORyIkm5w8nePQyLA0pFdgfLQbR1S/QcD5y2bIWnmVOBkS89j2IZHZnen9ANzuFn
C2ORnx52B9Xg0Ma/r+JFoqAEAoJ6+n8eD5ZoVPN43Fza0lljkVpOzoRCEaxvOZN5H9KVR5LWFpaW
SnbceRDHpArSU9DT04lFfXbR1P6LY0VrZOkUnKlIEHIzuh3p1FLecWbkMYi2laCyvu2OFbRDDge3
h7m8USi4MLv8snwPbLQO2Uk7W9rEmuvjJuValab6AX8qKiIGhu/dz4BaRaJzOIMNTSycewalOlQ8
fz7zwd/bcEnVKwaVXyC8M8B99pSHWvfUM/PNj4ZO7lGglForjU0U0pNRnP96WsgDX7NambzZLZfj
ltKgEced2caiRKUhyTanhtYaauOZOLnpEmXVPJ39DdJOtG/dOQcXwj6HjTtBobtSgWMVZSfWgP+b
usuEmPwavrrUVBXwEXGx8MQbdRvicz9+HMUzziEmKmGAQHOPj+N3ywTvwgmri054g3quDJdT/4AT
fKftWVTma50wX6ZyMAMc89vT7+g/Z/j/7bEsPZYHgGMltUcgKa9U/XrRWwWZeo8eyg2K0oSpFPyp
R0XJhdDxrj8tWBs/PHokymssQku6GCzP7L21rUcCRCj6G000i493IIkLegTuf0St4ZSP+LTgQlum
UbMUqdyIWohHOJU6M5rXmDNYY2zu50saCqyEJC9sH6PwRjy652iZha2Xcmyd9R8vZTiTvCj4fZ/5
af2S04N3Y3zO7UEMpOK5q9jeueBl9/trOaB2F8tFggfkoZ42M9ptbZypM+HdFo5YXK2RMTyKLym7
4QH9u3RTwMdAm8ne/dI8yJWTHhQqrcwJJxNX3sDeEupBi913ue537ZXZQMJ7wi+khCbrz/MzGrz9
ynmt9N4QLniWIsHOsM9LkDL6bQW2LsXjGJuFF4PkBR5dkP4RVSk+wr0BiqM63lgPkaD/YQDNe4Js
XDVNHiwD7BhTlu/36aAl+WWZuTLvO1E7enxKIkSw/ei/3m70HJtj1mKVU/bZty/91Xdk+s7+yKa+
jNlSKCoAjz+yWSEA29I6oWHZtXwQpoDKxq3cUAca9cjabgBlyxKSv/FMmczZkrSXHTjbZhRxEpck
5WN5ofc/WJ/qVwKYFeW/rHOI+tStADhhMKydrTTGYxUBPLkj4OJHoeDH0uX3QCZFq/x5uAQr/wGG
iYzxfhHqd6S0JvP0CLdTNS9+TxZav2eYFIpZmV+/j3i2gazcJwgAOJgUlz34Uuh2tiWLUm8ybCQz
d3fYd4npx2FpatYPxLBoSzRXcLxLnPOaYpghMQyvj9R1WJe0yEIfme22L80cy+T6qRCf9bK5WflC
u5U1AtLkieaDwC7gsoORC0zLqtUqjk8d/g2JfCNKB6DcOpGhTt+EgHKVY8wIxeHBKF3wC9sBebNW
+baPyvyyxN4kFtYseN+7mqbiKHDNcViAKt6EYnzuWx6jSqrKseCHMwKxIjuHzAHXnFXmknn+JVjx
DZ6KietEMO8r7UfBzBm7ZtMmX88wnsRjuTdKjPrMBmAMQgOFE2wF9+es0VWsJWsV+HTTjFE7MqUL
otPIasXyvEDd1ba6kw13g04QQcW7mIVJ10JK+DVtRN5dReZKAA8qW14vwoC3mPFsi20Zok7vSZEd
IalXv8Ayltoo2HpWpGDeUw3Iavq0kabxzU+xBpa++uDPR9wqxTjj0swhllCh8Ux44iUK5leHYS8j
xj8MIvw5X19OKVEeDm5bRYeB2jJGJboAhMluJvWv1S1wpFTEzhi1TvSXqjP1vlZuI8YaMcgm9UjD
D6TdZ8YY0zOxSDpqg54qGYtBdLLjh+Mwwj8rpBFk609tr0Tz4A9DJdSYcLkO6ZPsFflW9G3Z0h7R
poClnByztOvZiNbQ/uumqQ8sJ95mcAm6/cOJxj4KY1H+Ael1Ij50Dy5CAKMlF4Uh0asusUl8kNnE
c8hK38mo8uRBxbVeR/aheW0w7KhyMx0JF3yoPv+VsMJ4lt3qST7NKscvcQdXmbQYMXUfNphzz0Hd
+pfFOE3xfAsMQngsGns1R+cpheXvwEgK44vYKSfCf6DqyVK37zezNlw46DODlyzh8N6gRKG7kowf
6nIgxe+cnTivIZiZviEvMcARHNdxd1k3BpcQJmWz8rQJXMi/7D7POL8EbexXIGJEk9v0HsZEa22/
yckYg3/D1xaIooh6M0qtgDvdcRZtfZQD3RCYVKqiIZVIy5e4IEjOhjco2nEL3d3pv/Bo6uv1BCRo
Wxn9tL0dJDnrABUEuJEAvru6MRSEKp341qax3he6xFlseeOYhZIjkrOZpYkFDhcLttXi1HX2TnYK
0jX0nJSpNXclAGn1KUYQOeRKNuN0zhXrpOSrjYmZkNNPnZgASyhPsvlVGmeo3vwmtLygUpB+7D9x
J6WfYm454HsGgzEE6SZPzFnK3d2bddnLmqjOhV2sH/X95xRuh13jAyRkPYSDOtX2JQvgg2B9HxY0
0sBjow59avYVRZfRtqAgpulbBvh811CMiat+HsACnZVxtyXv0H6cNzt6hgCLMlxH5bnsyvtW1WFZ
roGD6sHIPV2g2/LBhqORAGVs19+Lcm3iQJeQZT29iMV8oYwHyvTqLZU6FX470ZMzGFDr1kBMzYom
X1MqYQGBGA+Oa+K7sjlfP5yg2k0Zv75vKcCv6xPhb61mfRyzGkGB46Faet9exvLsKYIkVPZjDXfE
ewvX+CTyaDkTcfzHGl8nN+7qowz94y5GM9AdjajhzAv0oPIFrJeGByAhci9u2CB3ykm8QfiHYbPl
ZQIjl6xdOi0+I5aXrp8/NFEUSKHQrKx1VVR30NEsSmQ9lV42HxyUzE2vivZuffYRrki7XS+h+T4n
YBdyk4uJegKN8uV5wle3PLFAECviXFh4PpEB2ySWrwWbP/WIFjYBXvVqp4CYEUIhvQBETd9Ru9Fh
komebT9huj1sYHNnSzBAQm2YGABPneV3SWeFTKwiZz/6O+HbnolEPhwzPVKOx3uHUSujBHy02/Ib
7LB7PoMxzMGj8sL09s+mcqycWBq06pIqH4lv4nEBsjaXPhWNe/JfyT7+vwejaRB/4XbQRBR6trtf
XJsgtfR+DL7dGzNNE40uU/8Lc/ehOiWkNYfa+7puy/HitoutQBSTix2/Z+0sBJPVdJid0GW8/ctM
ieqgCYMfzRvAsoOPayva5Kq8LTAelSt/9K1/rcsZrJBpssJ+2PTAXoYaAOOGf4oh4YQgjiircsNV
ZvdwG16zUKJPKpGeWP7dCjIIXTxoLkdb8FZUgqFSbMFT/Q2skq0Ia/M1ZU8qg/uAdmhyvl1TA1Bv
SigicaTk6IM8ssOpDi3hKU+JHEljrKePRHVrl+L9fpRQ3cErSpvn26EVX5YG6WkIjtuCVxUPbDby
R6gBY224WzKw0LxSw5lzSGHhzbwB6i96V//Txrr56nKR9Bx7eT6FFpbK8bRQ0bsbLmWECFZr5txi
HiNfpZgAyBlp6N/9STD9HMbhMTjyfMJl4FquWfqB6m3rcZZK+qK4HtzPwilT5xHpLJECYcPtPkSg
B0UrR4RtTceFL0ATIOE6rFQCg91l2l9Pio4xUd0FeQuw9sXMRP6n4fvkyajiSVFEQ7UBiIQsmaSR
NENJ7TT63Ks7922t/1XqQgevzNpkPbteyCiJkltdbHszxsPWE7r+IDeZuYs7cxALAshtX5zWlhCA
wc/E5Hr0iDnn0Hcn121CLpajHz42UkGeWVvMhW3kk+ftt2I5T+V/zdf/y4ogphidz+9SKcnAZNiI
9+poBLTpdca70EjRqQJVypi8lkYC0wFS9iLeQHWccAWB+/8oOLYBhzXszC4dbq3ilLe8LB/hIyPu
a7LIIdzeLK7YBVbKlK2dUmIk2+EvOc84/3Jg7Qzdpwlzn1F27iTdWGfulqWpQVr4vYxIqsPKUQqA
zNR9uDH0TMLB4HrWzwrnel2Uwksasih9xcIHpve2W4n90Dng4eZoIha+xjT0uE/RPV7dviF9PaC0
MZ1UbDTwCWzs7+QNDAMksjcTNzHD1zjF1XbDsE1bgz7Sol21E3Dl4va+XE0jWnss5JX5SMaYLOvE
X5OBHUaVZmdJQqKJ8mBfA9DBqIW9xYoSO10vM0b7hwyK+ud+Pi04Xj9c/96UaRlXoESeiEpvn5nq
m9QSW6UKD3kBryO7VJD0TFiTo+b2CrmGNAx9vb7moehhsxVhSbOvNYfBPm8jd4iR6GqL/rLEs7uU
29lH2WZG/FiZDlWxlPHeG0fhRderrmTB9+Z4QPYjV9CUZUQqz3h6a+q2w0m4HFEsqda/MoH+Qm5I
566NMk1GjhQH6Ms7tYUKSbT02eD5T/8H2e/vjmY4b1AMtFdxf8xTWM7rsKqnIJlpuBmI7BDgVG+O
DWubSDoiSk6asxt8SRrQKiQZDpV/QDcbipC8J1+u1wjPLgcBdN3p9ATu46Bju1CMPopIAfnHREEt
nh9cAe6CA5j/iaepTyBf9L0RLWQWt3MLiFHYUfmEa4N33tZk/LpDxEjJJ4hFg+TQwBfXu1lq9l2t
DLmhw/Hq1+GHyjNQToLOOuRrgq3iQurC/hcXeek4Oa1mFNQtvXICnho/LeQgwIev4xQKNWiuhSZI
38PozIzwXgSyCeH1o5vtGUWUvftUKr0K4TClWvmUpRSO+Dh5++C2puEFiq1DcpnDjFgQGb8TEDGg
YY3L5DeIuw+HfvrGiQbcw50abV/BdANhzgzPT7P8T2hRKOpGHhT5rm6s1itOsol/Aio0rdWHQjIQ
+CPf6brf6F2ABgpAPBZUt+LUEWeeyi9cCW6iVyHoIDC0/R84+tTlBJgUT7h5vG7J0anMcV3MvTWP
7+0BXEms/mdzldO5loNPhKI3/sWWfpdDd9lUdfSMhz0FnQcchqBBC48oFm5khQWAXNrA/2PNRZd1
ZXtAWES7TTb9JUpzpTQTAlLpVUFPnP91OKETroiDw0c3t72z/vj8jP8FvxPBgoxED1mp2NIw2kBa
qmZibjsThJN5tlFO1hgkFh1Ber4LmZBYmA6F77ynwlHV2DDzq6NZo8rxQpF/xOYbbBueSXmmriME
6e5tf3jryUOqxJmsnFN9QgkiA+bcppN30zP8jHnFz+37gi3QO9SC2O1TpJsK2WzuurQUsyCiFHb/
1Qj7Joty7Ik7ejD2r2TSK10UH8PHtDNZVfE8gWyPiWANfBmtbHprzkPbG/od0ukBa6swz3WlkiJI
t778pEjfPIaO+BY0BmInTg3Xer0Zz0fTuHsof5Vh8evRdQxmXOCkAZPTuO4z8iOxcCpcghKPkBmQ
o1YCVGxX6CCmLJo1sskvniwpSRJ4NCHbQn3K5NXG6BNN+MwLTGMGFhmFnH+svhASqxQDkoqrWvPP
CJ7qXW4dvQZIOQQ2UqRIvYYj1EBwe62/0orpmsPW056QGwrrhrEWAJsATbol2tl6rmLV3vlstRZL
fAW91KGNJLYFlWLEwFiMIeTEaKpHsYIq8TbWeBVyMcOYNWNvzWCJv6nHsUlGoNhz0O5XsCZdjhhF
/o9yqVJ23pkF6uBFpf9Y5Rj3se0NQWU0W78nYBoR2bW95vP+Agf+yzfhTyNMzTjYXzoqUN0mxxHH
MnsDAIM78HiraQNmCDD/rm9Dt9wY86jjoSBF8q4tpJoNRFk4C11baGN7fk6F9XIJOSY2jkedTihG
ZWyqAgSMUabZuMebpaKRP/ZXsIC4HLfcuYhAvLS6sWXszPjnrikF/ccUFVCYCRPJDxea6sb9VSG4
7+rhXUwRUZi1b3g4T8tvqMUeP5JanK2fJBH9W1ntwI5d5D3WOUYC3sgEbEL5tDuV9QExYLNCVTa/
aZkKTPCnhgQiDRD+JRSuv8cKlQeLJm75JeY2OCc90/EpUG9flM4eyVvQFQjjwR9Eg5MD73eEj5aF
CikHIxQ03aemiZyqTrHI+gJUIZ3dW+qy1Bx4R2yTe6/MathsCFgf7R+pGNnh8QmS2jZ9oLSlf3TS
UYfeR0s2+fZoF4y4eYNi+7pEyOBGU+iN2nQxtarq5N8yNDLYt5IG6/ZpR4XOkUGvg6srnBmqxQrL
HpefOabnOsFTB9/hXKLCXf8/hb0og5bEYp3470MuhEIeyMGW4whnJ9y49smyZGis47KYfIv7x3MY
rip36bBzdI1qKKB5SurpJaY7fFzjIzGxK5uoCk04aP7ALleUpnRtmPOZ2NnuOyiQ88nEXExpMxhQ
0S8lKssxqKkTyz6pFEfhfuIJrf3alsNL9RYZ2CKZDK8S2nTLArHd5D2t4uCdS9p4+/6xRxCHRprk
EycwsEqgH3+5ddo9O+UMsFnqVnsOCYVh29ZnfFRGvGQpr6Ja4Hup90Qz/0zlFWHrRG2/DHG884cz
AbrG2NlTNOOWeVmSzygKALwbzl6ysHLiEEFtviin9AB2yiNwFOVNW4ZJegn0yOQ+CwRRLp89XCMf
h5p5mUtBCpkg5Y1ktsmDgIsoVAsu2V9nEy8z/xSq4e45eZUowEogJZWM2U7azpUlaCSftcwTdmk5
KAXAlRlxZxFT4j2+9Vgce12+RU8gpFk+d7RJMiv+ntr/isNNFbYNHJNpMtdlNtK5IO/lrAHD+Na0
L9xHx6otNvi56wu7Vae81NjEWHqrt2GCKldIHtBzOkeTiU0t3k74j4djDAQnitwtHNEDqZ9GGwq7
OfpULpfmq2b+AmOlMQlkFN8lKOBHIE6MbZrW/3jLh0Ux1NXMoYtHdm3j9mv/7Sr9zt+DsIy2AWv4
52qyIxA39O14gn+AHd89IAZpzbEC1026oHVgH1ltAr0PjXPAW8duimAtf6VNhj+0rfSE7CndIAj7
8+SEPrYFX3aMwuQE43vF4q+BXQQ+1CBwbKkh+B4iMlkUkKFF1x5TpCUdoi3bSOfeheR1HtlGqKuu
39mkMXI9P6wZEzflqoY3GbS04MK9cnT5IyOSjAuuDRArhWJgk2uUXcca+78UIfsaz0PEQnPJQWgp
ibA8sAg1BlH7JzA3sxRij+04qcikOCnhwHqqsp4CPoqFD8hbWk7X3QrO08DA4ETQzqEhBOpYTTLe
qjWvItdJraStN8raE97V3oYzp2UlM9ZbcaZ1OVAn7Rd4/T0o4VN3YEZTsGiTNSNijNDO1wMYOhAk
32axI9As0VzuJojPXecurNUvIJ932J2d3XeTThzOhjob0lNzcXTWUGzFauXepKGLkEldXaB1PA1C
468lXTSbUOWGpYVY1228gZpwIBvJ1AAkjXSODTFKTWXEElkj4CQNz842vMcwjBjVE6a9Az4E86/k
zvkPpdL2/mO2RJO/HkP5FzC9JFEWrMqBHBdmBX5fN4gOKUg2zw12cwz8ZHnhfvSswTz7oMpzrFj6
GdNwmGjBqEsCJYrhsbCfg23v4vpH0xwp7xiZG0os5FlGeqPcduFbUt2VtOJOJnklVSJ9ua/7KXzj
qP2NJqHOTcu6LdqQeSc7zOoNSKlMva1/XFciREtwZHPCiivFLCwY6LiidM0GRlPTzaAGlb7udgeb
OizNL5uW1ZsRIvvch+xkR9NS+MfHbzJT+VnZc/LMsucteePNGtiXNTEYaJAAXUPLj1osqFkkZ4vw
zVv33TNYLMcDpcoIOAYvMi0AQXAJzEisx8SoaGs6jsBiz+nTTolik0F+7mNN0PsMSNtFxzk6rWUQ
ad4n9EY0sq4TzRhAeqBjql3ObgforS0VmEMFNo4AQTAz7v4BgeF/6jX/8R9ZTOs0wLQUnY4DGe0F
ZamrwwnBmhB0sLbJ2+euY/it4SRd6LnoDQqb7KWE6l0w+ojLwUzjErBjj8mPYS7mFZZarzom4ZfT
gg3AsT2BAex1MMZpNeIXbKmyfJk5DU4knThxFcYSde6KE1X2GYub1CoK7OyM5e/+BsEAG1ZB6wFe
23RDSKp/XFx00yCqTJnOwV49jm5TVXj1cKMFBrhl/XhDMFQGPPxS4BRvSiPIcJIDnM9RhALRtqA7
bjANoHJHnhcXbZ9J7BINew8BbdCTYNRohAoJkyLnKZNVJ5qsmz7BP5VAnNRkOLBVS6wra/F8/0+f
Wg8X1h3ir9AC6hVFUKP1nbeEqUleAI3ckkHI+gl7Ws5I7a9FQK0djKgTcPzfxNTWoedNQvAboUxC
OMiWSrudzHm+aU+BeVRa34ESQQYpw42kiiYgZig+1Rp9yZ6N3EYckdVR4KLipfKjUpyEmD7vgFBH
iRuI4NQ289GLhekugcnZz6XlFoWopd6mY2fjwPOY4cRXCfEVJZo/3U+BdV+TRj+MNa3cjlxZUrQL
Q7OI31g+pb0kJxoFIlTE7uAyJz+WBcq6bkiD6jNVls2gN6KPDO/v2ZSnL9s+vo+HVT1pHfVFKm/T
8Pgok65Zt/1jFdIErw3//OUmq3SdESquKh4cWMIyOye3olOb30GnoGaqGBwDUpVLZQmHBPkFw7qk
SkRZ6rqavbwWZV4ckXT5TuAS1qc+rD71jqygXAvhSLzFfMmBqu+OVUF2E8L+6sbHBtIuM2R+m0jb
XlybG9LpGaWCJYtZQW2tylT896RpKiUnzrO16gKFKg8cbvp2YR5BpwNZ5bJy9g5C029Js3KDAOGK
XDIMAAP5ixdvJvLs8wlhdGLJXoMvGxruaHBOZ59P6yRUbGhanh7GUYVXCcCSFvnWCbKi7qfOqDC3
joPr4mmbgEchifjhYenxQQOlSi7CHckHm9mZqeqhLgyrVeWLPyws2S1LdH2aW0q/olXQJrzBiWXj
B4HIKXEFwkocvu4zK3yB67KsBzTXlUCqkWueJnTqTP1bl4gqKsDedk6kOyD1aGicGnO+ZYBfGwjA
83XhiVUm7jHfHK2WJcp/DPK0O8W/3ssqk0WJktI1YSYLZvvyxV30hroOyBfkoudfy4Q6caFbHdoS
QzF1nA9c0ijLy5d3gELBCerH5SfiSgKuhyrbCT4+q67UjTdTEHz6M5v5ppc18J+d4vBeatnZ3xtN
AojncEcMXuHAWB0sLX/S0uDcj/2jlBHIC1C1AomshDHR8J0UqwFN/UFzzYTwlN/OaqIDht9wd8B8
f7rX3847UZKoEbZaKKLtd6MTCPYP7SzKbrXfW/aqG39G72kDbYCAx2zlcxdZZr0YGki7cT6Q0zAW
Xzy/Nr0nyr+2IgQmxRSYyg4KRXeuqlOJJe/tWoYl7cyAGP3yDbtF/54Q+dRgXSo0T9Wh3G8hH1WQ
Tz+TfGFLliprpd9ORpI3NgJ6jPHlGcjKA/gis5TFEwe2Ad2aTyYJ0iA9TpONohKlcR1gmXOIs2uG
socmivukUXUwD7eVGY4LkfqNabX/WieH07zJG7lBIkzp5yFU0mb5ecj7SP8OBHLgQWjzQycHnnjK
xO66xjxwtO69vUb6im3Y8lfBt5cxZo5yxrEC/o5d2nFGRkAxEQTCLBD4XCiFE2XCbtafw6JzE36Y
EYMt+QyPIFjU0rwG26wMu+2hciErDzRVak+uR/DnsIQkJpdlv6ROz2geYpJqWnsJcmo3nCYxJLnk
fwif28Jp97v+tU4TVmDeftb8KQplZPihNjwS+nameJTNMUl/D+NV05C7uP7v/IVrb9ilsF2YkYEZ
OCrsthwuV94qcrHNNCAVsYCSP+VfCkDnSCtn3I03Iyka64EkuBnLyXRbmJkOVnU3yC8w6AvWKNqt
oaDeYIir6nNa54cEfOCfo1NX+9YEbhRbe/fl2mwCR9IO3oYxfBhgeZWF7+OtZVrJDelsev+IiLTY
O9lr5CrA2Uro5fWG+zLeqh8AL3KW3KskvnLn3OVwg1wxj6RfiJnwPVytjdho14RHUVI97U/uaVac
4DeK4yOvqvxkNwgvsLDLzms1lhDtq4yvo5TwlhWD7aZ2UNakONno6Fr7la58C3u9opSETUOrTlA6
QSUFX3YpCc721kpd8l3Ma0looFu2T26UnZuukzhK+ei1eLj9zCWC1+99YzyNzMdPUv0dWMVAq5UL
9YNVC6a+1USyNoMQ0Tzo6EdqUQ3epoJlTAcqAc4TeJQjEBzlK3P+zPyj+xSVKtGpXR+FuEkuWsvD
Q/D4p2oRwh+z2ufq5HqpYOWELI9ebmTbOJbz4B3EXi7jGcZXJvGkS7Thwy7R99fkWpDZzZfsoJHb
amOIg89POaqkivMi1MeGxQdl3E1V0gBRvzm2HtCZqY4M78WKCjYQf6BORFP2ROBhkdhYhLL804m1
O5EGqMnBc615x6mDBRehyVaIxNnDxrWPSgS99+oWFfGmJR6FkJI1lm35Pum9xnLfE7/RImUzqshw
gLqCJ47nqy2yrsrQ48uK9vxtxUaktlCqBgtjtI0WiG0cMbT+d66VEpgybHtjWDNV9nR2KYx8CDeA
zHwdVZB8fzoWKX8OmNJ1LjW5toTm5QknKuotWKUowRvuw1QZe4J6oOWEtloESkUV+OQYhVFzhiFK
ci32QgBCPVGELl/Nki9luPeAcK1DoJ1cVdp46a7FexDbdItaEQ3cm653g5gpk3p3WXA7v7nka5ZQ
A5lEE7ptGpNDHQf/QzG7T/vMAjXhHpbClI/EnC1QTXY+3uMNh5LTqBWwZouFfuD/uS+a/WdOdi5d
x3GNX0cgWrovV7L7aFURgfiEK7hfgJgQuN8jhvztlxjgmPWla5zwcli6YNc+RGEQkw2huBPioGZS
D0+zxbs+/IzkzcMutiYgbFqezw1MdxxOCxnN8zbZDgclTvf4BLUlERpgtGQkbBRdmLorlsXFuPxF
4EKr21/QaiJv6225xLsXLVfxYH8q6dSsUYtIg+KH2OfRZpTEUWiBodm3ABJ2cM0cLkZZgVV5Y0sG
gEv61bRbSTp5QAx+tpvbROYiZ0cZ14BCAYhZExz21MFE6GKBo3BhmWZAvLK7imuTYHrSLyqwFf1p
hV/PkIcRDE2YZaTJgt+5oAI4RDS/HRtK2bwD6dhCjPeVlCJklLZmbrF5vgJPzdKS9gvudYuGYPdl
T3WMrTEabJsTpVJusgPTH44C9XuOnl7zuVy22mRfTloAuzGEBA2DPaihUjoLYiJfe813SzDxaH4O
P5LfLUfJXhdBVjtSVGZ1eXbVnknhYzTnh6q4MM2lbyODc5AhBzD+Vf+wigiBzElY5sb/J69SdnJa
BHpuVgvfUGKTkWLizYcTcvspGx/xOTLkUAow7iPZiCGRd/x/9B84iTCu89juYBEtIj+z3CC7pcl9
w2ZmxxgEEAKjESldoJtlesHN3SIXC9M0qZ55ABdSbHz79MhPrbf+Un+48R70C3TcKrhNy1ppZCQD
gz0Zuy7NS8zdrmp4LcR/hIF2TUI0hxT5K4lzTZtA4AMkitV7EbwNW51z8w6N+ICjvZYYgKLJPLmp
ZVMI4WiMDYVDpNDBOlQWsXq9uBVh+YglLPeHDDyINVVeDRVOXrJNa2aZN56+5I1hUBq2mIUZdF8U
D9qND0cy71Fpco4fD+EfY4+vPcHoC1L6sa4O8zBo6nwNCI3dPmV4ND7UdB8XlhVcSz7UQ7kBR7IY
bdhS9d8cGgfW1rTeG+xfKqHL+w7MFh8Ub89QrX2ekyYWEOpgQ3ful5JxnevFPju0yoWwlO9EZmCZ
KAPTvowN44XIMAU0EHzyo2QlqEEf5p1nxz2Zo0YCtYD81ewk4+Ssywvjfzy4LW73XfmfOe5+cfAy
Seeamw9gXe+IeE+n2EF3nBFiSfXXOtAN3CjCELZ4SgKKlPArAb5LjW2SGh6TGgOjVATn4xS99t8M
+NxvhjxFtXjw5S4uC1kB5WRbnSIwNbJ+7qTDsj1hn0jReO9s/LnvoR8f19RK/7mOAt+kdDXQ31A2
/1hqR1aImZ2E/FWpQSKAMDlrABVPleu3/DOZ286l2W8KOCk4toJajAnNJLs9V/WJvRm9PvwsRddi
Eyd6zS54m8fqkYSCpHtOA9kpfrcoA0xZsBJApu3kBr4MDBgiYpcjbD+rmZAy7urDwAlF/f+Y/LvP
t2miKDeG0ymklZgiR7iQT2kLqKVnRgf4f/JBEiWS25vR0d1ncqNqdNtXouqPXK/xGBxInihXk+sD
WsZNr6qT7VWBtEn/JgVKzZVxUhTbMgjFA4vcWkCajB/i9Yz3dgm5Od0dApwh4gE8+GvlYXVcNLt4
HFAVw12/i5C3jVPKqdRNmkov4klR0ScbBTPyes9SJBkPqh8iBypZHdOBOW+Ee+lMG7xjHx6TIYOC
wrqPN7r5v2lICxlSns8OYsLj6yfOHVl09ji6rZs9CX11f2gSPmR3w0UUrZuPP+dXX3OPy/HrBbkg
qjK4F+GiuChTOa/bx5EwvqgEolDZEvU+G5MQXmlgrDwyogwyK77J5+yTsSke0sL1SqjISz8iZ9Wr
VW7ANRTDYVBt+CnQXsrR8iq2djU8eelEXiEphNmuonwBhb0/3GpJg7comvI7KFOay78FrCsywznT
pjYDdEGugtAuuRuL9DIjF2VHkXlt/v4dak0qkJVZ8mldrvQt3kEMTeWFfEQwA/ssn7m00BURSPVS
N6IOfgSWdCMNW7lOoIDMJHX1t/WPCZZaoYuSJZq0kIsGf9m/7uOPsAg6ByEBwyduXTrnVb9IfFWq
xszaz9OCbxonVaOcQUjMOWY95zGdkS//tzxSy4dWpx81TwKKXa2lJ6rZPcHenK3gDQybjL6qkLKm
fYpYLaa+1e/xJyTLnhhd5hwIc6ElbTX3JVNLFbLHXnqGSZF7sCAr2uij3kIks7pp8BVw+gKi3nEe
KoTtkD7l08EJqaTk6Om/ZjyZUUZvLVRReNZV0lmIIkMxqzaEtQeEM7CwLaP3XAf6gNXFqv6yvuzG
1gzPBSGsRwRJWgxsqUwtTvPuuIPMR6uLMyE98IKOlzkoWwYcoox91b5LYGtSxJT6cs9y47oDP4ab
OsIF8uU8tU+oEdpQrOs0pidMErSUSmB7dtRQVLqgO6KVzdcStLfjU4xRLozh/z7mVv6NyXW4AIuR
CHYXTANboYInDJ+29fjmsqDzk/zJTjiCdV6ae6tdmOaqLuM0s7UwEfJ8mrr3+hIDSoKMCcX/ul81
lWhxEAZG2NDEH3+3o/0SlYB4hziWPXEcWJ5BsV7zjmhPnSalZwup6EMCaxV+3ON59tQy0VHrmEHh
glz5J1B8SbyoyXtK8Pva/Z/s0CKu8NdxB2RpS4lMUrlfdaHoj/HS8JL2ATmz/dMi+8zAK+is1Hhv
hyCR/qgMEO8HnqZC2wqhNtuNWjN5O7DgPgl6T/yQChO7g0Rqoa1LAekDzL6qrZl3y3HawyCcBp+R
UakI+yqzTog3ZQbfrvt/NwA0sB9kNfh2q6+q6q5wnmwTOnybdXgQu3KA1+mDlfty4oZuU4bc1XsM
fHyNkHmQrU2S01rOcxkE9/X6l+a4qJWKUzczwUdqCHzqWpVb3kEJKn3wGLBmsw3sWQlp7X5qcDYN
EEa5l/FztuVQuGFX/kjqtMJS36g5VH7PxSxQfY6B4bJOC6wgjE13clqz2VNpUiAPTXyPU0/nU0d6
mz4xgHqwFSAeVjxhpo8qvCQO0iCU2YTi2mGymuYvEeectM2ASDSZ6Ri4zGvjOOcPQhvfSOPb295p
IL75IyPOXU3KzZNnid9Ns+qOOhV8tIAMmffVhkiyvGDoTOdqU17hlflkKeS9AWI9ZYlAWgog4aXW
eYh9SpFWNwNwQHBltktW3g2O8fKANhMIYiFy1i2Gif6Ga/XMQmqCPsp6J6Nr6LO+zquTOI/PlShC
sOXPCgXhV1sQNl363R9y4HL1DEGraMUxPPGez7OFpR95QBZXgomIOhNv5RtZdGRRKF6zmsQY8E9C
cUx6hiXQTzLbwzrmykQqzSFn8gic4fizMrYkODB25enSIsSjK5snuHR8Z5WhJRe/czPrWmZyIE3b
dUei3WdSaMkodeHEybMt2qzRDcKEeZWc+Rr8h+VNvZgesUOqlDJW1479Srijet3W07n/rIICrQQX
1vHqTPgVSqKavDPNSSdaYQ98Ci1ZrGXPRXY3ew4MYTqtMMbEfQhlWMvpL26oq/wZUlXOU6o3z967
Wvst9qaqWrgd/MK5mFUF6ZSY7SnzgoslMEzTOtoKLMrOgx3DeEY/Hpj/lPdzXBOwgVf8y9Cnj8Kb
Tij2d1aehLffkAyVRYMemhvzaC+i4ToK4xgFxzfxicuh2DtOFjqyPoE7nuSURm4wYbcl7JiAH08R
vp94KxU0eDgfAaaMZNLMfPDiOG+SeT34uNtlAeX7HlPoo+lE61qU4MMOdoZH3K9YheIO46AY+HcC
5aBdnOgoSW97GVAFG8ckLyqgg144EmcDGRJxNCWSYgoKigWukC97+LnCtgWw8Yrvq7S3cO8E49Xf
WpDMlF0n9Y3LoXKk/9PYV8KnfyCgFsN7pJP5GNqHNUqqFaNsdriCjscONgr1vMRo+HkyhgOjmVXD
AyOfrTcU9c68OcA3TnVUoq/UyzsRMsiJCEq89kxTD/6J5vzFufRDNzX2PwOJIhKSEm1WvmC954vR
fVFogEP8D1eyYTxFso3XN4Vf+Jox7kioAdpu2RRwAif79vBWeQBwjCQO8QD4gqH0XEDidLiEFgkt
RHTbRgTgBlKSxcqSR6chgNxYmwTzS8s4Ks3Ilwc0HF/moPwjmt1DlelsH9cUPwNF8n57qUV3l3PX
V5i76qTim0tiNrHleVCwmvNv8r65djwwtRADQnNLDJjD7Agev0DeR4T1v9y6kctPgrFJVxVD8aIV
iEpTx/XgHUGbUAkiUhXKZkoR7Hq08zJXaBXshuqzK1My18bEEukSpON2+4G9Bo4ngUHKiRlMwjMb
IN6bEkqtYLmKwQWdBW9Mx/bJ6bQNgxpC6z8KgzAxOBPZlObgqMdqhZ/YHAJZE5yMPoUE00GffP9Z
XEmruIawgEcj7NK0+k4mYa4V0+RU8K7Xb88ZVvM9QLZDcns8Zwj93rfeGhl7o8IEnSvP3szhkdAv
wCVXEgcqPc71vqQvtszmO1dEpU2kiWB17mKXcvSSfeg/UJbWWzggm2rtVogVd6kZI61tVZ1yiRMt
48rdlEkpAjxwTKYmzZ/g5C8wtfOS43szLNA56NU7kQx0n4KfuBFxraWS5AbgKDiUUKYp4L0hP+P7
HqLTPE4WF/t4UWXSEZNaYe4Syk259LMWzzyvWJGvknLBwWIViJYQIxAKX/QtUQjI/2uiwKxF/GJr
LiPvqzsWstaKTfzNZNQjsF7lnfjtunZGv1VSVINapHgsaznEguIUivT12cxqCKf0CMK+F0rOupJY
zW4fcHk+IlWasizKGtaRZhdMtPWDZUABXq/xz2s9hNVjHhO5jrVAQ1IQKxQa3KKQHEMw0dWuww8O
XNMRCxZ7TAwDqBXQqH58K4tdUE3HLyDhWiR1ht6ohdKIP8RtRh0AjpgodMvB8htoyqcOlOXBgaCU
rQpV69j78HGiQjieQWk2BRvYW9rhOdfpKYQZLXCQdfprQZHZCW1LMvBL23vbXoVHcUrpf+ZJVjv6
EI5FSJb88399shFggGnDza4dIWmSUVfvuutYWw6P5U1VFJVEAP9ugS9FYFuvxH2gg8n+ovxAc7i2
ru2OEVvvsCPaZQ6iRY2w48LI5tty+qATvryZ4Zk3BEyNy9sJN8xZ3NWe7yrbDyce1S18chNmYZn5
JktZVUwJBZKsx2m5OIl1gz14TdhiEYDfbn4tfngUIoz3sFk8OXXSp1lex5C8S/ru1r7/DzrugmGJ
oq50R7Ls0ATyrydkYxJ9hZvE0/XCMbsNpeLzb/kU1yWvD0+/PcG5u6t1COX9Q8ZqgOjjMr2vLkur
20NlHE2GZn6gVhhySHhiXj24wOzVsMH8FGMcaOOGTxsZBzo/2G/nUWpS0TwGahychSC5lMO72gAl
xGFoi5StLQTvmKTtJuW+HdjLQU6tSKtDRqjnCAyHK2T0UbuBb5jszcXV1h5wzoAF/g6dGWc7qIut
TQu7Yi5BNSH6EO0i9fFkX2egQtrMFGNdqSUcwMkKftBSwkJSgox0rAXvulFLrkVQfxCUkcpDnH0Z
F7YeJE8JKkdDKIRCXmMFyIpudplQRl2aAXbWbiPnE0SbeLCe+wqHRqkw5cqyOr5LnaVn+fz8lNY9
BsMIWQP9Y16bHF8eQoFdWNrrWGJ8jXjfjf5AtSTddCjJfBnunTvOQ5sLFbshwI0WdAzcU+SdChfs
B3zTZpKsL2eDpvQkRYiL9hc+W4UEqz+1Z90B6kXVjgICUOJLJhmiR4OqFfkpX4bFMJRrrS+Zd1MG
QRmwzojezXK4m+qlwkbeCCmhe9wNSjdsmPSHLjoblhXagICXuKd3V8VQoScwpRLqOglfKiuq6z87
4edbjcaWYxs9CoAojbhqZ8QB34tqk9xoMJFjrR4h73QGbwGTN2scjXfL5+ogIqY49161n2/RWeVG
Ge55VfUCN8wYAtMT+xH3SEABxL+NydN/adQVZ1kqAMUUoW7Rcemou7gWiRFDztW6+GEN3s2aN6uB
RuCwZAKEBIg3sfUwWLCZyYFk3/vZa5WBSvcq7Ij5iuDFnFlZCzkMBPyXFbdHr1IlwDjyhSFEA25L
pAujjDIcSynjjwBhjwVY8ThsdjH7T1bQ4OZ5vqCkI39MAMqGtmv9ESvbnCgx+RQynPi1vLwuBbLp
ntFHFXsn7d0Ej1doqB98j+qM852YbRv3giaxGGSTde8o+XzsALHY/PdNwJcfg/OJZmZhbx2q92Z3
/nOA5brWA+evHsHU2q2OlVsuFIA3yBMcyWCX7LV40/8u+5Y/404jfq8OybdPPYbrvivtOu7gFS/I
vCOwc83NylYZIIKOcbjTE8vmd3Y6oOFwXog8knVNCVlhah/Jsgs//rVnrD3mkMrBxKQ7Rvmim0BR
B/XyqPLhilR+ZawkXUmHy9AnDoEag4WEOPn9w/4Cff0J6mJWIorp2FpYey28xCdnxye3aeJys/y/
TGFXyQo2TWvvcFElXPew5F3nnSEek1oiC6oMOlhbuHJp8Z3I+hxVLjlutU2yPxeydkyPGu8Hlyj/
SIWu0Rn/Ew8HOouyukBbOBEmLWSkOSNEzVx9sfsOI93P5HPpu1SApqgEvhXYlfAuO4sX/NYsQytK
clWWMnDukUtoyOR3xyygaAeL622g1Ri/QPFQ87w5aBeo+hhGunvI8B4kXptPSRo07EGeqdma6kea
dJHip0bQc7Vy0bDrUA4OLa2bq1ldcYx2NF9fAjnm42Kj7PGOOpzT41QCMOlEuk46jyiiRJhmOcLk
7Ebw4VpJ9Ky8gPsKqT1XPtsmdewJPb/bDzztgvpXBnxdbknhEa0igVRh7hooj7pcfKfC3JhdEY2a
OitORraG1mkIv+SruHFKqXE8RCLfhQBZRHMsm1IusOV1QWECabn8fr40TxjxLI5qdairn2wujWWM
sI/p055yngXjAmNKCS5iPB1cqfkCy14SeGiCkLAPLpGNrj3hXHFy6hfiLUoYzSW4GF8gz+U1Woyl
Duo1x/PQgLLctQNpriEiBumv5HpNSh+rfmSqMR/cFUnUf2w6Qv3MN3W4m1HcNkNX1gmJw+X7Eh06
Z93O6S38/6oa/HJmPHDCjZFuonXEi2HGBEimQA06TRXL/rVAgJgv0l1W+BC8swIk8Be6G00dlpi8
jxMsc31f74Udi2aXa7DtfDqYEH8vyFH7PVurCtz4tuADP5udBqNvSQtDf0xyuUZu5zElPNKHddLI
qmTqyVpw0qrJ+pc2Iqf/pnsE4xDp0rRhi6qDGo1OHXMfUbLzLrsbWTJUgUjxmBHONMoAj7AjOSNX
O9P3gz0hYBa9NLUh5Wpto4KdJj5bpePUhT/wN1LZ2qDvO30OA6JgUL6n69s4f5l63Yw0tBZxZJnd
1Muy2jCjK4aT23L1q04jbcjAwAw4FQyWN04ysXTwYykXjFfadPGWoQ5Zs71wC5aNBuTQQi8C74la
0Kh3up2/AnV1fgQ6rvjFkMW9pik4o2AwqGrwju8jkBCW8a9qlprbBAfZ8x/zr3YGXdv/PKgHTNAA
zOlInc+8o3F87UjX/aA5T9cStlSr/EqRDVRSdPGflULufwfY35ceem5aHq0qH/4EPXgBsWfoTajw
K96Ab3g7yYABGsRYPEaUw0MUczBJ3bXOxXYzLDGFZX12ZGfvwIh3YckuhfLryO3Ri5D9MQx9exwH
d8CL0tgiG/SQz79MTXVsAdQNGIl9nMysZabRicgRpF37Nr4r7E7modQxX5F8nuebtG1YjfXy/5ja
INy9SCZARFIJ6rp+Yidm4xtgLvMsVKfgr893BiksSqZaEGNFqNygnzqws57E84rWZi7ENgH5ld4V
Ed3XYrR1p5Yq3cAjZJ4G44YyndbKIAaUY6BfXaqF0RokzDByk6+Utr+JLudsKyuIA1w9mlworWuH
VnC8nxgDmGjAbqd7Vu1phVF2QVvCv1t4ucurSG6CfEKNHUSqpxk6UTRRq5fjileu3oFinJLPd4kG
pBpLk2qI8lua2mqyM3O8reSfP02xZL9eZ29vUYaqhrPRclmbWrwTKC/WrOg3ZpZ1IrrLidF+zkg5
uhgutPz6BY2+dJ5Sqpx0saEYZsMxyj7lkDUj6vBdEhj0u2i/ksrIBLT18iWdIjiHKufkCx6PBfsL
r8t0DRa4B5f5oSP2GW2b+frNKgYUq0/M2rRDC3+AiaolJOwXNVcG12Aj2uIZZChMySo+4a+R5Q5K
6WZZQZG9aGSBLYLkdgQW+lmMUL4og+zkia+LpmN28p5I9v4goY3dl35l7iArydIqhwp5FlXRKfE7
j2dSiYSRC8eOfqCIxw8bysg5z+k82Yjgg2I55SD+90mcgFOaLOo/LOSlytztVwe/GuJpCyAdsLoJ
rkXt45hC6NZCpbtGRr0qwEG+Gi0bJOLxmW5llwdZGweoVdrU1inshAXHHqtbaY9B+RZ4yOM2WQwb
keVBLPiPDvlH+0YsWz1Tehys4H8yX1uNO8bqZEYyX+w/KDB5cCSDvJYN40/41o5BD0uidvFz92/n
YPRv36/kDdVsWx6qc1xIlx2n1iubSR3U2I8C9dln6E4k4RTT0lynHSnTgIyn0dpsBgvT4mziAUEY
O4rYQKHmbpOXp97bslYhqKGHbEG21DuUCthPUsSCAjgbeafhvurvgJhCAbtMBSYn7IVbzBXQh+kP
GW25jJuxLsTnYclO1rjdaGKV7tGk0jmjynA3ndQzKyhCuXcP7rUsSQicK9jZThqObJs/WX6aOfgw
89L/TGwWxKLwgJaWi7qRReVMygBjlxV2Ye4wvGy7FfAx3PUZiWJ4iwqsQ2A/9zksYvkxYPWYfkJ2
2evo7V48IJk0Tuxt2l6slUY2pXlywbBbZtW2vji0NGepdcYAtujMKSo9iLq+LgEZ8uxXmhVY7/wA
E6BWlni/2bTPQbfTJ8JAwO5qDxNMQYC+1/uQFJna2rNNfYfB8Pod9BA59D+te/lPFEvrrvr60sAs
bwKAws+zrCo91qFKTsAYIKEhd9BlI4TwK9KPaKkt6G30zpdCKKms9CbADe4TULHyIrQwaNcOIcl+
axFJJUXf/OgcfMwfAp1Xb5NSeeX0Jed8SG8yq6l69rcQ1QjbtHfGNl3t7TXlDXJHVKG3mQQqczbo
tZ+zVgXFLGq+WMNoLr8G7iQPsO/70eDN3kydoXBKkcz40efhFj4RR2SjG79Pp+lnrf8m0cBwVZ+D
AHgLF0GVM1QcAedT7ldCtVsHsPjWvbYmepYaSS/qMc9VmAwzIR21VjqCj5NAyOO5imb0W/vbuP6d
H6fb+yo9oDN8fWOto8lPku1bGA1DC8Mfdd5TVCEv2OtxN/R9dpn+aMViCiX3RrLcYR/mWGuTZsDh
5aoznh+jo84cC9sBWkjh/D+MzPP0hBxoLfpbI26KgTN/4v9lwp5mC6FUNTkbMcS/l+be6+kWR45t
O8nzIDPi/Lsuk5N2MGN512MvVBqd5/cpiBXgw2MNh5MW6dN8GBMwybDWD3oUfB8W6FELwtVgDrp+
gX83/d056vpbUiD6DzthHUaC8t0JoE7TOaANaDFixnPwK7rj8Om/tzU6kbtmrjQAKfXhCEG4CNfG
YJmnNm2LTh/lOKBImTmKxHO+810FHNvpR1AgF0H0wfmzcZehL093OFpQnZ3bwZKGKtnRyZo4odz1
gw2EBbWK9HpcnQItW3lzJ6A1NxQCh5crhiBRczwSOpwgePkuXJd/EnE8M1bF2eOJGu7ZNNLaBRZe
HfZ/CK6/BYnnRXYp09jUqwGxGehjlxIaplRiXatpxTNYmUXlvld0eopvSnv4P5pJOJuO2VuAfQyJ
9/9OjsG4yE8bFpzSoDKQD8Jr0N7qbF1MgYsrv25XuRgPzLfah+SAkRKkr6iojc+J+j7qdzJcffm8
zHx+QCK7XSY0F5w0Ct3Jruyq2yGWbyasGtu6mKL90kNq0+K6vhl4MKNazXTAm/qNkZhyXHqh3Fw4
TvLoajPM6boAOClw5qtgSkrQZ2kyXKoCvsEhW+6oLk7yhtlQNUvPG+1uoL8EpWqSZiwhFFHaIQ3C
3HDj1cILTsjm4VZlQP5WZzJRb1RbUW9EqhdU5SbyyigkboVQfGH3b98L5iOFHCh+FCgt4I8Tvgk9
yGawxhd/pKSeT73vnsX8rZUdGMr8qF8UPHkPD1z+Q/Vln547lFRAmndeFpOCvBRXbBP6dzpJLdKW
DCXQca/oT7N1QMOJUdHwyQbD1vr454WB+cAxWFtVwOwoSdYGJ07kh6D6vpCnZ0m33G+hJSpqkbXX
V8s3N7AWR6WpDiUmzMpNKRpB6FBYW/0KQEdveUPNVm+BqCmCtb+sTfUHVIxZ58fT1IwQ0WlorgUj
scKlwmHGb5tzqyipdnMI/0nHYENs2xWhIAF6/Mf3o5GTIZ52ks0oXeyH3R7cKnY1jjgwHlAyaXoz
/TEmM5ksPKoJw8J5DSfdmOM4ssCoUGTuQAjV8HOMVMBnP+epNa2FHrRGALlpcl7kOHF6xvnn0d4L
Zm391wbYKDBOD1DdtO0wtcUKLLwSXP4ttXknrjPjyPlihJC1Bx4pkiifZkh/OTnDMg1Ynx5+wXAB
n6uGuIjJTGiMPku4x8hp6IrhNqWUx/qu0+vHR8B3KGuFrftKUl4PwDbHqNqQ9b7453CEdon+x0yx
Iz7gjhX/xVcTvIF6NOvrSjWTLMKpbJzq8uj0rzOl5lbV/pGg1WI7xM1djg36iss0TN2CnnNPY4E+
ohZWd/DSENHfDaQLsPtVbh4WoElHvEWRBrdKxtOq0nHK33p3qN+2mEoJ6r71qAESydVTM09rYxx6
9xP3UMtvuP2nl2kqVJSWORDOwoW+zvfaGv+lFfN2A5VXgDyu6sAcUiS5MCQBysCQwsTiANZ5+9ma
+6NOK5B2m60EKHiCW6Esiyihd4FYBwbuc423K2BRE656A172GUCVAafI1ojI+2EzJkc31iepK4kE
PDCX/i6UMyhAqTEZk1B1C2MTgcokfXN6GwukF1iaFR1H8w+J3u5WKe1/wXn7/GkWDXLZHd82/5n1
qvcFTaMusfCBd6EtOBE5gWtOKntVAW9bvGIHeEI3qDw0060K2itRXmTyUeUPxOn1n0+0CE99fi13
qJOpeBzxaW8fDPMilypBAKQChkqip5QA4lAjesoZ3TzHoLuBf0oITsGNs3FQFWIJ0NmPgexeJ/o8
VRjzPQ42/QMszXWFaCYr/NOQOm+4hov492i/Lb5QPZtOCiArtqmoSBTAkjsVq3q1hmfwMoybJv/P
F62iMezPDbxgT7qNhE38Ml21i0R2gwVSk1mu9Xnx0hWITP+xYEsFuysaDmIOzhQZrgA25yaWisZJ
iPAeu3yIzYi3F8Frh8D458DiVIdBsF2P2xs3V6E/7W4zyBwp9oEDux0I5MM7d+IJdM7oFnMR8WbM
3smGlRzDSJnIAoNdKul/J/+9wSwXGBJM0jxoo9h4uHc2Pal8fIZo1fue8sqFSWFnaqlWb46yVTBS
M194CdnRx/FkwewSUbOPrvXLGDpDBgGHjGJ+EGWA9rFLwsIIvpM9hqOpiJ4Oa4Z4Ldew8aYBohMY
WOHAfgTvLprm4JerHSpThjKgHGb2lFEpWiBw+uuyQoqcdq3EoxpUE2sFcm2K+E2SLmiojDpX6ASN
N5Q7e3gLVvo7vKNttJx4d7T2pkU1cjTSpIrUzS5Cup+xuigXyNyoz8tAy37zWxA6aELWwdrAInOM
pzx/3iWoxFeCm6N09JsBBjsFgIYnSromluoedyAh4E4S6/AiGTUO6tN6V2lRcB+HqyhL5a8QPmup
dGEAsy2KVMmhc3Cx86gdGZzXnpi4QDRCn0BFbfCAAp/Y3b6SLD4ZcwcT2tFBZA9909/dAF2XuWGL
KY+ZicP3l+3erdjjVcpxAsSrgz8Z4TtzykQNKcDQQCNfEfByEp4MstSG6nqMIBn/QNwTXEXZsqdl
2gtxVS+n8Crc18+WHC3+/Irk7K0Yc+Xa7P5jvyr7nDUZXFApXSyyYMdGpl9gWt+Gps0W7Gxq5IoO
KenKL0BZ1I28/U80kIQyL70KpQbK4UkIYTX6O3jaMX3RUSeT0X0DVVENiKKuIez36HQTBkKgOvbI
suA5+9Iu7HxjrlLZuNwXJUXIjx96Ih3M+8mA+GXJ3TMXk9VQnayCQJuaziN65BBJpfW071BMKSQc
vQJldASC78/2nWKbuJg2YrYaoJ8rzzl+j5eA1fH5fKxWvirIui5xIRm9nJFzAoczcfmZ6r2zzlNV
1XbQdpSAyrMAYDQPEq72BwQFthJrzH6gmcNYvdUGJ9nGb4shpqZSCzRm9lvVjXnT9Hf3St7yNiq3
1IruRMtk0oDiIU+aL0FYBaqLxbkrDIr/qV8MuU5xwKseyrKk4ZbAQeP5hwsEGB3tY3ZFEPGj6qBx
rWdyb5J/S4CjmsEXKqb25zDzDPfN2rI2/RL2znbQwlEUhhOZjfwpW29DgX/YH54cgKpYx183D0ka
xphjiFCBozjpS2WIJqknZ/8ykxflnOax+d2t2bU21o1jVsnNdzU4y6i0unBnMZarfUg4oB3MZZeV
OV72RkWjC45WDX7twORO5cz7TWIyCiqf2gCsiVp2OwJA8ldmzQQunrfFGKQfhZYy/lqb+PYnZYme
IG7wVa6QvXVH1uzKA7oW3F0KVKg0CCjb0jFysUL+BBwIVNE9lgs4CPvOISxkTPUxJ4Vj5SvA5HGM
pqNBEEG9ogYOJYGZN+yFdip5lLcxOX9sAFzY0RMOg4UTKUPY9uBb/752DZ+7I1RtCb82nytjVbUK
T37wE8z5ND2aY6v3/Ez2YF4XQX8JV+6rAd8ZSXLQVszFOfI6qLKsTVdQmVIyX65WVxy7h3YnMiuI
qd4KEIl+xSBZxzmLeUq7QIeWfwCNdCgm24NmCr974XVvMWfDYw32V+5omcNPqoSrmoWpoP/hvCxh
+rrXQRLwJzHtx6W0OJ7wmrZTiyX3ah5avUJkUtuh2kKp1AtWcCKnUx0l1AoGjUkmd0nK/b6VZNWG
CHa0d7awyXgcC+m3RGrjNlxWE5jeWfL4zSsRBiJ9yPJG2rHQX4SBOF7Fknb5mhRp6ogBCx0KHFgi
La4dA9ttisylnPhR0hnPZ0tHC61Mk9/hTAJDHRm609vn6/aIWj/oGf+uk1QYwFI4LGXDKaJWPILt
clwUHf46EPsUJrV+LFCbkNf5hi+7sa2pUHiCEPEvlDZXn6/TT35N7j578/gDoUarxAVfoVt6td7w
/+lmjNstgorB6Uecu3g+J0ulKcROZ8GD2n3ExD4C55y6oDJclI0SsysEwu2f4YIrLAxF/tKr7kia
yAEEtjbz9DakFRLi8ffHxBTvUiAHAT2YBJ9lyJv5rGm9kZw+yn5yTlNtEWF7gAvGkt3JGSEVM8i5
/2yPY2gbeZkAwm4mBiVEC3LUfJJNwFfmNqs8JPQwzrFg/vI0eWOAVq4YPsjBVzxGnKcBuSGM2mSy
cQBcG7qXAYOE52zTcljlqBuWpfgK3Q/lazZvN4jBH2VVCm7XRGfysrlWs87eaNabByTK1+6Onv6x
02cPwdEtFxu/GVTp6++0GUEP709LXJHnZcFqkrd2JhH1hqhcnMaG5EPR3K3WlMUMfMIQRXRYaVRu
I9xnsC0/l6Rh1FsYTGdD93zGmqqcs3MTY1Ea95fDpqOEQmTY84Y1wgYnLlGa8o+H72YajFQuLQOg
1tzq0gcE5QNkj4JvABY+TC/rnU6WGuPOEzcu/q5G9pcwUiIVfOvrW1b7XCw8m003Z6pE28qiz94O
nzKcd2rTnQTr3wb+3enmNaQutjmFdrgsFe172He/gtRWEpwIUvN3oGZynet04ldF74eg9Jys1pV4
xiUtm61BAFmrVC/OJTng8vtgmnAqi0jG4DVkDDy5xD5O9C/Qv0gCfRUGScCI6MSQ1C6G1PK3I9dd
+9QrWNA/H1xKmL4iAw7KXEZLT0LWzk/kerTB2BmnmAzDiPW/gFr0ne88gAScpN66APrBKiQeOanV
B8j7SniTCv5+GCAQN+nlJMIxtM6LJ3/WAgse8hxlOCl28WFgAd7jyV6a1vKUwGnHHQ9oKOwKqgvA
EnzWj5OffCA7q7wVlMNoV0tuTxE2blbj4CHcBx+vgBghYt4EsU7/JJGXKcrVK+PMfyfluNxcNsTL
BTzQayOtoqSIdF7Dlbtqk6rEgrrNgOvHf9x1fScGLPc56puIrwqutzWyySJDOy6OccYVCWE/wH+8
4lB1JJq/hLfhuOx1yXUzO585aNk41g2uz45Nf4Ue324L7zOBvC9DUblmYTCdqJtfM5dbUZJ/lE+n
slnQoq+q5kF8h2mD7XvEl4G1mK3xyk5tLCFbaI4A2HnNLA/vaEQ3ejUzqV5vA5lBjAtUYmMg9lJq
8ntjTDdlPWAOWwDaQVTzvY+VgagrneXWzS5tJRCSQvj+X1Qu0Ex7rlcBMahcrAaiwY8Z9yBMagBW
OELzn7NjzVh4GOxCo1nEBJPMC/+v8IO5S9RGOCH8lNKkfc8Ratoyq+x3xb316j3xOXI+pzHlCPjT
ntiFzjtPTf4h00C82acIzyys7yYaRIaMLewoodiulNRt2u243qIgdffWM8LcqsqvJMZh4RRRqsfT
T3H+Sia9FVNVYg8cQRldVIJfWf6XSjzdkb+r+uJHh2JJ8GDhgPb+GXkmp6nnr0YeUYTe2MHUEuxs
OA9xtMIK0e2saO5njYKLjBFkY5PZGcsrRte4bi4ELGPgpztcu7aQ9G1ct7M4mSlyrC800Z6ooLb+
x4WZjaV1PcpFcXGOm5W2FqIhXfQRpN4ufL+1C5a5+LNQf3i5Jdojq10mCqhqNlp1vzZlMiK7MEES
UAqxRBjuBVLHs7XH5MwmrftSLmbtNi9uzgtBVRFYl0fEHd/HhLYmXGIg7RBGNjhQkscEZ996fZiU
aAG0mSrcM/5jbjLh7WZIzQPN8i4JJKqOahu6bZ5PQ6y9w1Bwtm+k9a8WueWrpp3Z98b4KhReoUSk
AeqwOw/L5pWD+NSrpakp7Yy1dBw50M0kzWr61SY7uJhU9gn5pRIkqy/5sWRslpGXdetMjYAt6djA
69x+8WrwP7x967XxarPI/Y4zNMfw7CezvFNGzEH3O+6aD8K7+kqHMfsPJzt1o8nNYKshTXmcE5pz
VFA58hKO+zym5O7RYE94k3HnJ/MKQVCiNLqejWSaboodJqwyl0jX+EGhjM8+OcwS4bzPjFxYFr+/
nP/3OtKMB7voIZJceO8YZYY0mc4xUPmVNk1fy60egILCtSlRglXBPr9TMFUgSYf4KBDX+MN4vQDM
oR30A3e5lw4VNMakC1HN2aGNgxGntFl/zxkxljT1aEWB/5xOskESG4WtlmQQl6eKOx/jIOZLKzOo
gUWVva3i5CqCozk1IniM96JmXPGDrQsw7Yswom3jAgoMqkBFxlBXaSm2rYnJlmQy4vz4yzpbxpXi
49W+rNzm1Y4UOEq/2rjZ5hHJTcPjW+Nd/Cw1sEzGbC9zETTthETbYO/ZObBkpcVVMg3cuPiVPuNo
pmjYtw/MbMnrEMw9v0V5F8k7gvpoBYZWzcUrb1GxO+P1Jj3gKNAue6BtA4nYvEl0SU3xhHcVUjgn
qG4RDwYx9xFJ8v0vEjDCUGzzx9AG1VpWDx1I0WrNThlZl2HL7A7gyX9V7qHCtfcn4JP1ncjq7OCz
hkl1wLlv0dIOzIQnESY07npGQHrrfb6bq3PVxCxYov65AhNaTfX5TK2MnEOyfDtal+j3tsbLtlsW
uYzJnpAtjCZHq+c4+Nnkl8PKB/SdxkunJIbgZ053QCHCawAKNP9z81TTWY62vDF2toElKG4ErXBg
3z1rkOv6oZINlRPmyi5nC7O3cumbOPK0lz8JeFMKPXzvjWQCHLB1fom675TE3sF2G6vIquf9iP5i
YBsNB1GjotrITgcKRCrivmBdDnUn2x9sUU2/mFkz9D1QLMudz+u53XNty1+NMoubOCKdW72y+KFG
HxWG4B9jHz5vnDycYjEVkGdBEFXPplIaFNWN1g71eNrb14/xSmPMRLiWFPt2lDYk9sH9B5dKURpp
Ymor/qPV3naDQhk07ZyfAQhCNfAhy/4vN3JqCzlbTZb8nUc6mpl9NHfCknjMmAhvTEtxlfIIq7DW
L1HnMnsFTIwGyB4sszJePoZlY7bEbvjUHm5ohuc6OQePcXj/NcZOBmABWLVIqEuKe2dcMZnDnEFb
qc+fTxGU+eq7L7HsI0urNgeZ3ffSsPgRCAQajEtTqh7CaRcwuhwiMnyPzhqsJ3q+PjWZsc22Mms6
tifpBR6Vks7JwNHD6GaFn3932Oj873gNySba2Cug0hSC68LTKNQQHqhv7SYZqXtctnmCymbbPkFH
DY8m6vypGNDT9DOqeTMMHqErF9hmmrUN0wYyIKoZ97yT77J20wpXiMGV6WPibx6egT+Z8kxMWpqC
bBFI+8l+5otyR3ZMGpg+1z1cvXK4gsWXcJsG99GLD5cWd5fGjm3TrmTIBXdqx22pSBHZkvwJeqV/
toWsMifWGa2i/gZrWez5vcv9jvKlhx9iXCi3xfatq8bRbOJf09y0JNy9W/x0MX/kesd/0OXyfD2n
bc8A8ypcGuS1ZACdPW+WulGJc+R7t5LE+MlkSKrNbUaGlBUGI8VMLhFH1xS7DtqiuMERpR+DjzuU
mEX5rZlr97FuqjR9p894yamp5ZZYLVkH64M3rEgQ/VLcMdqxUwzLXStM6GzsMUk7nfHcA0goam0X
Fr2umLWaIpuRZOElrVKC8Tr6gKrS4z7S9n6b0+Zxf0B0wyJbpAFXdlew4U4ENyi26UcDttlbz/g2
ikjp+/FrW7DMvFtU/tqJzSQt9BCBnIfgWzYF6nO9vozmvM5c1wEv+UAZt0dNNIv38qV8Jdoj9e3A
Z6ftUKnYsiEZcJCCFTlRrd6AU2EMQp3cnfnAFat/E/Qa1RrhYG9lccptHSKfnD7rkj85m8KvHta0
kfc/MIVxhAlu5u/0ATQAVNbNnBEkb7P8OiGFLpoRz1sjLtUmkNzZtXUA05+iSr1zh7NvsrimmGtQ
liARH1FGnsmXpWUgKHVWVFetF65F1ROdY7RqXzJ/SHDRTftA3DePiNsB/vU4S+F4JBLy/0rETh25
WsBGxMCqzbO9j5VwZT7M/YERlWqJgexlcR8NLLVFNr6C3ch5l5S82q8u0h1oo2+3NAYVd8xl/yn5
1TwHgW+EOFfevSiZgJSReYK7m+EqY1W8NWHCQ+Lw4/1g0GQdBmdsjBBV/5Rq+KI7qr7dSRwVP2Bw
WDFBEKpEvQj32/uH6XlDSDoA8zZtKCdmIxw0H5ZtQgKd8e6MQaByMN22YwhaJv9Jntq0ZmMpCNhh
KNcSq0EDI76p7yCkWwH0dsoMNMqacfiagqyPvBCn7cNL7APH0ziLY9GXxUQ5z4ZrK/GbhKm8HVKT
8Km/u892uU0TZnBNbsBlDAvs4E/Mo3L83CsodP8H/hAGGAfpvG/Sj/ykI6Pc13M1/I6BQOmo8G59
fdSVMGu8EfMV6l5KI++z5Hju+t++BpdKkEENETbNK2TQlmMtD2ojWxTttpI2fXLoVrjji2vR41Lp
tl7kghHE/37mFdybSxZAzvSyB4YbxPeimoYqpSqNwixK/kF/DyTe5LxJjewiiOFejiS70nkG8XJK
pymuRVqHinJ9TQc3x5frKaLlmQXodWBo/fZg+p3gbSFX4yi8rAd+IRIXu3aKJSgPsMvp67L2bd4S
hZKzboxQoWrfkqLi0bYZxKvSwuM1Ffw/L5z0VGb1XdzlfkU9tcj1C4KVzT6j+A5JYcXKtAQ56rOK
h7R0tbpUYvu1YLlRToXdkmunMaQf1kH5wxtXrFQAfH+ZfFdlnPWZC4JuAC3jzO6TClyoHjsjG7td
93emhlQnCw7d0YwbPssUUHCWshiVTBGOL4brBGR5Mdl5JbqVXwkAiWN9qMcXNMzh8Z4rBUQyfcml
0dw9jPLyQtDrd225P76lR/2eCEVQ+ecQm6a8l8O7rwP45PwPh4yldSwimiNvoEjpkwYETQTn5Vqt
JsPjyI2gdYSrLoaWDQkXWilHb6CU+sVPoXL/328hy2XPZeQl7qjMZIGnwWgHle3SGl8kVxAJsNwB
AQcmeW281d2ptKbPJpn2uBJslRl9GyQPgf1iWT4ZVHNBGcxXVwrGJXj7BEZ/2/9a695TQGJQ6K+I
Ts9H+sIycYIVXC4qCqC/x3R1fDq29BLOxyy90hDPsPivgcmIcDceFjAd1/Qdui0pHPdnRxzBw/K+
2AFkggAQgl0rPEMVtftOPoAIM7nU9/LXwsH9/i8c+vykfVFeOF5bPbr4UExyU0DoH0hUORKhXcjO
UiJYSxynpGqMqgUyEV9QLVMjY3Lwque8fzblyN3sLzk0+uRyNZmcGESiA+sdyFrrrz8GTdFafI/c
HX+NCM7UDlT98jYKzSPdYbxgRlf57x2aW16hJTCNe3+MY6xj2xIBnedI8YTER07qFL0o+Y8+2atO
PXWZNr7rUpv/bhDOjNmA8Yn0N08x2BLjIc9v8FiYb/q+GpQ2qaA9qxFr36bTmFMaZcRW+fxzmyoM
IHbPCFSiEBkEQthoIxaxx6bA7eOXkUXB/qsAo6TQemaYU+vAlioOImgREl+5I5+Y5I6EHF/LJT6z
U8HjZHcnxd4OxflD3XSJiMW3Doy56LydD54I5pdOPH+U7vMSyLinq0SCrCySmypvhIr6bXtK1rpF
MmOOthqM5IHsFtUpke8I6Oic/3Xugo9H+zAmaEf0xUvsK7j0DQd02caZpYs08PPyKkKwgP76MZF/
BTKKyuLl7RctKvxBbER1T9QBe0oB2KaIKZNotMhdbb98Ov+vhPrjVqQLYtyu7NqWhpZgTCxuym5i
hMmrrTTO1rzwvgUjUanY1BDRGQDeQH7NUz2zSDKR9Nr4vLsJSj9dnihy5cmwhKk5M8TipBHlynLh
pfcuA/DsKkGtyE106Tdj+vHK56y7pOOFwgEB11XcijNM54IQDi6P71paH05QDmmfMs8mUgbC/i5v
8GMt95myCdpUjdQ6+L3r0j4RgaXmeBiXvVNFpWdoDNu8WGv5lh8fTZ6mUYhMRlciYjy4Ndrh33ru
KGQl1ZuNiDEogQg3JDtEhcADydP7xTopEKBDjaFirzNjAQJBXKBvW/H/hLL5sIaNWItpAuacgbA/
o7ZLQDKOIwTGFBFEg9pESM99FLH0twbT1OpAYD3/MrNoWCSnkhm/ZTGgm3Cx43tFYxVSJgglzekc
fvWvNdqF3zQVCOUh3xhd6RtDqFi8EjWu+E3mCAozwZkdSr8/XGLEhMDN20OYsixmVHloA9Ojr+Zl
j3P8dgOFqp2lAgiDe8uLSjELMMqAc3MwAC/PEmwVFGK7rmGtXYVlvhxF4sHncY7LpeOfoFYDAITT
3euqmJYjEaAAnB2qMgWYgAVmn6hFRLMhM7cmVmrXUqOZDcwSwGM6OJrML34+yfRav402/gpl/i2r
XfO7bTsghOMPcFE4reIm2v6shKTX8zWc0nRBazzxxvOB8lauz2gU7aHFg94ApHO9VowbEd0PPiLR
oZ+Va9QqgwVjq0RC8mLwdX0O4ZzaHVeQcxqZ6B+VM5ZTpZO8tJXgZCA6SSYuUZPttbfKCPhBwZdb
WN/cMqjjtWUaMLJdTo1bL6zyzMojIfPpisCR+F/y8pHbrFNy5XvNOsEakSYV4m8mX/LLguBErZ+u
LSmbFBD+br7BLL3ogUHIbL+ui+kSbd8UzUq6OHbmJ73uN98eYtHA4wjIrWNs6NIG0mBqgu4Xaugh
LQHlBImXwnesEQOxxV7y4ezHAhrj/9+qE4QuUQ3Wjjo1ktnshUlEUge7CBJ69x0sTmsrm4Pl5g+b
t8xSENvDovIIyqlV1O3XqeTmR4b6wzIyFKsRWhiK14X5TwKWtR/M5HVrOcHv3F3SmTbSzjnUfUqX
p7e9xTFsEr5vuXw0h9i0gDPMHwt8YfoYTvlnOMI1SwuqLCu3xi5TPN/mdCSCYHRtLWts9yUetpby
7E6/bF7V+MsUn9A+tp0RdxS6XUTgX/zSCED5ctN5f4bO/eTHDI59dI6NG8XeME0dUhcDj5+v/MB1
OVh/Ns9dbsm0hCzK0Qz5wRK/+tJRIEcZhmXw/2HMgYdZmmA+pS08sUkCiHZSd2JEpjS7xWaNPhfE
H0wKf5QifcwxjZrgkskVDiyrgIL1u3Hg2Ghi+dfy/w4o//815DK+oDRln8IFwz6iWDh8EWgyYkYL
SVVDjZ/2hlGxb6ftmPq3lqINDA8wkByg0Em/yr4uXsG78wmKEgWzwTJXX0XDQwRT9X+O4azkay6U
S8DL+TZ9jAhR727Z+n4wU3kcsKyCUc1pHxUx6YW6JnuOVLDAR9GwynrHTIJz/6sIMXC0RngpmGNW
gmhEB4gECFbQc++oObpSxAc6B9qEcAw3KenSll5qeVn1jyt5lIcqLNJh+ZlcuVdj41Bg2CUJmigw
KX+zPfXzP5rN0F8LWY2qb3nYpXmxb4jJ3k9ZnxWWXuFu1c8c35elh3PRui44MvFwWqg7mwrn01C4
FxdSUEY+WQCEKtgHKsjGd6yqXfurBV9M7w2o/A2XZc3HnE2HXj6/CY4UXV5ASnVTw+0j8MhhNhtp
d4O3zn7yuvOP2Eb1queifJiOw6tsLeK1zmE3Xl25h/ZUHI+CsLxchg4ud/M59fMRo1L54JBrKBk9
Q2BECF5Onyup6X4xrgZZYvRQ1/QhtAyWuyMrF7C3ADoQZYiOhKzPxcoPhrBH8KMkWW2nmn+owgAf
OkkeDGjRniJiJ+9HYtst4tG4qvIWyJ4ZkkBZreJNAiSvvajym5Kmrdi5mVn2RRX1DRBpjae2vYh2
JGBpPfRBz0/+U47lk/mjrm7s1Cpfd05TYyztYgiHXokXAvyuUYEEZeUGmtDQlzHAfUTXAv3DaKpx
qGLeVgSLxp1RsI/Vw13bBcOgMFd0Q3YIu0BRUXdSYtIZgaQ7WveVAwCJprB0PRu+N2ugPkkeiIbc
Ac26MHFIXak2dKiISblO62RAO4S6SQu5j2IZrnre0EebaN+0wj3Conpe7NGvBurjy8Cm8o/ncebN
cPOH5Y9F/9+edETxf/5BZZaICy/1dOsX2YsSqZedpAjTKbyj6YslLfxHVWzQWIGhcfJy6/crP+MZ
zY0/g7gfNXbSKGe14EFNjQsADgpx5Gh7fRBYGkJ2kb76TiqD/W+1Py5MWJmX+6ELjy/iZNYLvujm
RVGQbrmYoAs8IpdfK3oqigQ6r32cEBA2DfgGwQRm3/JsXWMuucTqVfrZwgVRBBWyOpSwkhw5zWPG
t2DRL9xWMpygU6ZLgD9YcKP2IJLsJKdVWP9VC4E44dOEC94tkXDnVnieT2DePJMz0ISsEAt3EUF+
S9+H8fMMPAjbY+FqadJJugfK47zE5M75hkSxa0Pxlw+WceMZQW8s0iSFpjuFM19mjmkK+rzP+fWt
XTv3anDIiH1XTnPNe+gSXcR7q1SdbXG1zJW8wKNB0lFyoYwviLC5ZAYjcyn6E8yBz79Zljb7lHRM
/j0DDbo3t8NInY0sw/+rGGuqz+/AaY1DTnj6mgxUi8SDajZjxh5HhovjehRBm6Jx5MIjHhhgCAlD
VRbAFq/XSCgb8yj1JNBTAnN7RiJLHb0lFzFtR7rtTKQ+EJq1D5U/agZBynTNITY4/1Dho6hziLtC
kq92EH3iUS+Rd9/qWoaugn+nr5fBOX+zfVGjhclaOuiDp8ZDpys2dCs+qwIEVwLLjjzjU4JgOPBJ
AuEc9hnuxy5KwAtEGAGrdXqoIiaKEXY3T/cM8oe58tZS7nvLalKY+Ee+D7jg0xrmugvyWW/YDa9G
FBLG/9a0hJnWUD3cX31USsSCFc+HnoRUKslejMCEPyTa8AeAVoOhaunaASc4PvIMQcgVNt5CnKBd
qUpzw+MlBIpQcvObzR8er1vCpdJP1PxOZpXE6+OOg/q6SsCotkz25iOsNeEpfOXZ5F9Gn6LfNpCN
WNFv9OOJNUj4SQCeo0j94tfSVSt/ewcaAoSvYkuBC7csANrHkgZPL6kwnoWO+vbwpJL2Rg/wgH3g
ckQO1QhlI6tyNxXz1GVzjzo2NilftZVgMuf4iaR4JOp4CESg5dJo6U6/H740xv/yNPRxdC3lgC9X
01H8tdOgs60ukEe+TcMJMWQ4hXKUQpDWWrPS8Z2FB1W0Vq5lQLVVWCXd/2BUfWV5wfwI/SzExVk6
S41e+wFG5eE08GpaL5LtVtSqbc494WM4aaUzdwW8XyBcfLdvcM92m2qALPt4NhWpLr8Dxx2tMN4d
bSKzZESkoaofR2xmjd5l8CTt+K1jti2PqUf4A39znrpZ+erXnt8ByIwHdbVifYgWnHLX6Z0nKIAm
SHSeVfLu+aNtPYyOIMSyYq/JKiQsrJpZMdSVwWYQmiIhU4uO2zLtcysmyEuOnw4zPhn7Wf484GiF
1t4Vhe2L6mvQWpihFN9KOfbcH0/k3mo5Pa1Hrqux6QNwwDc8Dhk83uZxhGXcMav47gKud3aOxR6P
iseyvOOqO/AH6mrKfeXR5T2eZZynk6uXP9aMKu4SA5+NDBqhZTyr8sHUUuP5jt0N64pZ0cPyuo09
g7fIKV4m34pVYjRKTdvwxJUBu5l/sMwBUwrG/9qO0aeSDv99sIvVx3w8F8jANZECpdl9rUiSuFqE
C/izjnbwJy51zkEztllhGbNhUpo+tYM/RiNwpXyRIyZqamZVkRVQACrggI3F76vOee/+FC/ptnr+
QNBIpr32OG1Yd2Bz7KLmGW2+h3hvvpvAa3eCmlshfxdHcNSIX8EdpvgrOghWfD5luqzrkvs9QADE
JD9k5l8hr5GP8x7p1dxHdpNbW2mScbQ2nklWZo6hwSqcUUp7mbVTmftFpU2+b8lQ8Vvg1j75x+rC
ANkscFWzMVLYr3ICyIpH/2VBGSz1prWMLuL9btoochZwX2k+g33jskYEJx5E4qOTYEtI/CNXniju
I38+NnH1mkbFqh2zAwfMS5JXIADRk/fXXNkj4MRxMM+nEKzTDTpy5hXTTCgBa18cbt7avmpmB2Pa
Jdiu45xQzKIh2ct88Sf786CCLof0QRXGQQcvcXddjcQIMop0IvurSF8Jc+3JRI8AhtYTSP+Tv18q
XvoEJnbEIejZu2ga1q6ndWBnvoDvlRjroF1xxD4CpH2RqKZZ5AYFo8Axn/gmoLbRDH9hjBJXht7N
aBY0S3TWJ+1XODBVkjTAeQYtm4KqOFdN4cMi6RKGLXp4glJwoCGxIMXL/0VGptw80206wpnz6sJZ
45F1WAUuHjDU05y6iRXcS4R414WAGwIEk+YUXdkj/Kf42Qe+UdH4e38FXuB3wwy1HCHQb13reC3D
aWVp+THI4QLr0NcanWYHxK12Rjizw7TtaM8Rbaj7vaor8uxhgYrdAE23UUQgcJym/mm5Zmd3dQ+J
WdsfAj1z7wdunhTnX7+2klzsZgzMjI1klwRKCek2OwpPtnrb2YwNlktRRbGcvOm7JHm6EheUb2LN
cvxxmhtqjYty7Gi9ew37AOGITQmFQttzt4HScloPcbPeMUPM1GLHhO/UiNl8t1jNdSkcPWwVernS
dNLl5x5XIirTgXqOwsqvw+BS6oUUIj0if0LEtww+L99OIkMcDmDG6qxYvQGBfmlHr7YHGAU1GZVz
8bnSy1ynw8lGs2K+Q410G1e2/UnyT+lrcEW1QDdJIKRyKIqPdYrv2COjJJf8sRibfVNHXCvuk+nX
fKjHSRvvulY2m5ZjbEIJFi3Vrs2CdgKMWkROWZGL0CS0s21XiZRenZUvPBq80yhLs1Zb5BbkA7ff
TEu+W0cPnWQSh1TDRIEwOCmAE29b9udTg3E53KXOOg+885WWuURL6V9jQxEimLub+Z5Gv96jXuGh
NdHh3h32YAtcRaVo1mxaKvDYQaeqF1oZVqgNucr8DldQQSjIJWgrskakUVsxm8izFX06+U9F/Xop
IhFIT+jmqfDx1w5nyEOiuSzKM5czX/6cGva2ofhSBd6s6rjoWQ2jjPy+F+DwS8QzKxzcX/uLz+/m
Y/QwRftGPChG7rqUr7QWYIBxxKfuQ4k3fp6FdY1r0EwE6QAukLSulGeh0+cpJ2hZLkKyWtDmGXEP
0Ach5OJUw66zAD56eQlYnZiDn21PMZi8qnEwcZ9IpV+f9c6bXqguERO6NoSVCxKrOzQiTOfyvX9W
4M2p+SuOnzjySb6K0YsEasg7EqQyCZtbVv4pMkDz7/WNwWCrAwzNZTPIxJI4CkuWUi5ayIlYwX8K
pyKwMYhP5Bz+VV07HwABP7ao4fMsrmZwN1jLzYmH0J7HWZERa0TiV5XnnAXVBzD0UHG3+3+Xa1+1
b3rGdR/95+0Cdv69pUkBt0R4JyJwEqyxhYUril5SWod+luaCW/NUM7PDPoyzUv37Yx8I/X9kyyc5
a4DqgM4JPCSznQPxiVVeHwore4yuyWM/3PQYkO+TJV4iv/0aF10L8yjXHr4jkxHdTVqFkc4WGoCY
4ZYz4riguEQQeqegHOlal/MeCj1yWNm502ERPoxpWUKLvBczeSQdn3RH07ChP3uguN35n3At74ca
BSiPYCOpcqpawEwn+OOZWb/Vp4PgBnjQzRArrrR6LzXLSdk48KS7evmDiez0cYP50NFACdktVjEP
aCgWSrXNVs2SUnjBmYBIowOyCNxMO87ywCD30stfYTTPmZqsd0lMRvKr2OIP8JCQcsbgilyfsvg5
DeTRCJEr96FUkGIiXvIGBNBwbYV25V65eTmhXSAZWZSr6oI0uNuH4c7UYMFeFfKyyjaNnK+bS/qS
GtegIYXKWyMLCf4lBHGMyLJRDMA5ajXQxmdsWjXm+dEXwPqGqhx39ryn6hzFikU+d33U94KnDbgg
uTNPtgXSsFNQb4UNva3tMxF+RTEkwWe6chpHAUT10wAa54rDd9uZFZL7/qFG5qyMdY9KpY2U584M
DaCTELXyXG3JbYctPH1RMdlBFfa2jEicylq8lOd/T277TjO5KedoiI9P5OczSW5EUBhQn+2C7c6Q
gOHAw8woDifBH5eveIrLHiUWVMXxheaRkN1gyQXhsqtXmSXQ6xKNVKVMbO2AxqBeFsZ6sR8cE9Up
5TaC1llA/DtphvoZinRVaxBV0sjf8z0iWBGBQPBPb9XfQTEr7GoA8UulA4JcwNyRQBoCiWLmnJG/
n98CrL/3aEq6gE92BWGBqMDnvThD8fJo6FtrI4hX90VYM1Bpe5Spz3PDox9RxL2D2k+zqB0BbEpP
nq4De0scPjXlKTLQfXM3WGN5+8J+8gGigPBjYULIY3F+h5vVQxbFKHR8uNbYYo7rmnBP+g1SookP
91bCOtB2qTsUCcXpO6tkI9gfRnHB4KPIxBJ+Lx1U0PL31NZhQSk/YoIpW/qcugTlyj0w5DeV2vVh
2gijSMuk9xEI2AnpDQU/YeEyXDPedCL3PnGmNbm+r6kLvkPH3akEPTGMEvBahCiPtMa7NaPjdiKR
MAmSawVI40Drb6GYf1/vXneAz9l1iqrSsNwm9Am9qNi/dIoWWwapHLOl05mK94P/MF0dpJ0wb0Cp
yWVw4Y6dcWNr5VZuoiQxzkGTc7E/umURBMmpu7vKRnTI11t1oWkqakys7vAPCnJ3tK6OcI/Z68Ow
d5O8cq0YKN4YkNorGTCdbUOBNrTo0FUyzHRPglZY/giPHgzoMcghopkpFToKyAm8ukujlZm5er95
o4KDb8knLVeHIx5J0I5Zothu3IkwUcQ5cK+wjmcAcoJkBC6DmuqpMFpHFiiaGj5DUPBkJID8bL5b
ZJztFjH0ztltJrArZ0OvrBeu7ih29VdfgpfH/08sYZObNOwCvHBvBcE6bUzc6VErRJF0zxmZ0y/Z
oFIvK1X00zFXOrZIDXgeRNmxRaq+K/08VeDJxHF3xEzQahlX82Y91pVKC21wbuYLEQtubTlBZVKp
gGUH4ytJQIobltP3qClynRqO99yR/R0ISAeLKJcBlbLEae8qOdiHTNkXtAHfW/rVX4slgqBPQc2/
T5GB4ynXhvq5Qii9YjcJvQjeXgkbYLASMdwMa+owOU+wsJ1qzTk3MZ2tk2QpPutEmqr9ZNtQqvt7
12wQIYa8QhzM4BxKEYBEJgcY6wnhHqo39X0MbuJTvcezR5D91LYO2ewtPfajXTRtAsSwDj8N/X4t
7zyoVODQdci9ckIlQA7ROXpbjaAupIUUUiioCvgUYXSXz4wlpXPhmYgxC5YVP/TfS8fyq/EQslXz
9lyoOP/WxuN2oGTw0Mwzakw9cT4LvR086BK2bnoYoUlqh94zUXLLgHiFkQ3F6+blMP+GMNYogct+
R5pGZJgBOCHHecZ7SKPPOI05+ndBE0VzXEJLIboRzzp8TWj5PgwkTD5YK4BMyEnklvx8i7hQJfuL
2CPa0ZnbliRnZy0RiQXzPxvoMhCV6aV0lD4syiTNtRGw3YEb5Qur6ZpBSxS6LmdCO3mLtzQQOnos
0LjyYTDIcEb3fOaPTk8w6b5hWsTWojgS2HFGIupLl+c85gtAxUMy0sVpK4slJypgbvl0FJ1BWJzg
p01zYtwACVECDa+H9JYoGXmyyUSlehwUmIyWyRePNKX+xm8h0pqCdCeFwohhiJJMcT5mpJq15J3t
3dRakbu+vcZJ68HPKSuzDKuP8AbCBRUBWIKB5zds7vD2PtNyk6C6dxSLuLcbtp8yCt+jGNrMbjV5
MUxMCu7Rg2DUDMhbTwhR7WXTrswMRkwoPI3bGfcrRAr0uL+eDDjtyiTqkYO68ivq7UMXw8GdznUS
06CwJNG0yg0zUOTlBA1UvXK9aHCMytCQoSgPDK8tAZ3IzKcKlISASgg8AIqj+ENxTZvsbPzjgjUM
IXWLyyLsZQ+jsM+rGhHbGk7CVZUzZXZbGobXtisT3znAoZQMsJGEWcVD9E88biiefKMjQyEuV3IJ
x+Icz6G+iskDvSirO7K2QsKRBTHXxsMy/emXhxrw30V+7l174AxL3TFPhyFAlIOKGO53/M/fvWHy
q1Hup1H6pysmrOxgXCx0IPapuCn6QAyHk7Wqhh+ut8rxgUeoXtnKbFBN74tHZksxx2nSmdGVXIvB
Zydnc1/HxxXF69el7BiInGXm6FzfwV1B/R5fx7SLjGHlg1Sx27cnIQHRiIec+D+0ltK530bYv2ML
zZuj+++KtUVnP6G1d9cXLhfCgcdgAGlsAimcC6sqOEAvtHTllbCH8wtns6SNzKPrYPfQjrNbgI6J
ssQLC4UsMqmCTC3Ji7s9OpHKxBfvfRSC4wbRUOLq1772dx7iW+s83EVwLdNo4M2rft2bK3c7Lhmk
tAVFV89rsyuRS50tImBvIZPRIftzwb0B4RY/VWPYryCs6iHx6Pv3wlRZfBQoCY7iE2/cE7e6K/K+
/u01X6X8fNIXJxcCmnGqEK9NDMwyv3ObGHRklneHvR4PTr3oi04aLu3l/wXNBj3Hz1Qfe2wOrl+y
h6I4OCu4aJX70m68FhKOEBeoKVK/biE4zgk38CA/8kjc09u0+9xK8RZ5Av1Z7JwhdkO5cO/6F4aG
nqiNGka1ZbPayHGZbX4H2YC5DL5ZgMCZMdjnReaFXF41fciuijEgwKsvQZgVkZf48ccOkrHaFOqN
bAht1CAbsRKvBXAI0LwWi6xB9ZCEZxW7fJjHPDsllPtUZ91ERjCXUclk2QxwfuHd27yW8OqHjOaZ
TbJvSrnKtdMB5PQjr7cdclOOS1LyPLPSiwJot7GYMVxAidQCFRETQvONqWIBMayBi2st5x01v6kH
2ESZWTV+Lj17okQxhVC0b2rda8sgmkuJMxm62B/Vme+Plj9dweM12F7qlTMFl9IRlT86dUglgaV3
PN2cQDZ8yXT1I/N3dZ+MHZDZ+hNoShSsvihxDrETevl36QPqsZoxnHT/Y3dxW2cWUn5RBq5NQxqR
yODnpVSTwJ00V1aK2HZmN+GgFVUrNOpjztNRQCMGbbv6RBJfbXlqdMVTqZyEsOkv1SmaK+WfWqrC
EmheRh7TiDJhL4W2qBCKsyXHbH3yE8OOVJJsAy7Ljmp1sLSlAtQN/YABdg2FXEIr/UWnNMkOWzKE
39QkH8y767Gv+VQDoaD2NFafhvnoK4kGJfPrSBKB1XS8ipEUCwIDx5bnBPa+a8QPpspWHgI1faBZ
Ix8Uf6vDHWCbu6SAol8gPCZ1ebAx2ak1P7XzQ9m+l86RLT6BZ08OBPqPlDk4izzCKlE9tLzUdT3X
RXP52x73r2MKc04A7bII2zBUPs/dCA0xE6hDkA5qylVccYitfVyiAm38XUcFRJ4vsL4MXwFh5ayu
EtwfeCE4q1tJbTwv1NuS9h9CYSH1xtrPyWCjvItiUJ/zELpDZABvLrz23fcaf/6wiKF0JDbYVEU1
2L9hyrsysVVwMvh1CSasVwxusFr7GhGtitq3K5unjl6n+DW4Ck/EVqRVa7Z4sszvw/d1LUNNRYoe
lud0pfIXhMqW7ARFffM/EZ8xfpkJir8vrKuIFexlYL4x8jBDHQAokZSp4IjumoALUlTMb7N8H8LT
pqnhprk5ac1ROtB5QwRTCh/G+X5G+/cMjFWk7FxBm0tcW1oxg8ZG3rqNcQlUeI22pTRSaz8cg4Zx
BH4ylYe9bHKmCFJpl7yP9sg1SpPNV/wTEfoJv74Kur/cUAF6gESpyQ902tCKKdPpzf48WBrCW9W6
dKAILTYPd4d3pol0qWdSPtQzMP8ss69Wvml6kkrJNPhsXQsE8sJG0HdJwNOQs0QIi8+K1/RXWGAD
kTnOT9Uz6x1G3OmHhGSuG1upuoHeDUdKWN3QbeK1J6yLl9yv7PkoaUp8C1PPYGOmYwtJddvhZOpU
rl1tVg5jDQYvSm6lZr7zs5jn3J2bpJqwnd1AD1ytBX3NvsidDE+2OfQcGAucb+CrgEuVvfG4SbXB
bnPmuO1FsKXeJMd/cl8e9+7GUkm9Pflt0/8YKPsgp6QN1WlyP2jD9jFvhSya3gbuiWm7jqXtqxyg
x3T0zytaVgTBw4jZLKBakrOz5x/ir1fsdjE1Av/uO7Fdjp/T+iZ2c6cXVFYzqVD9f42u96tv+sit
J0h9Lgqz+wOm6RvXHWoeSxAp1Hf6TtVgOG/Ec3Lsii5jzZwMW439TUvvDMu3whEGr8Q1VejffLl5
eEoT4b1JdOQDf3ZS7slZiO6iWNt4v4zhmPDVfShDC7CU1FKQEpmM2PWfXSjeqK6e/bYGjjFsik8s
MjoGpkaMtiHQEE4ou2U3IDcBlzwPe2i169a5uPs8wIetfFzm6z2FNwnNGIKbos4ZSrjNt72sSPpk
wztPJYgkr9vuH7fbguk8JXZhg0/QZyzCuPJ777hAozCfLPZRN9KnauJc0XgmQQsKVYwCv0ZBuBFY
eJbr6g2vI3I30R6yPOYz3IvT9CveViyb6Q5Ng+mUPkf5B+q5FM9cl+2XKJJFLF/b5pd1U4rCr84V
j+3Q5C9dthD5zUzGQnJ75uQbnU2edSJqEh45IKG5u1YCCGpUtYN8xlCURRMsbboWkK2WGCVniPo5
wyiHq6nl6rM4d+Zty5uJF3wB2e5hybLYT5T3YPn6ugDEJLVuXjhFJsMk1++lYwI6lRk1WNK7ZrDj
V6xDz34dFMtdE+ZHwvrK4PI9/LvIHcoLKCPaCLwqSZBiKl55j4Vepz1OIS4aYYJdnQpEW4pUnUqX
cXsHjTWZXI0xx38kz/RYRlun38tX63PNaGclQrAJ1mXAvYDJYOUB5tuJ4P/0OAZIqNi5+gzKK90F
eksGpjUoqV/Si8X+vk7FOjvSNKIdPiPHjJ6golAh+KtciS8nhb0VNZDuMlsciWe2MsaUjZLE0dhp
KhNTGyvEf3VlhXtD1pKr9in2lMTL2qqxH8fHaWYLt14FKTKttdDqKRhLZ4fa6rpt6+i+W35pKkOb
tgwwyp1d2WsLx12PwRUA04Z8YTAXxMkye2MwJZ4dLJOp8LADFU+7BrAj+QbGm/BXLfRPRL+4w1r6
ASO+lK/LApmog/Nd3MPCxHmgrkQxCYPmTNYLjaWaPjFil9+oXj29g+uU0yQD5u67wv1htEN2OetV
BV9JUzIDk9R7k1Kg6eDlHS755lAQx2HDFD79DfgAhuhHPWt7ysXIoOEfPgFo17Dejf/Y1jLBCP5d
XuqsTBtjN8LgmNcigsnryzL6TbI7ZukFw+yFPLyS0P14gKI30VeshVY5I7wWAHM74aKWrAn4M29O
48A4vx+EjduuWd4jQgoEYAp4xvEy8mDhwOHM1ra0089SAJWjRO8c1JL4OAAeZqrfgUEHTIwa73eh
w6EobBp/MMXY1rul8kQmerxkh8knsu/cvX4Dca6pjJJfDPmhPx5QBZQ5K8/cu2n8sm7BoLG8SRG7
wHGJR9k7WqXS0Jy9jLO8twTMEPty6G/RYxVGlMieTbBjriL/4KMvzBF0VyciPm0JRw/kxs60lLgY
Hg+dxMmP5Hp+vgk8iI3WWyCK38EtE8dElJuHGG5DqthkJmPgA83hG3U0jlSMQNef1hA4uxjMoi3i
7WEvAOR1HBPdE/T7nyl/+I306IobsNdP4H16FFL4HWLREHEl1GAyAU2rFrbQ2CBwqh2S2HsosFoI
AZ5vIPSj0181xIe9yqqotHVwFLcPBpJrkQ55TwLOnomdhMChuPdcmDxKAlT0Mo3/jBcY91B0BZqL
huL3AWEnjqKUVfOgDaqcdnFCF5CSYHLYZPjjDGdezhxouT0O95iJQNheTwhBcodvjb/3QmuyiDr9
yyosRqtdthx27gMGbVDUOqnSybuKdqvCI+yU4+tC8oYMc5L84JWWEyfcTVTs4gbtCUkZjBLdj0iU
9I0GcdvJTAZ3i+mzstFJxZ9EHjkywVq4MLPuTBvf+EN5sNXZHPfKhhZnhe6KNFV3mhf4gshryJBk
qrzm5rO503Cjskj2w03oEiNAdvhLJ+E5pWvsdQWVw33SMJztO2GNXcZqL/m9+N3YTN/zswr3wSK2
DFUvNjW5b0z8+Jc93s0Kus5VEPVVRLmVZH+mmJ5+KviL4n3//pNP3ulb8ZcaXxprmJQDYIsxSk0J
yKFvLtMFGh2xfso/mocJttqkYoc11igNIxG10bKPladlANJv5P0or5SJhXJMxgs2EfCoDfrGVvjv
zUOgYwyn1W9UY+bc4RyPB3ZWQl6KbJS6E70AIPcjiscETeKwL4HxRfzGLHBhT/xOwGn+OoWOYW2F
txIm/90ZUb0Q5CWmXbYAuGjhTOqq4RJ9M5GzkgmIQQgrmiTVSibg5FUM6J2WYU6d9FT8LvS0WIcq
tA26cDwf5wdlY4lB0TbOjhd3s07QeNN5FnuUXdH1cxK1TWyO+4xMY83r4VOfA4HcTj62CNTawZY1
qhcCkr29cF3Frsov/iLt/H2cL7NNwIbuhxxqLjSbwvHnavNH/xHKBckain21qy1ORkPeLrw28jIb
BFhJMEVFcQmG2hJMb+qlPfTcfqwTA63Y6g3l9gGibiuZBqWBJBmT7ewo1RF5OuckPo4Z/0wt5inc
UGqPHRAa+o6yp8jvWZloocPwiN2cM2Cj+jPckwji2VqlijYY9ZvhceLlHqzYU4az+wIPtLGWLvlH
rBSmbXc4eYR/OgVAj8Knlg8rl1gzlx62+Re0nQgy8dksoaXDj8EUpJJcAuqXHgAu5iVGBaQ25mTU
qgAbpLs/t3gYGXaBaTXV0zWr8nip/Ss59XA1iQSdWqNgdQ7o/JQZ9L1wZUc9KOJFnpvad5UMSgea
yF7dsTCcWSy/j2ZLc1bPO0LZxUDzV/RkT14fpbIygCLTidz9T0Pu+NR7cORhY7WB4JimMdSRH+j7
2zP0zVFOsuJhTVgLgnV6zaJA1C9J+izFI8vkwXWzPxitVj3eWkK05M3VD+AA7rAmS2wWNr2hBxjK
SfbRAQlhIh0vVP8CDNiaVBOgGOXXtO0+SqxM8f51XHb+8AFakJ1pkYlsPMW+9FdrfdnxHPZgBqjz
eQkW4Y7c62eqIJXUmLeqO4DBGhgyAXZ5Urv/HeLElmwhQ+NLPUL4j63O2sJBu6NfrNSJg8o1lypM
mFZXPvwO+ob0RYGL786UY615Pnobh+57rUCmgKFHQdtgz7hqtnzkTnfqc4tXNBJLWiE8TYn0OuoK
k1c9B7W95gV9KAoWVlAw8fRjIWHVpCYmL/oPEC6v87AqD6ww/Y74jPiNfTlLY0K+WzTu7FJz9Byp
6K1RVrjXoHl3H6KK1TatyuY8Jdkfuas7GLADVFlCnj3kXarv4ftsbOPxefBDEe6QHYhEcJcx1qIR
Y2YNT2LqxsYBMKX762Mts4hnfZFtC76N/ulGmtSl7qrjxOmzuPcREAb2P26o2hBa55svAPxi1BvJ
GmGy8JAdNfv50QMRaWiInq0/a21X9y2/Ijx878PXfBvOuuWK9zf7mxVH+o5ZbGR+Ul2DGF7iZsPn
eocYSJyARe/zMeSKUYIKBIkMkyR4B9hjgeyXPtgn3z2CKiPeCDDI9ut5I0CoAyLUA0uTRIMJ55AI
qxXg9yhuw1FA/MZMllBbfzVmJRuDR8eHXZP9J9h0CZqEBL61dvDy/Q6T8haSpMwiKvj3ntApW3xZ
VSN38Xbx/HdTSwJFcRwbOpPJIa3VDj/d4amK25dazylEyFjJ+U7PvO6Xk4OOakZSa+FdMd1qT12i
NuhcTm1fBKSbmgilWnZ8Wmy8UT42RrZqBaGhp9FQ3WTg31/1PS1kokPVTc7tkySPAW36v2xSBdJx
CQt4SDDlRfoBshIUGiRz7ieTuPwXEwiMvPi1uWyLqdJx20ZrK69sEtXksNVCw6Lr/BT931SMcal5
hiwpfaa+aaOdXc8bufkGY3eooiP3aZ4kww8rF5ARdfESQLMp4r/WRyF8zT6upPFwbn25D34Ss768
mIYD2FH8zDrlbNPf2bxv8YrFhQ5awDBqb61ZYBMbKW4DL96wVeFYxOEj3eoikFnauzSHIt4wG10B
wJYGNqN26eZxDr3/Ubks6PcQa8GlZ35g9VzErshjGDTNDtL290a50yJpJMZqScCEaF69ox85Q6nN
lHPzYjVK+gypf3FiGpepeZMBRbQ5YI1VrLh4wJG2/ClzDDve9H3j5yTRXTUcIQbvDYvEZRGVZNh/
i4yaUfKz/hLVxwA05h6GNlu7qThBZDObwWiKCVh3DRcLE6ey9JRU/xpJXPUXN8rKzBgutqgIQe1E
G3fDZCqwYtkps85mL60qJCtwQutN238VG3Jpq29abnOq+TQnNbgbkZrIh0M0ZibBMmcGOvzeJDnA
GDBe5LtmR7ZY/VFyH0a3P+gfhpEsQ4Sv0JxotYiwlWtWHYxKKogaEB3+U3VhaBUTAcQBiTlyHwu+
Av76TK6bR5pFcCxlKpqs61QCuK6fJokfRV0a8t9A6ZzUv5GIE3XYtmQk7mex9kPVOXEF9XNyEkIW
hznl3mMphy2bkWBaAZgpI7p/ed8MKXn/w2eDtPnU1ezPbucbAc/bpFh8uAmMbxEVPP0kvYPt9dIP
m4Te2e4VRs3tq+hPgdXoVwV4UOv8bl94eVnNBUfo+qmFToFORzAV2dEzfU+3XDmmD1//lpGiM9GV
m3aGy3Pb+pTSpsaBJ2KLoYJO1Oa01Dnied/Ye52Z8nrfH1bsl/uAXHxp9walSGY4kJtEoCX4Fkuo
YNF5Edn4GE9uY8uCsBkejYjWMBv1jJQI09GrKZpwfLe319gqgg3WwKsugz8+qnKtxbXPupmfkrUU
m1sXx0pg4e0iK1Kabjjww8amQ11CtF8MxOTZyN6uwxmJiW+ixME5XLk9dOK+tlEQ8vLx+Junt3nK
lrxrjO+qP0vHrSloYZ7IKLrBtAzG1yTkPLnn9KMPvb9aNqgzE9voLkjvpOSsz+4eQnEaOhKnEckA
jGCZcU1DjtB1D8IzsroPZCKjhmR1zCVp+EbWodafbbgvtkI8/+coFcJq8Z+MP9o1CUMgo4ZKSUVM
K+He8gl/8f8ccwLsmgkAj1n2MZZOLZVJYvobHxAQ4W2W5XbGiFIQHbmprnn8HupPW5BRMoRKHvGm
NgzJoJ7lBx3r49t/NRRP9J4RL7R1H6oF5oC5E6PnsZlkWjwGR5Kcc9Pgl31dyUaFl8KjUvz/mXEe
hGX0BJ84pnbFiY4tTfUva/pchzJ4RRLheiNEbcerQaEGUmMFnjVvPyv5Y4kVjmf7begrE3YzIWnF
lNUWYWk6cnAnw7TfYBGps1MgzO5o5nLCgX/EV3PwBiLL4HsF5Srj6ZUSKoC2SV3GhUSVMPScGAGU
n+cDmxJqSZH07xP2ao5tEu0Nyhd/AUSTBVUUit7HBFPVUJDkbcPXQNOZdS6s5AtxNxA89N3O1sOp
v2BztrURo6r+u4nljpZba91KWYtIcwmekk/Xhnq1yoFWLTYSE+UmxxNOx6p4pn8PAKAJNfdJKJKv
Q+b7ArfHk6VEKa3n9496wmIGUodQPogELiMR/yvlL70EQBIM6J4ppkVQwKTz/jtPrXBotIJJdyiD
Aj3tZsihPtKGQRI98k38HoTUy4SoqazYHAQ6u9gqmPEolfhbhfb029siLMA2djP390kXIJ44LpR/
BtghH00rxHufV0y8WDh6cVzzvOBWbyjVKVNkVCe3uPCcR8FSrCEXIRCNejaBgNJFMNsViGhktPHs
SucFv/YBh6B2krpg1NZ6iFf4v3HnNYhFe0rNsSKUtpaaccSFC1r8518Lj0p6tAbWnVXYPiRdUh3M
RxJLc6u8Enld6GDd+qINNxOqTeUUtFFUlZa+7hHi5+VgAeABpjbOqrwGVTy250pNm6QbYAMfcMnx
cUF2J+RWjW6+B+8PFqQsTtPUIIODTxjX94jbw9pbTaR4nVJSJ5jB5phgmcsyJgAO26PQIVB7g3bB
GqJVAEX9o7yv/fXNUbDOkyciIPaE2JMsJO+fKDZxOOX5JkSGXF78y1RLub569brw0FxL05+4ZEdr
OBbMormsmRIjro+b/sq2lClLQz+McsQG7Id52mZlv7T+9mYJJb66I5ZhMgMa7lJd15afUZo3D8MQ
f0PCGCE9b7MQXYvUl8rYwcRRGUtF5YYcgppCY9BlfZrZ0A1SnmZOT4/y+JEcOBkbgcBohdPUwacB
kisPghU/Jkl7LCJucLRCz9J9296PGgI3+Wcxmt5gXsNslhhDBwAzg0Fj6PKQ28EooVCsX9VrtxEH
AkPbc6W9lffEf4O0rKr7p5jbFeC3DHxlJPLbjYP00Fq2Cj6jjmzh318NZcBz/ttUZfG/Lb0598MV
oftbr6ijypuf0U9/F5/6LK2/T0ah7ysJEi5JTRA54QdOXgKUJZBK0dEH8eMpFQyJClnYGXcSKsQc
pO9Af0DCthFCppE1991EYKO+r7OP0rpcKu2MzYcOOz5z0o1k3eTn/Vku0AwE+tXYvNI/yQUnp/aI
kkq5FjqY45YTC7gyvkwORQYz55s+kmp6oWhsD4sRCpyb2Q69xUr6+0nblUBsdsgnROeIyyBSSx3D
429eTPj2RXnmf2rw+L7BBSL+g3E+izRiic6nyNvNfenKxJ1prel+fz9N5nO0nf7XuaCylnl1ikAV
13ahAN+Wyxbrd2kbGB18DAGcdZpba2CNfC5KcV56XX88CYgRaMlvTinkretF0z1d1lRg7UgpgoZo
K5uhu4CxxVUYazTwtTV9TEpO3W/GOxnygYtLp5WWEHb/EOmfZY8zJL1gtMI7CxEsqeVHAAGg9ETt
b7wjSEVIgSPrUAsnZfJdzybd8svVR8xUjciVl8uVDZxjjKKJjCqV1bpK2o1UkWWhI5GM3gZbcErp
CSKvYPEILK6rXHHJlDEiU7Nymnsq3V6NcQc32Kub8ZALDWa/ciGc4/fdJKD7ADg/HhwjEJlNVdyL
vUDl6KoueP4f2+mcGJBLWmmGUUR2ZMBhMNY3xEpWpmK61gzXWHxa5rklSjOVOdN7GI/51oSezFrD
ARtEm6TYePz15QtJNN3yXvlpkrTcZXxLaDKI2UycxNTflQHFETQiJvdJPDDCbUyStYfkF7RRPPJl
5PdhCRJaHBeM1jShQfMVFtz8GLB5NMR8TBq1B7Wy1wKM6F3D67D1SyYMxtvN186RHU9j2baDLmiR
z7UoTcD8WIaUeniWBBoNwPbW4EC1PTZ+5CxMpt3NPE6QFY+FECDerWT3qyy4fQIFkdyD8g6/BDEK
EV2jeJKXdTuEo/qFcKqrNSAOtwhma0Pvl/5Rv8JPoM/L1fAoZeIeWyxp9XgX4sDDrw6KHeYWSCI/
Jd5kjhXNJ1Gn0EejX+FgY+AKTM8XLn5Fk9nnHejyvH7PL4wJvEH4vVxaxaDl224SrXAtdKnk9LBV
UGq6YOs4yhw3Z2B6xriQKSaQTYxsK8NIwIR6zfyWDgmrD1bsCnlALyxEID6Xb2V9Bb899YTaCq/v
hp5qlCGeJMZzaZtXDz8VaZG78exN0ABpuUF9KZkiH+0ZuBN1a/MmYugHMU0w9t+TYReuUj0Zd16F
efju6xzM7o20s7q0FOjsnu0bJjt22FFm0nlT7W6L+AYUrZDsMBdYwwnE7WXil2maupcZ/fPSeswa
bFe9mIKW7xTak1oLDHacC/P1jTAIEB6rD2wuMTHMT1iA9OUnvEylDsONmKTjBLVgVq9fCzeHvD91
fXYXh6UY6XGJlX0pI1V2hTyO/19gHVRo7TSh/Sqkol40MJpwEncZwpJ/C+s7SOQzuWqRLO5KEaxQ
cQJtNHwqML/1xYwwYcms7SxxgCHsFHrLVP0lnmJzZNk7KK2lrMHmnlRVKi1cr1sWsbwd9GCIYQPY
R4/NWrIMdSk6zNVPWEwR9K3ZzqiNTwtrWAZJ75GlOMUXwbACHEf4F7p419VwG6nMwEIQYrndR/dy
vVHrt3JFx+US3d4KusdForVXxhHXcv1OOsPYgbERV+B/dIy8siDbsq4lc+HxLeVps881L2w+QikN
VTaE1wjH4oDIdq83B7zeJrs8ElMxKyZXH4HNdkCgIBNYUB6mwHfU0IfOwI/klmS156xV09QNqyFW
gIaRXgO9uUchck8Uh2JXFcWQfaSd9X6bVvUVRAt2gs9SZDlMYmjDKbn0Azflp1jk2VGqulLl62uJ
ZogGAbsAFiNNwPpN+67gXnJxZBzuJ56NOINIy9p2pK8bcOWPZadjCn7qQZa6sw4BkrO/SP9U4lPG
BKpEPtdpw3+afBn+Sqblz3fn+pGIMiUkp2mEEifeJYFCsEEiEeGTFIiaRCbgIz+wae9Qo758uSGc
2IZFamjnN9tbJLQOmrpGhud8hvf8NGu6mAfxAJcOIOyrgdoch6Yx582avDH0AWwk47WehkKTbAn1
tfN9/ntUqp1cLATnxl1cZRHLpa0Qka57w4TiyQUedACvm64Zw3f5L7tFkWbuID2tg9DOupagcBJw
csIVXde43wAl01ZynCpGZ+RTthfnsqhHMzS/GZwACLEKHNCtjPdt6alD0s6VU5snn4fJU18wjbHV
K2gXFOsl97fzPGxJ0sG6gHZQvrsYuz33EAmZmOYkv+ZZLoaQsJ7uax9tdSn/SQtCsa6AjXqHvBCr
BBNEpHaTCoGTwzL09r5nYIFo/rvnmEw7Rn7IoG31+TFYVK1WoJm2644TlIHxfRGyvVjIc6b3okUS
GJ+bQsOj9ieSuiw5hYJKACAfultYRYVnVf9l81Vi0YYsR6mEogIsKhigMTuweVgrSaQvDtAKDUpt
u6hhPIbmTS+pq/QUbNb0ytoyl2JlUd1lk0i7isArGoD9lI/0NLT+giUBMh2kDzYXUEQtMtzmeIne
0uY6qC/R9XTP6yIUgg6QZHn0JyKNCSjajylSOG9V/h/aNn/kY05t1bVb5jik/BQA9BuXHpw8vd8y
fP7VMCOiZdvCgmC7sGEJwRgE98EKV6u530B9Ma6j3KQzj5jz+Ms/PgZZIjTfcS6A2FIBc274nNCj
J2mmNFs0h94kUGQ0S8eS0BGMjXqUscvMzgwb9V/7FS0HZkPczyoEzbXdyp1oB0j4pqutWibNOCmC
9KTmOvQ4/rMzanJ2YZx+kVcD6cG8B0OCpAzg/SY4iJIYhaAL+yUG3taUhDwMMKHiV/ZGY7/MmPQN
DO4qRbejBMGsvO/D16VYpS/vxs/5ll5o2vYT3c0u7YX8Jk5duuws5uMytJWs5gN74QlHa4DrviE1
EdewycMtUQKl7TLrq5v91qNm/lE3GtVHCv8o3v2yBnq7O6gW6fqJma8rHIhUOhrWGQZ9SZYQrbZ+
SVqjkLG45d1TkxT27ObOvYGTLkH0MdwcFC6JUPURY9xJDHE0OOMy1MPj4RgEdgafDoRPHEQ4QClm
rJXLiuKLh/CgJd1NX688UxSxpHh76LNLOqgyhIZPgyBHnqqMMo1qttW2IkWW2cYb7MpoW+BkSODx
x+v8KDqKZ0fmqPi1f5c8Q9DSLWn//RB6wdk8SzLoqexwMyfVhRUcwNGUEEVniDC1OdME5eGfwlhl
b6UsGUyXzbxXqduU0HHqJBu40JUiNDX91RJiCv9SbaEcCa72uypxeo1Xb7+1+tOQcgkiLhdjudqg
/8ClR6HmFhUaYtda++UaLKBu1F15wtWiLWG9ONXSyviyA/6qRkVdYmFZIQA4nHSUoeBu/+GP4pDw
GgpM6iUHnQP1poQeiDq3oevjiyzr0QjqDMGJSsTkidSGapxHxU0sFGyrxlAxSlfmsZL7k2ksqKAi
r2ARIyE/YK7RrJl+Kqw78EfvRChXiM5N8AR2x1PkMf2VHeCReIK420rj9NpkG9GNaUueWHBjVaVs
Z0whpGv7sWScsDrkgf4xY+0q+43ipRTTanUxVDHRuIYYCvlU/eboT6fHv+Oa9vpPZltim91frqk9
/rpUhgMdKYrujUCIirqPiZbOPw4+F17wgelvb5Yec3ZjFyQdRAo61VcyXg9oOKWbK2e3xBRIRJHP
14DWTGt2CicPdc7S72wG26zHK1sJEkLsvWI8EDbtH1kkpHXwH9jA+kLp+97b++wI58cCs6D01tLs
n/i8eS4zYTTToVeHBA9mcyCGVzBK46LubVhe14RoWIma9h8PG0Gx07jZj6HLc6nP+jD02o6fePGR
s+Twyb/vHGhY2Q1AR2QszpuO41IE4RqfTQ9YJyGPiiNPNWRrBupB4EPAZYyl/PDmwyJOBknIVOdn
d8FUQ6OtP8hcTX/o41e3U67u9+cKJBjvBOoNE58VLD+3zT46hNAyHP33gff+x84UTkeUGTm7HNtn
gu/yZFH4TRsxgL+8kAFbWnaNBQKv+BOl9X5OFOmHwW3OuIq4y58FY9eBPE1DCtK8PwOykEttPbv4
rcJxm7fpCG31L4pkfL89lTOMMmtAcgB+RVUcotAIIh38IVC6Rd+6UnT9igIYlgXPXujGwA4eCUn7
XfvMOsZnePSVPUnkOLpYAdG75eDWKavSxnL9MoBpStwRESFlqKe9lNSekbXrUE5v0p3Gkk9jmLaP
TYjZDaUddrNBpppEamRHNT4KSiP8V4N2geOooEuJQxqBI7N+PzDxDFWTmsK94B0yp2gUtvv0It1e
FC6xa0jj5BisGQtcbYh6ve9BTMskh/T4pxj0hvZvomdHw67MR3xAZJeU4huhpjvb5IwXDPdenL0E
geZZc+8k2fsTnCfP6URiqkdWPBzhxRJTjBwD7ts1yrXtIo62kqTMaEwGquxJg9oMe3EwtfBRNTmn
Wz3VQJB8OZKbYnEMGDc+hScr6uwCrpfPoR6P/8wVmdib5ZMYDrY8xDzrb50tjrynUTL01rRoBIrq
D/7asWPJj4ZwKlktbutIOcxaq7akNI+uDC13vTEQ92RHUyiKcbv3J3kx8m/tTBxkPqz9z6RlOOBS
SAm3xSPKyvChRPlmSYOebXhaDlrxV7/m6c4HqILLyqJsvCICa+zbLAoGMrYVERC9D52s5B+3iSm5
N9/l7QwzFbSbNM4RFuBYHwb5wwwbzm3i0kwqUplRUS375HL2mjQmRnkz1sVWnHHcSOKV9hq/wegd
EPtCOdyeEy1lpBGvryWmCuVowAY7kq7Mgkk6fUv6Z2nT8IEspTdtyKNpLIzMWACiKNXozvYkbn7d
bdS1brdKjNczGX7qbm11iHBANODYDySNagILZFxhemS9LF1Q0Q5TS31T88Xw2msO4JvurICeK6mD
R+Ss6mwavfwBbBGiUR6U6XukmRKhT3Zcj3ldi2BuESNR/po34U9SmJtua+oKpI5SPWubFILj8SsX
oaCjrbStK+K7Wql8hiTXpnwdSLe+D8+9jY4Y7V4RL2kdWRZz7TmBTAy29WRLJmx/gqT8nDrmV9Cp
pj6lYF1b+XpG9oxyHWbSPpz8eyccAq6mQN6aQmhITg2GuhHYf4GImqgXbQR94RQ50WQsXIzpMn+e
i+V984/Qg65nTGRSpH+Y4YppLJr/x6H1nFq43H2lkEHOSFFQLQhjJwhes04fk8cy+VdsTVicfDHk
rFMdZzKOg+Fpov0bKyNXLFPlmo/BHOXsJhWwVwuNhG8HbguLKW1LL/eLGuhAdJLHkec6NSfsOjO6
GTRBfJ4vbQyfl23mUD/1Ek56EZfC8bHTEGSqWf4Y8vJxXYNhCapXBpurnSA0v192JW8ykGVN8+kJ
v4mTZhyK18d0adjivtN8jPUiRjMd7GxufEmP+lAk3rdbx+hNOUql2XsTIde8F2Ii21Kqkmk+hwjb
+spiEuBRzEagVraX1/2WGvG0WGs5Q1qHsjc/y0epQf/ETLqpdcp6pNTqsovO5Rmx9BwHIbhhYff+
mE8e2NCQj/2RlDw7fdr5owEWh0GI3g1YtH1KtYzzSJRkhs6g/TXsMUcsktIIn7NvlAJDUmIpWhYd
kNT6vbKoQyuDHnIBbRIEJwxdzDxvhceunRB1BzwwhKSCVpJdY3dz407oFX3Y7kYr3YTlMucbRpTV
CZmQ61D7HN3XhGy0oUCO4kJJ7e3ZEvZeo2RaAwq6u/qwwi83OZ3fyswucr9j5jcoy1WfmPmh2Reh
p1yaXNTCwH8PJoJ5sOBDK1PIsf65V3eA+Fx6xcQN3t22AOebcd/WcTWAeCPWbBBK5lwdaLbyOi9I
8J2+GjNHw7Sai0FwIrQma6txzyADC8FYimHXvXESO6vSnXsAZ02RgLUZo7MSUabLxtWxlIZOxXHM
7hUGNADbHJiz2hwrLTZ5+lcvpbMJKn5Sv9PEiOUIgW9oLR29EsiZCT6qxKN41K7rwVmAuLjIdcOx
tOSYXJZ/XhtghObrswQRS+jS4NesXtejRHddeSVTyuk54utLp+nATzwRP0kZau9LxroFJM8uIETG
dHdx1hoSgGwubDcC+zSzm+eBdukjrE5UhbW3j5Kfn/LyUCZC1ChpGMZtrmRYBjPCLSJsgehl1Hje
XHDhRKaZfuJBNlCMUFD11SckaSeula/R+FYh1VPaaERr0i1qUq7zD/NgKBnbW2DnVuuCWMYrQooA
LrBQSa0KCdIBwHXRDJGXr6olam4DT3OB8Be/nxtzD70VggGQCKaPvqUkqSqOnYaLZz+yEU+uTePr
M2Bq5SSMwpfV5KoCQh/TD/o2vZdhygJ8m5KAuhACOKS3K/+V7gUSj3H77YC3n8ZZl2Jh/T8Macp8
K+e61DJuDTll2V9hWqKNR3DEHIPv8CgzwnW2xLuAbRCGIZZFXGJTh2zoqtfYwOT0dO5D29JHefR4
bN4edw0PZlQf0zW37sXJU2lEgGwmxoreQfXupMjCU4PsUBhZbl8pIHSDCFAVYv1JX7Sm5hy8dcah
GhqiI/8mymfQ6LIC5XMYBbfXn1cK/7V5MNrbVpCLlTi1QYRji7GbBxE1zVhXudXGrwVX0tjVAeFt
5rnmPtPCxhkdqAyjZ08N0BdOHwhbLWIvS0252TkKgt8DIBIyft0mOymMqir2rPxnm+UleEbpnJpR
vhEfhMQ9CXduA6P64ogcjRPtEhnerUzvcVDQm8y253pMR6pzpQeArymAmkdC9LC/GBAvU3MiNo2S
8CL2YTIPEHHvcZZd6pN7lSaMhZUN/+OZe8w6qvllvYWEr2Q7JdBo39+iDKSskbryiIccZ0b97tuA
MtNcm/C664WAJabLBRi3HH+Sg4fGOFfg0mIlnA6opNO6P/hSU6vrsW0CvcTnzjddl/OnnCgMJX7x
CqREbV0vXFXDjtaq5xAv/f8L5IUNsgGUI8edjmjsK3SeXI7mEnDywO6Q5RvSeDQBYjulCbP78c9a
0KrCQ5FgeBOswnhRLKBTqEK4HbAIsaAFBV22f2BNjwRGBqEWlUlUYb7rIN9HeIw+1HqTMyOGG3Kp
DOJ0M1RYFQLI42TM/NixCxNpFFknob9owRZAnVIogTuYF/oGl4Iop9hOCh3LhMRnrHZxekhaiVvu
1NAVPloYN1dGS7LwUo9G080qpvy4FeDwg7LO25jkYYtjhZLi2tP0pUPhM022r8QKIoMjpvjdrwYs
zDtm+/waojS5reMn9NaQ3Uh8Y2BljoGjdSyTNobkHuxOytxv5RrI6Kw9QRnIaPCdGrqbw8+i5lxc
u+V45t7a/LTPGg2ZYbywGTeVO9+6I8npYs2O0mUlh+zLZliuH8+gy9zbDSYzmGBrhUAo2FkfPuEH
yVBPNFKn5mQHjpTZ4up+6qE8uNKPtWkcAbhCjE0NJhWpnScsgavdEq+BrAr30ZLcTHRAuiLnPXD0
0vwNSm1RuQLyu7Ve/ohHN8jJ0Wu1ZocAPJ/taDltCX2/t0jMHyAIefDWDpMY+g4xWcUR8wSKjY1Y
2xhLIsHIcT2eNrJo5iW4QdHXBLNQEPev+d8qCwWjcbVzK+F4BF8cC7r9R+iV/8wHJhrSIKR8WVRm
pDRaQ0MlvBko4jQAqRJJ6uMhd6a86zH8C2OcJue1nSLLT9nXN1vx5zHNpDvvpiUjn770Ec666/EA
+Xu+VSvtly6YHdLYGg8qxH33VqW/2flvAp23FrrHS5wkHTOF8YlY4VQETU2gXYVJ8+Mw33kSSj3U
fU5xTeUkT12RehrFmR7azk0vO1RRa+6f9SQZVcF1KQr4ChUCjW/bCebXgzqvL3qGL/JS+wgGFsxL
Y17ggm8NdRY5m9q/0Qixx+vlFYUnBguPuq+1SvKBbko750FH9htumVFW/GAofxpZjLkgLnFm/+/t
r+1fr/0DWuQgX6JQJGELvzyHEYxL+ZKQs/4QPxyIW2R383oBSq9HNXG1j2PKEggPvWoMRMwQKkZK
BvVi+9kNoAdupXeqA7iKR7AIIZvLIXSlqikZMP9bwtolskLI1hjYGZPLw/vOHgB7+nwrhJdJl+KW
PFog/e/otUQBOtWJOPEmnhG3GBdk4i46/IH6Cy0Qu2w6OnycJlqY8+peJ7giz42a3I+R0AfwWbep
vWSmS9ORCh3mk5FLfXimmY6vK7EFkBmxm4iC9B0BUzO+NgFq+qWcuCSoWm3MBik/XvGKVP2VYKK+
AZW1DNJ7ANVmzK/1oIOQurZK6TyngZcrIbUOkAb9snndov3L8kNq2iKitVPg0K2YN31Ua6D9kGH2
xDl7XZxucpDMUKyUAFtnBONlCb0u9vLIwyFaF3MSZgBNj83eYrVJ9BdMsVg1AVLyqSxvBXHYnj3m
0XCt9w4co9Exg7ByKYdu4vKxrp+a7Z+V3zNnLn1s241LMv9nyuvm9aaqJwai3/gT8IdcWU8x0cF8
wBiTVfWABjYRVTWr/5TTxYDeD2YvDzF2rLCYFiIeJ4u4tOJR803unPkNSAvo+bmy4eSl5k/dAWJI
kDpIV1ytO/1C9/J8LpLFIRcCNLuiNZQwrDvc1cruX8/Vq+gajcrKIiSB5oXlByxt7zDW9xps+kvU
7E97ZUbifHP/xkWJP0zak101QR4UR6Xu1lELeb19B8aJhBU6ym3CU230iiwo+pObxBN+echt1dbj
J4fW0tK6GoL8hYdmvnxmxfceoHQqeiw4bIAORrb2yYKajaQVg9pW/YtJOlMB4SGBiGDU8E+PAkXh
OLJ26HFdfnNnGe4guB8VQtPRXk+piSPYiylxZkROgPAZcudYYlIfDXWzngf3JcPe4nd4/UnmXMoS
JyrNOteANJel5Z8765M1K+uH0/o9ttgpvPz5pKB8P3rzgaiezCwsDC67RjbXhuqGOSycNXAyt2BN
Y+c+sG+5DSviekCZc1+mENKbpaomzACWbcmVHb/6EADELsYSVp8Gq0+7BJHw6c4W1yX596vdrrcu
l2IFo9UUvJhxDjlO/6yp84EJQ2WqbSweuKPBU5MJ3m+zACjTMlRJZfJwBXbpjgD7U8hhWhoNla2Z
vDXLm6Po/a511UfMx5TOnDzCeDa8tPA3FwR0EGeE4FWCqv3WJXNngCP7e3mC9fpxK6YQB2C+RDnN
kzY0K7eI8fBnZhCv4gxWOTzs3ugf+DSjbFnO4W6hC+bkVpZByDCqQwSnGaARyvSEjCHuaIksTOkq
sIFLo8hICsNW99SSDUFu5CV8xuVfJTlBfv2NeX4Q07hrj+AzD3KXEU1blRGc4JvQXfQ31GHWXBT4
7XRsfonzHekkrk50Ju+qbO7/ufQ01ss2WBj+7eiHhelVw6ZDI2DKD3GxsNoOVLpIhk2/Gj9E7IrX
tl6bS+EUmHs/OvKFsNZen4ryKRR2tUQc6BiTqHV2yGkxPx/M09hWsz+BeTZzd2G5rWUtE5icOyAu
flDGDIFxi5gNcCKyWE3t0WzNRYFX/DmOXI6xXyBuWk2gt2Oz2HLVASDKaW1mpX0ARvA8L/DQUDFt
WP02jLT1S2iFNzTWBJaQ0smkGVVwYrdXgtFHiW9qrmY0BL2AU2W1ij58VrHoD8dvh1oNJ1Ac7naw
GwpQEua6VI+Yws7NPAAUjm/3lf9lFyddjjOzJ/ScEfKB7XCT76XIlo5wBRmTdp2BH/EM8WgdF4HH
Uz3dp3R8/sYVMoXSBPPdt4MfWApJf6LOOIheX7sZgJ/zRlVHrSQZh0aJAbC9wzFvx3ZxT354ScXj
IGVJNSMwM5vYvLLfvluH3yVk0aflIa+8FWH6vMJ9xKVs300yYkQdnBCBAT+P97djuTSeWHAOOj7I
DA9K4IYOCuzgCHUIKu7U3PWs1hkBPhQxx2KyOR/mSBvuOrv/m8FvQfuIeBR+F5Yimkwm8okOkWGm
WRdd1mNXAvvaMXXGQHRsACzJZhSn48GaMr6wFU+OXTfwDj7QO21y+TiWmr7XxjKSrtUVDrRWv6/L
N97iM1hLl5bPY9LxC7XWM8apPpyQ1cNRr/umfawrg6BD5BvarkJ/ISfiLH9v31q7KEcjeWpshBW1
dOyEcu9usTBqV4mSosaMnKqCiHFAHEi1eK16UnykxdYeotloOoZF/zlsyZmNFVT5BM60VcHI7ZJq
7fj9i0DFDhkTylMYghzJVLWawX9rhicw87Tr0ikHgVNqSxQU4pwyLgkZL+npzAmY75yTIlomGusQ
ZNSZSHKLjc/O7R9wzds4hG0AD8szlG8LI5MHQpJduDTf+4REa3NkqXKN2pETIu49210wx2e2KhHA
2Om66xku3JIFH3BLTSPYRVS0xHJKfKYPl9ckH6Iv9iK5v+14jHLly41vTj/i4LL4ebEbIiMXgSIn
INiyN/PJFNyh4vdKH/802WLMzJREpJH4glg+lk/RplRTYdFYuHIG/FkXRPiGYeNpFchC/75ftkFa
IKIMNzxXrxvG2Dj/qm4E93JnqLCYezfHYzBnf2mVm6yjGVURs2h8j3E7LE9IKxY5ui7REBOTXXqP
C3t1CAY8O5Wm7wUOJtTUxleeyJNmMJ7YuvJbUT5HQ4uIykG6+9THu5JfCOhCpA86XzUdVyNPdUAI
695cfbZPbhrdxp3bpu0AKZkKXioEM3ChRzaIDdFCotOeJe7XMRwF2AkDci8VI0i+oRFrFWyoVFoj
mb5vUMuNezC1D0rNbIxLItvmQI3grJ+2/IlZlLwjv2vabYqiBQF9IPOwkP7Hk43vfcr0Q2UT94Rt
lJMBz2SS7exg5+FhAxcM5BdLVOHvl0cQ067coWQQUnukq5LdoQCgWUAbL2ykremqDtW0z7UYW4jB
CpHa5lFWjs2Rb/7eXlyPUGlZK2gSFd4/YzTTVGV6roT4CerWtdYePLr5pMApueDYuMlegqR+ngzq
2kdjm2bFPnpGWMA81i+zpVuRkqqpO9ATfXe+rz+5oyaPDHXoEJ9enZAMuubujk8l7XbUGtBYZdK2
iCgiYbHZrJLS/I68FWgGpJA0TWlqRq7X0WVQDwdei59xn9j4cTzNYvQTUWsvaOc31KAMDAUxh7df
wczna2TIgx7/N9JOne2MSaGwTSygx/9no+MeAsGyOyiPuBEHHYPAC24yhfaPd19+S+KOsnu6pZBs
3wzYUuKcXiv4GLOEAzEZ7eRDraDleHlfcReeuO3RzRb98RsHU+jAyZ/2zuQqibndw1LDgx0vzFFc
MYVmpC4eETIAGwyxLCsMXBlP7EPNoUubzIsKF9KKjCn2QniO3GMCpWemUt+0VDZ/93ztSgjLpefj
J9eXnoD+67YAgvb8z/3e4WucLW6iujGrgGohe7cui8j2bA+oBsuTx2Te8OFRm+RK14GwADkFi+kV
t89YsLBvG9gpawkKYvq5C+xeRWaEB4AibiwFEqZBXLkeMcA5w7Blad0q55WHKqRUL8Ge7AAD4wQe
qr5wMNHb8fL99etVZP0hUpbDc9/pBLaQArYsjjKDn4V54AIRZEg/CUicyuKU1+Ceds+xWZntIHNf
VpYqrHdrVuaWWemEEB0Trdf4ceImavYL5g8I8zplFFLqO3W9F+UpKyw0lE9mk6kjyO7jX68TjhxB
H885ViaTXLMk78XdVoRvPWXSclY5kLH60CzxYqP8i53FeeBf7b4BnClLa96QvSjON0LwHaz/rOHU
tMQyGMx84PPRZZ2vYT5RTBDOlOEW0PF+VvO5HY2xD4+8+6ol51z00iFL9qyQq5DyzlbK5EXPh4Cj
dtE8jyrKIXznv/ATkhOZi58X7m60bhmTMC79y9TEu6mz+F2LEzs6IrTHfqMBHQNfK1Z6uLnkynAB
48xjd753evaWClt/rtiH2QP9vFr9wtkMEIMtvv2aVhIpNxRgIDnO0sq5WBDkYTXvLMyiv4uckJYa
nsHyESDGfyQlXKYW9Xh65YHCuGWrtiExv4CEpEDuahacPwFVtbRhh0YIEg4MLFbvnNvMFO84IPsQ
lL0SXBhoW4wdqtHavETfp/fR8mOOj6t1J8KZxBDIuL4tT9LmJvwaK0HQPgYnidXLouUVFuWBTbdX
QzX229nDbUVB30I63Mm51Oj2FMS2fVsZJ1qwhXZ6YUrxKY5Y0UfJSOrxGLoOrxEprdKbsGGAQL4T
5S1iabHmRHZQpbH2YrzbNIPS/G4PyRFUtVJF77cz2Tk/CmYvJHg4r8iVg27ltMf3omR4ZG/CHm/k
GgIeywS39opJr1bmTxsozJco8C0pXFPDfq0Eg9vrrnGcGaMJq0jmHtagLE907pRX6frQ+CUPPYVK
tNj4Dt9/rfBUQKcvM27zcRS4RWsJnyRhkQfZXduaOSBmdbK2g8yn8umTg1kfsK2iAL7n8Vyax19G
ut+RDGJgsZY3ektkrf2oZTwK9MOLGyRVOl6C9Ccd+4k3sqLHG0NeLYY3GWFq+Zx2Pxb4T2Q7IBp/
6iNWZHmS9Lq+wj/NYdAvHlhaNTyJv13KHSOBRdkLqqec9pyCfyw2NTAUcCMbK54lWRHu9gC4KlWM
6armFATnO7LFD0F7MubcqdcBzEeTGCd9rP245+fkhyl8s4jDByiT8+WOr4VkzLoweZOeDdV6mE5G
6ebljEBBRLyogQj+JEeBHcxsc0rkTjsSri/hs5K7EapSFKSMY63pJTcyp0Sr4O8wx7lFGcydJx+x
gNr2p/w3ZC3HduutPGgCNMJHCzqEYM5NSZQOcShxIrQ79wpyMIT5WnjxWiX2UgOgvJba4HQzDCmy
gsJgVk6K4kHxibxtuTn3a2ZU9J/rs1m69dTxRJa3fIhos/utcbgUCR/vrbv6yRo4bevzsbvRoD7F
BPWE4UgieUBle0P2w0Gv6EqxCquUqnJx/omteiaLurQRg6Rhl1kqaImeCchjqa5okebbDI012VgP
e9WrCkodOzW6UI1ZGKTGs8Rc5lmYUrrSUGgVJc+SoO10tFTPsY8Ul5v4AeV4WvjP2wBWtJ3YhfmB
UUissham3K/vz65RhIiipPxsD9jedyGCJ8vmmp8gA85xdCB0JOeeKdpUWxn62iiLWhRSMWF1axHE
+LsSPeBLpjV4iRAu/pJQ0WLa5zRAl+EKJFA6iLxW/d9Cthsg1FyxMJveoT7XnIHcZlsern7a/RLQ
vgfzLbkyNJBgaOoImPDaRopQuVqUfLEX8HPU+TDbkeqXMs+QYf7NE4ciwl66zIif1BFoYTNJCl73
jhp4QR7eQkFgYdZ2WhLuEYq/83y94blrlE/qJjVm/c5ticyunNPRBi5lNa8L/JwrrMHLeACYPKQL
7H6QHAZzOVa+qzncS8o6o/kSf94+Gk9NFw/cMFHTSlSTUoTNms7f28AXppAVXI9iQAtw+BZp9p3a
NAh34TCUaJEvSVvEIywPqBHIBKxmgpa2b2IcdyTFAZx+6sxXDa3QU9vvX79VUe3Ii9X0OJmQkBbi
IcnhOp2OuCDK6Q9D/kl0zP/h6cmLDCGt5zM9oszAsXtTUetsxr067mieLnVDH3XpOGuWIftI9WNZ
xASdIX0epIjypBSQNV3nk5Bhqo56kDnULWZ2ky1tMVA0AgPcaj1Vom3koBDHE54t6yMz1XzipPEn
AGDLKMrevSz+B1sAd4QnkXrapPoigQ0UgOcqV/s4qKUpK4aZ/RaZuH2LWC9WjN2ylvJLGzSn/Rbz
tn2NQNtxWTPsuctIiIU5o0foYPdENr+Z0/JW7qWrB1Cm+ipaDlPWZhiyMvk16pd70Nkx0Afe8JKy
BZ1FCEq1+oxH6rDAUARFs4qELrhK5eD9M9yNZ/m2uzRe234vSc4hMiOJKsir8uxLCsgR/YazA85K
Y1Y6KlRzsKCY9CDLJpT4MrK6pREDVAFKsScezZbqzuk7rhwwe8Xg3z6Kuj0Ow/qQebG73muVpyNE
ORHeFXeJW8EQSIVViPkeLc/eGWb1ScUBfGKUMnMmqJ7plT8+ey/ZSk79mh64sBcMS8fuuWn6Jbxz
WQ/sauvKYduLhS0sn0BkbfG986Hy4penJJiF5qPs9hoxerf2CGQUcZzUHPW+qBftGlOMPwoOnMK3
Gi/ajFthYzz0fjXP8lmKc/PehtRvo5iFz5g4wM56tCUMX73QvtUjhFaqKbJzL14rstaxXhsyjsXy
636pWig24UbqjFVmg1WRfPqIyx2jZwBqWEHDEz5jcbmfbuhJGoB6NNxmE2wulf5LNeZazOce5GN1
6+/NZkxLFRGWy6l5hKfYU8RW6c3tQfdECNw8nk1eCLOIjcW/ikiW9ZlJ3AM42/rbLgWI7bj9QJTp
JnWcbGjFkI+qCWRIKPWxcNhP+b/9FJ4AZ7iFfScHr7lLrMSXdcKs+PmWweaJCw3ohSt44eVdM3TO
l+BZYJ+Xz4z0RJFPXFX5NNYg71/3sLPqVSDjT72CbgVhkoOvMwtA4eocTBXJqpgOmFgnj9H9kSoc
yNPVWbTbmIan/m7fdJDXHC2eVwD/OawxgCdQ6LCSTbjXmWHsNsFWpl6ZbIiORDBwtmfCvOFYWGic
NSDplNQ/Q+CBP+Vlozn0ll76uG287AxKVt0KWBwsNXzJeM5KcaK9ACg6RQMtf6k4JCXIytP9m87w
hBi5x4o5LGZAM0TLQSP+JNVa8qe3+xEqAY2GDLMJOKjK/P6Zuy5GV4XMuLw9sQbPu8wWvM/q2360
o4IWKR5NlDLT8BUTAf9siUFf/vMuicykSXvd2tzW40LFNJz1nzVldT0VXIowGttiICUfvL8S9vZO
GnsUVy/xtTqFqhdPZQoK0k7bBIEKLofcqUTOSd14zH9NfShqG7K7qqcfLVfhMRUl/ZjbQe5FZYzK
sRqI1eT5KjFLTdYOLp+mS7331OpHpLp44TYgoVup3rfJ8VSKOBiuEY4RKk+zdD6WzJ87OZ2rxwX5
vpxvjkyFbnLOq6ct6TWBq9K0pEsfqN9sJ/IwHuEijewoUDf6vijC6bYyl1IcwwcclPK+Uxwi0meb
q8UDvuNZVWxfEkMk9MOyVyMYNXE7A3UhDudMrZkfyQdUWT7D3Pb9zI+BnXQ3qmIXWpaCJ8Njm9Ho
febQPAfsZ0fer1msLm4+SfJfg1x0u+N9JAxuolmos71FeevoPvJx1mVsgcw3nF7akf8Ocdbi0qA6
NS6ByplpdWTcjjL6h8hrzG2OMsBUzv32D3pSg2uqmu/G54erimpn9mk5o4JscT8aoGxIbHxgEBwn
Icj8qzhXbLLFCaHLVaeOwspPnNRA1YgjjdfTRSZnbath6EwDggNkNry/Yz8wh/V5oawtSE4cEvoq
8FmJgC/j99JgnuqqCzHkxrZEEArEbbQweuUoJXB24iLN2H/UM/i0lCajEljaeC2fusxkzUXsyrOg
tT8TSKZxsDcMu87ITURDJyL6U2aI770glHsrf6s84BzBQ9JSU472QjGTpUJMJXCrp/NAlN56Q1y0
YbaBEzWYz6NlPaX9e/LI5mALXrO5kxWoq0EUlVSQk5yH1x5zrGgUk26GMX7eTuAvgqR3MhxSeGTq
w8MweUuWDyuO2ohJIzkkwHgMKH1f2hHfXOYZjd0+gJpiNm14YyT2yQRMBbNU5ale5rclIbtj1+xJ
a0lmyqPy8C3iMk9vAOLaGo+uVMI5tIE5XyIlIlOau1a1hg+RfQBIZIzKbI8rg3lTcDCah/ntutd4
uQXvtxqgVRVp41t7zT67PBDp1CoClAmfq3uTUWC57vULYEBm45sYoavgRFwYuKD2RN7LoAl+mUyT
zpx8upzoxePENS7G4cCuamtysJ5FNZ9QTjnUfeIPCv0yk9k8Ib0ZEpg78mMyTSA+8kAX95B6m9Bx
6OSeTUaTTtMy1c6Onje9uQfPuq6lOVDIrub7ZYpxk2t6JMpDkMx0UlpOYYUfpEn94b8s5H2YYfeP
gwgAfGdk2DSfvhiNOxLXN1AO3S/k9/TAj5APekk6cjQXHKFVKRXr1tdwQcIaPGMCbYrOAxMoMAbo
Q6dHwMiSLkRUztAOHlfy2pCl1Qjgb5a2XQ3oqMYAANReiR8fBQqSYmLo88wR/UlrwljijgJI1S5l
Bb3ZRMC2+mEdoCOlcE1A5Cz60ymcLbc/rnLh329mBBms7JAeiNkvY/sAy459VXK+WGmnBr534QK1
Yln12adb15b94E93ofl9J0fpyxu2++0n+Q2MPhDqgY+pCM2BkWf61aAgLPmCCUeUB1Bnq0dmaa0y
eafazT8wRmT14VfKlWb8Sx+taNw9QldoHugclZw+SvnEcn/9Of84tPsM1G7Y7H6oxEHTZlZ8yHPn
00j7XaM/h/ihLXxMMAg6J1/BT+MPtlCKqIIVOtyF6NW/5o9tjX/rsQlVOmRhIemMT08hhLvMH+Ea
cm1ej0CLxJCPratNo/2kOCh6dPJzPt0Duzxv2hkMGkFfEtb9NvhOIK/6fPP3JEY2746o4Lifm9Pw
qyzHJqGwtDTGylRu02L8B2yQZvRQ9OqVM1kuzrBDjwfqgNMl8F8in+o3kW3ts3UdQ4yZbY/Evtk0
hijlmzMx5oscyjtiIB/uNGRo1kohcnt68Itz/61Tx/m4RUlRsFgs9oEUuvWLm5yObaWBWDCr9hvt
SQ+TMxkB2u51T4Ga9e9z7EPAFS+EfFB0dqNEFDvyIBaJTSPdiC6qmquAvr5T96Rl0yJpQCoh3NDx
Wz9ekYT0sUuU4l57yzbDbrDrGb3F1xlNz+jWZfdJdp5NJ9/wEsSAT0/PE/UNIZH/zsIrbFWM6Fi6
LgVkvY1gCM7qmAUdPVi47/NYyehbZZFw/HUz/AywMRN8oNgd5RELNXVLzeTG3xdu9YLU/cgCd0bb
7xz0izweQq+AXqb1ZztGDgo9nXU6vrPjHi6JqDAot/sAiiRbDx7NvIQm5QcvjPVWDXw4TSpp80Ky
krVEk6gfDzX5Psx4mpIwDtjAs2eIkSDuYmLRpJN/2oWZnW1ROlLJiWCtvHEbMmwfEz9j+Y+KON0E
1UnFRZQP3Vb5/bmFatJSqD2kAeUYycW1zR0Tw2+AJfA4czuKD6SwcH+NSWe1xbRummg/YXcNIzi3
6ROFnGjFARo2nE4cXqGYNskP/tqskleSn64XOcLxIzFjdcd8xaPbUZGJHx7X2b0+ZjISBsSW1W44
zXr75x7U4cuYIxuoEDJl5d/2M6Y6ePPZxIIbuxMZx6C/QvYKuH8AAixsuyQx8/dlxRJ00jgYLAcB
sJyGASpBKws51Kr4CvCWMBVzsFrqg0TxwhJPhGTJfHc1Fu55tPOQ8D+3ZAhuh+/qDHFS/Bu/i950
DNa28XAeBGyCCSULxiZky1dyE8nOsMk/i842/cjC4iSNvjf8w3wvj7RlX0Q2yppC3z2TYEHRZQPZ
XIEnbNFUdBICsW6xcgjMe66fpg/lyjSFx2gczMQF3+I2x1zMzvA/TjYp+N5GmCt8b7WymWm8B3xr
7BXlO77W9FE3bOvxtcfU5VqdpS/aa6W9Zvz8SiJUBJTZwTGInrNbzyzxhfIy6oWd2rfz+7VU1Fc/
x57Zt/MF/N22IrVZ+3dgqMAX+xgPz+vj0Y8DSbk1mSgs+s0LDJm+dM4uoF7R+4TFP3bvmispEpHt
dzjKdLA86WX8tllHLSo5gcnRSfTPsYwr1QsbVN4oyQjTGKs+c8qUStZPcrYTLAgQuGyHnhwvkuNV
NiCqqaEMux27+AA2cVBardYe6q1vRE60hI72YNbgXdYfWdnmvtWBzB8+c0t4lcKqHiVULCUVlhLM
Phv7e8ZsJ+tvnITC4GNv6ELKjq8hdOUdes4wZDdaZCsVOE8Aj3C7OQNJ0NsGJcpnbBjykxaHMCg3
PN/TSCmeEeHNAvCFaPGYoPh+W6a3e4ucztmVYzZ6ez7qTzTy8pOMOnmelyGSfB6Qu8Mp2MXohzW+
XfIwUdDu8/4K/90ckCBxwATx1g/dzw9et4V6J3lwHMSFmaI/RSR4PjoSMVytMnkHMxeD6DxQmC4W
SqYrGe9NtBYLkP5Defrmr0FD48PHd6yOutZ+RIAYfxbIdYKGn/q/J9oERyES6v2iG0iujNk4xi/P
Ch27eNskKLvpbV9F/8+24UF2iMd+qKpM2eh0Xdii6slcTKnkJPMD8BUBpUbdbqW0+pxdub8H3JMn
z3nweMkkAUb026QIWSPnlY9xqg3TWGe8glVL38Q3BdnwHKqqwZbPCQtChcyjSHwnvLZlGaU20aMM
pFubpS7xDFGOs4BZnDQpiMQixf1UGqDbBUce+6zXPOmRlKiYVhrb6uLaYMCLM0KV9vuTBC8v/Nob
qP2xkzujjrYuHuoU717ATYlxPUDS7SfoCBshwnBr9ox2ehQebavVwKoB4vA9HMay5cYivwwG3V1J
y/T8ZjVeM/NL0CtvKa90fESAqP9MKL/1XJ9JWQ3lcLM0HDoV+rcSc0iMAXqkY+nxdAeHb/8z9Cd6
Hg+Ln2pVhcq8x+po3kh8CehoF2uRUO6/yQOeclmZACh0BZMuMcQXhFifBZCDHAOVo/aeS52Z+keN
ENmrEAsenAG9mYn1TMphg6gBXCwbMgI+bxlCvOys/DA6zPxJ9rExPYACccuS/W5SUnAFnRL6xrt0
NQ2yNrMGOxOkWqo0WyJOQ8QTX2HwfVJ45RG1xmCtF99lKGZfbSjaFyqYyWfdEw5CGjggu5x5nPTQ
BCNdP4WZnz12r/N0n2crOCXPsSTySxB9A5MN0K0IRnMB5aoIpfm95Bse2+xZDp1hinNsA1Ikt9r6
0b8t8K8X5ARVywDIuqgR4Hj6RgR0UHBwnT+esqKc4pOmXP675Y3a7540im+VzWFzx02nDmvqVSyQ
G4RPQY3WAGRNiFlXvVSOSYAb9QyO72pt3sWVleIv3csObFcHMVxrEUyswAVsuKEj1RA1zAF9NSrX
cSz99Ws4XPsSqcsf/YRLd/dvLbNR6Lll09457X0tdFotH3ArJXMk33gE14eCzaCz69subhaO8dZP
0zfrcI6bYwde+PbMY7r1AS70HUdIlmx4jaPs3tyDh/dCQcYjwtaCxgLO8wDtOMv6+L1IYgp8VdqB
XSYXXQSJjVYheasR2T80hUIh8NY4lg3qCEiAqxuDN26mJO0NrrLYMQ5g+rmJxtfxSv5hHlVNKPze
uhnmOKwqEsKR/+fO9/AHj+VEf54EVlzasayoLRY6uExRZshm1t5CeeJltTfWfXFmtjQTw8Vt3Huy
VnNrGLKfaHu4BWbEVS3aMXSk9h/iNFokyPbrUmD4cpXv94wFD84pi5AfMzH2FFZYAEPzLhhMf/5Q
ZwNthTbnwf36GkEVlYls+UMOb/KYCyYtCZbBuXiZePqrv2SF9AkLOWBPCSxjYQMrDu6QeL5iizPu
MyeHO4z/rr+JIIrrZiUoQYcfWc2Zrezp1MHS3RXBHsvip2dMyJOSx7wqc+Qe/WPL0ARHQXWUzBBh
a9e+NYtrQV/+7RmZyZaaSJKkSaRuaWyUboU/9NfRhSS/E9GXpVBldoJi3imIYRnw4Rnyd8wMiUkA
RUeKIDMz5QasdWDEYdvBfww7wG4IjA3wLuJ2aaMcWRmGhuoyHZMy3FHJaxNr1ya29o2ZKmvfm8C8
lrAWeb8WIxjZEXhWu9bjdIt0Pe7tKds2MdJ9CJi8iavhElJM7kHgJF6wSCQMShvWg6L8hpXrmdVr
qZ5zz+Ve1F/D68vLXRxjcKX56bBYOTPDcpWZTewv7gWFmbmkZHdFbwplDu66VH1NHtOIl+tLTeyY
NVF8eWdIFUlGkoiH5Da0zTFM/hn+zu7ijaWReIR5OzBg6vp7B1XbOzSlQ8lLaUSncqEWoJUjF1XT
YnykALjqIMYKUWG1WKro27koXZVAeSkc1HXFW3b/1Hd3K2XYi5NGLM6Sj+hLSysvIbEd4k4hCNw+
p1dQmoPH1U/HoR08vG0ovX5/SCD9H9ZojWCLJB2+IgTT54Bd1fYAFnTsr3484366gabjqRHFS0si
Ws3YiWlUUI2EIZUR3FTZiRyrkn0bIDknZy9nivjOpP9yKTK3MFxkSQZwTPWK6BGvu0Opu6y+C1pk
LkqKCX5m+OkP7J54go23Jv+jbFavWwOTE6PKMO13Pd3TaBlLuznYOcv+UZxtzVqda4vJ2EuLaGFl
TKnJ43hNJJiWWDinj489F/oRrs5wzKwkMnTbPwf9XZiP8bQz4gQF8ohA7hOzhENr0tRf2DMjeUeE
eYo/EBTxd5YWuh+MV2QE/eWu3C8FWf8PMX9XFd6ceuBoVfmRfRHIUxJGxYiqk/OCHgW5p7vm1MiP
YwCVkvpjugfd/l0+ZBCLHAlxdyqq60mN8jf8dyT3zAqzxYhLbfekmUVOzXecGCIENjLnZAOymQ5h
wOd8cgoYIslcp1qPacMD5IOLr6BdVEv/J/x0HWo/kBZ9QQETbNBnPpgcrE3Ll4wx8C3cUZmuVs7V
eKTbFMMogQKqAJSVGO5QcQgf6BNlFaEeJPYidpGbocZtrWKTEUOT9okeVeqnWh9A1vK3ecgY15nV
zUN0IP3Te+E1Vfc1ifnhL/IklCKLJVkpPOk9rRXutWgWJhlrsqpW2dyZhDH2KPTfD5Cu+DMgP9xH
YVoXjQtBav5mjruhuu0wxPiIDkRCbPOpMhbrh9OqUv0DmRBvOx8335mdyYNCjk9dsqFD3shi9CNw
wJ7MxeLy9/UlXTz6PdPK2gKvE7+3KSCSSAxvJ/2nVeQ47V9rVV9zbSIY5L2qwm2E1zs2bIkwkUq5
m4Exdm2tFrcNdWN+Y4h08DmlMhOsSuczDW9YKgnLYUGWDBzueNBWQ+gKtzoyP+A70t0nrzNxdrIM
1W97sRYDCt58TLfhrXKHw5NFWKu8IlRSx92AkpnyySCeZvnkBrxnOuCQ8OfjMoErR7lMUeuc/gs0
Ffebxuai/H2G+iDt64IiS+p5F2HemoG7DBmXf4D5vzwW15k/6jhWSw6dzjwbjAfSE9+NcJg03dh7
jtEZOU0pKWW4I6t1yF8I2md+PQz9qFnG44k2dhgZ24xWczO9fSlj3visQJO8hCLwatZJTYY901P3
AprxVraUIfLBoNeyRhp0RA0g4Kgqo/6ePzAdQxi/PG0G427EOd2mJSwmWKhtCpIAAl6WSkj8Z+Qy
5NI3iR8S3/Qg6S8la3oe3AbUGYXPYYYtjR6ghUMffZyHYk7DFAH2CqZZuYkCF7pr96jI/S3KMQtD
o3vqtVPTf7VjEhMNY26l5WHPyKJls7IfJJH2euHV0CbSOm0gN9ScmRlqWiwT0miV3V8f8TUVvlvW
V+d3fAIoAjzoZdtKy9WrIOu/FfFV63Cj9Pde1ymy6ddUCQjyIU8Ldwnf5ORsnUS/doKkRakEtIlw
AcaOu32C9KOEETTdETLsXcIxy4jurdO/1OQs4axcN8Dcf7lHSWmT1gfRP7EvXlQERgF8VD+wtfrM
JJGAPTU2E6v2TXPFr2DEf41A5/mCq50Y75xvESJIos4HiXeGR01XvXI33rVCEVWSANlpsYFOjb3W
0j8fPcylZORkZV3w1BOgaJqgy5RPhTJK2pjrZDIVLU+OvIEj6qnLqyh+7XCKmewnc+tllBUxTptY
QlJ2DnvBdjm6MbC1UONCjfN3/6pvWUVLENXMctaN4Fhz/Ea5xGkbBIFzX89+8MnyTl7eSx9ZPSvc
OEMcZW9Y6Qpae4G6eognq2uU9p3/u4oEVZuO/vi0R2vBf1u0TY4FdlFAlqjnXsT1xka+Ega1NBtK
zVly8vEmGgarehWJ6pWgP/XBfS946efxHj1tuRXih3Q4JtSikIsaB2E0QHq6eGdFbzjF78uVnImu
0co+sUckat2cy26NpgEIYVx39H73Tj/myAu62XIP2HkqlDvQvHr1sp8y+fB1d1AFNkpllTmoJv3r
zCJAIe7QfHqQ8dANdHrPwk1EdjLDyabKinu2MyEbizyCoBaLtKCGgqyptc0d4PaIx4zXFDTsqWYc
9udZpi/HMXnmJD2RDsyaZzPuGcrmlm6EmgjlT2VKv636f+P1/MEGYK1dxkzT8VwcE9WHcsJGas+4
1x2/7wrLss0iyxzZY7R/2UjJtnajFnmAtzsIs8An4N+A6+6eIDE97Pao0i3UbnWpZ75guZe0OOmD
eT931HRpbltJpWoPGS6WsuJZ65NHT1NiEgc198wcZ69gjerhj38xYmVq+FUnK8t1YYsJQ9JkDdPg
citS1DmFK/qjJ3KQpPsaaiOcqD5XHOfb/XpiZsaOx+8xUQCBE2ID8Ck88Vg5DvVQI0LiYwr0986p
b+nq2W/nQJR2O8dX/MczPzmq6TYT4suurkVYtdQdBIbIdwmE8vF0fDpY5oBYxtmIedblzmzo8s4L
37DrYwVXBtZZxzTkItkmS/EZ6KmkeG0GfIdTEtX6VYAY/7JOCSldiEo+2pctHsmipZgjxcd3sl70
8E58YlQ0vs4KBFsI//uwHH8TP5R98rg5kcXTieAFBMjUnVhvFVhtRgGpcDZwwCFY3U7t89b+dBki
aEkGtlHjah2Vs5iHhgHTMNEp5G1pJRdn2JB78frkR7xyJwoCBdvCL9TZIUGgqauKw0pc0pWWRTMp
JZiGLq8MeZa1xssZKxvBOTQZPuNtz4yN1p/o7JInodQmhwZMeJJ/R1TVcQfudXy1HDyO3fgfsJyl
g0e6Kj4DZqNI2+elLe0VCxpnF5R6s1X5tV4ZK+yb4ez+O04TUOCnP1mKZ+c9OhZuyrrFoRwJxxeP
aRZZa/g0uWALQrfLUabJKox18mCiP52La7We6uZJgn9X/TNPFypw1CT9Zdhb1P0x56jm38b22S8a
IiYmcOPSfo51urvQ/pYB664ZxqjuxlZKd0gThNiT4uM3KpyU0h6YQf6dNdbXI9hUzGP5MzxVDvFG
LZaOecdi2p0GG65vpE1BNL+mbYY/KGl1uz4Vhz7aUNZPtHY4qf17B4D7ZbjrAHfRZNJ3lLMiVP7y
x8LEFXczBVIB1RYTgcrnuXrI78dj2E/V67lbxQ75KELoGHxVP4qr5W1UlfBXR/Wj6FZuvTEtkEVa
zr+uO0gj+FvussWz9WEl+XlbldzyqriMHRYbVMOvxOUeHTQU/HjWmgArxmBTP5mzQUUXsIxLIWq+
5XiDO20IRK6fkbQLX/dm+poy/DQp+zFcMyucc8ebHsfIfBkkfzFs4nA3T2Q/MDiUkR5L3HfqqhvO
9WVeKYRu1r0d87qtg9/AHKH96vfnqXLbb43WDyIKxFORm2jb8yqkrSG/5qKOgTyfRKyA4CU6OC1o
iDW4uPQphAFnfJ1wNI1E5JcY/i+JgrrCB40a1gB7HMr07lydbi5QZRJ5V1KxZgtiaARGCP1mb1fk
NX7ZJraPuzQviOfMobcEBwOFzW2lrZeXMkQjJTYiXvLjQ2/9eVVq6a1QuV4yh/+vqaPgo1hX747N
S1np0psKm0pph5QTi5qgvmUie9wMaV80HiVYpGRLNNst/p5e/VqZ4g0h2JjMPiBt3SQP/TyCgU3L
DOc7h8NQdL3DVs7Whk8JVXyQS3JyG1GGYmpxrnt8SECcsreaDUddW07Q2keIe+W2qZP2/1N8mcxR
Gre8uIA4BTuspCrsm15wHUZ8l0rkOcUvG05IbQAveu67FEOtlqaF4YOrpuCUChuBKpbTsISBigyu
hbyUOlGLwpnADkzyUGWTa4kTsyKtg5zn9sItJG4S9eaykwhkKRCSgPysPznLRrLm1XQP+GJEC0oe
SuQbdvjdOLmz3xW03AFT5XGm7we5AhHbkFkLwBTOhp4Q4d0NLqf0z65ur6Au7dSVzfX+k9Fu8I9A
6jBxW6hEiOQcmSz6z5555h1AO8aS1XrFeogkyfdkZlCP79bF2yT+0b0bzX87cELIcrlfQAztrlkS
5bjDfC/blOSQGXdXSEeg1rfJ2IvaF3rQrn71XKD+UW3AJWi75zdosxC/vIE+ys0D2J92VgFyCAwW
+z27KjnWUNTN/PwhT6zrb7XA17CmDk45Rl1xnBLFy3HGcf/xE4scy//wBxUihb7Aa2fO3d2iPfiw
cI4sXpEukJhaL/qW5YAHDopmfrU8J+KWDCkyFO6NowOHNU+F3S6l8cA5VDg005bkLo6OiPqilsqw
/9hZ0XyArBzkMOaJYNgl1JDxUvLdSwFNGUt7/nEf/DnJZWv5ap2cz9OcbMeszPqVb90vIrhQapQA
SXoxn9LBBs/EDTQccpTTe1EEEyM3BMhvoZRd6pxI+jIk4zmGVd2H8vHXdK563s0/874PtJLLc2oD
CFpYReGoUJLnQfamKp4vgyhud1nbFdixRi8++GbpHMMbh1MU01EOQNUEYtmgj0p1X0by6livULwG
6U7Qv21Q2+LWAVKkVnzgLKAlQThiGVUqI9ExZgkY5tex6WwiqE6vHxFaSB68nUN6r90ReaVHPTQg
CUfhGi29A98nHDikH4tLVkBtwTH0NUAGEEA75MFseJYnijB83MoLLHFKD8NGZhuWhn8VbBgKxgUK
a/FFDnNCXRRfXEuW+nRN2y8wEdkNXCLx4kSR5+evKgZqeHRWjqxZuvz2O4PazZqwSPK068waSjAm
nV8Oi3YeRd+rCRMfc0PHIQw15puV219TgH1DkRFxtLdstgp9XW9X1GYYq3n40k1WO1J5D62uKyzh
IixUz259ypcb+druXK/DVo+MiPMNDM4586OmDtLxDhR/kE3VE2ZprUlc0OoMWHYg4XVHfY9eeJxW
EoKx+XLeJSGv4e2zu+FPXnUVP9pFnZ2HdbO8f3OzcbOrs3I4vyuiQWcPyVQRj32D+0Xz7WVkMFfI
gIcROdbeKHcJB9ITKnCxIK36bWSSv6hQ2j8Q3Z3a2lh127fhSkXghlta6LJQjaQaCDHKRz5d/mVD
avgMsBkFujvrYbV4gF8wQEeRMfIpf4tkEuspBdK8nzucWzaxJXOaPxD/M1t0O5jD0hSifpWAF3+K
CtL0hvm5V9qjDFDI7iWKWjCEnGDdqvz7v62yxTr7PNxe0nX+BiPX6XK1PePKVF0LdJcE/JIaUlYR
s/JN6hvS4EMPNGVF6BruUr3p8v/bZ8GqSF0BuSCKp4Eu+RonIYI7+gMzPBnV5HRExRf0U1Ds6asv
/ET3szaObv47AmoWabK3kLRuM1EY5CWND5JoJeKiIzw+8p7YP9f4x3Qqmt45Zvr9CgfBr3DXOips
BLmA11sa0UjfqOojYkviAjIEBts/GLnt9w7TFwkZn7dDOm4pSrjEgihuEFfcW35g85WOkQIymE3H
5Eix4gmnb2Z+0QUydEdB2KRD0B8OMY07cpxUYSdU2K6IwkBbgcSLyDypHFC4bxVWqu3id3vcrcCV
k+MNtcE5DqJDOAGZ+za7iEbuvchpgTZde+qKwqXgEFS8UwtU/mb4u69eVkKZW6zXA8z6FhdNQQkL
c5octf218RMhqI440CxE+ywgc52S5frO4FC5L2ImS4GMtxlrxe0OMJxqsnLj6HsvI3Pl44DXvEwW
G7L+Vj1NuE6cwTa6oZRy5JLJdaKUtkvvIfPV1ep69SYO5f7peIESTpTGGIERylj3GMaiu+bGuWlL
WcJ7uQtUx/LMyzHV1sCBdmbcdnsPw3/fmtD+4guWG4v+YzHEY0+145F48eNZw3D2rViCZ1c9mkEU
X9PPVzUpNXjl6maaUfhktLd+BoDvknVFWSviT/5S28oOMVbVAKoRzHSmlrhM96j23/VTN0XUxf5X
AMmthFXltHTC3VUp2n044rsxA8ciaZ/WfgVHOBWXn2bRV4meMLNPho8J3kZZPtytH7IwLrAAKlQp
dbrn6YDhW4oCHICS8zB1Yeu6suF9xQ7F0k9KixT4RFhw+Xj5eoS5Xt1QYX6TaJQzXBPYiqfcsT9Z
qTcrwk4FuHgNdBAgQM6k7aN38Axk3BrAgu3doQLZlAp7z80ezDkiZbOv1jiRViv877NS/5Od72bc
kRnXVFHPry6/b0EVcGHD02DEJPP1YUJ7l8nla8vPA2AxRRyC6Un299+4VnOz0zEtgeYrv9WnLg+T
SoPGHPaG/eIuepp/1v33ZEQEipmpJsvAzs7MYBa99VC/jt8EaN4i0HYnZNcXN/weuTp0+g8u7WeX
xDyMiJVI6YlyeL4/3d1G1zBHE6FhfPopoOEiApTgVvYxExcALb8Bvrozm0k9hzJS4XZHu/mCYVOC
tjv2DGLlP+0y/clHgwGbZ7xLq1FPkcxdtd0moVNEQXM8VUFxH6wx22MFGF8+P4uNzx/kSNOR8xmG
a6xsWAnGp2+Rf9lWtmCgbLSWPo8W1+FXC5TqfBmd/IZOQTV8IdHCvl//kcnHhVgu7Lx2VIhpCz3P
bAKWS4E8JvCqE/S94lN3CTG/kNqt882lL/6+pMPeJ/DdXASHHkldMs7lnyyloJglG8nYNeJcL0PS
hb7u+ep9bOOsz9y8ec3sPiLaX0LqljT7w+DerL7C1soBWGIsmSvSGFeVVd94gmftnLJnZRbceGWo
dZmLGWTDll+sGBDeVPgS52/ldOjrzogzXRGn36oWXAtUlOMbgD7Jtp+Bm7/VgpZQkrTJhf1kiPvk
IN3PeZpn0FJHQ/i8sDP9xIxW3DBntKFr5wwSb9XF8xtlx6gmNuV3qKMELiEaD1hEJahNNxxdqbDz
htmrV8g3yMSdrVMbnSqtebxZB59yqUBnXoBhDywVbQz7RposuDaPRiTfclicYhLh5oIufEaCd6G5
4VQ60q2LcTQnSbUbyXGgASGiB5/3qyjLttLv7IXqODAcbs04fK5zLYEw8xxsck5YZd56igUdJxOl
7ls1ak4WWFakCJoUn7zKyufV3aYpwNks7vReJxdzQMn32z9Sj6zeGMYYUfiE6QRCvqiUcQjFTDbl
j8EnHbXJft11WJ9EvHaA2K5Ta2gYbNlTQAP8NGyaqdKzIEIymXOGdtfaMa/IwMLGpxPvX6Vz92GY
U7dvUWZu7JiSqqaK0mtPEE9HeXT2jeimx5PdLF73UlDKp8hXmakoyzRVt864gcnE9Y633xbB/SL6
J6J8R4M0NEMbZfqzEqw1QCVlJxt6kP1Pmq//9H1711FIpf0jZKGYdkPoUWHslc/ANiHL0z27QH0x
qqs6e70tPke4cOOBpbeoI0tmAC8TcvvX8QyEIffK14Gj+zCyU/U7peoZkS0+0sVYyakjSJiy9Erp
KhCW7WUnobSgH67JM89Vb++npfBKzGgWyL+n81v1XxL1xphgsCgXtlKvQax3Ma4d0OmuFwel4jzu
qBTq2Q5VaKcxteFV2saUD59Y/Ig4rnxcuxZzBoEE9dmhR7M478y0WRVzrxFfjBJE+E++0CSGtqdq
2p7gnj+SGX6qOGm7mYSX0H20WGzE9Rm8FvtAhSCIM8Y8Fy6j3VYnvQfjAbipg/pPOdAEBKBYtii7
WtdhWfT7Ekzgyax7AKB5mcUUpQIcD9fKDR74DYtrEVsSIkT6u5jqGXpT3JG7RXPLYMXvP5rl9Dbu
HbGw0pNoVJ5YHKYk5aVoZRJkNMA3UJxgcal+/cyObZG10UlwbkamEqHmGo7YwN9bvK2wLSrk5vOf
nC8bCNm0G8qJKpdZGzbLenuFIZ8QL5AwJTS4+WY2huCcvnLgdplgPquOgv4AM87a6kYo4roavOjW
UrPi+z0kWXgX8EYrUeDkbA0w1/0OZQmG3xs4WxELJA4T2bvp4SSPjLOO41GEaowkiKH8LR5r0V99
9lH+aiWKOuYW9wdDOSVCdApmTWF4i3cUbIjW2VwCdp6uyJ7Xs4HFpafCPnqjEa56spoifMlEbUEG
GxnuCss587DylLPybFlTbTrciZPUbQGAw4c5FrTj60tJNKvNEr3g42HkOkt+puIW8GP298+Pmdgp
Hmos7LW61W9rDmesp8wzhPPc4crWL1Rn9cQK0cNogM3ngGowhaw4tywLq8zraDmdmapbd1AyUxg/
fDgLrGbAxN+FGERIgh478ERwVrLceLlUW+Pedruhf2UQphAxV4fuj9N8Mzq3Yeooo1zOWMmRgNTy
RpQZn39douoVNdZQFRaUL8FiJ/j4dnmxSs4NcnNokbQDJY6T+S9epAyviuDEUFqrgLxmBpX6iho5
9jvTkTZp3n4IfiSpmpNihtWjP3cqKQnblMcS26I+5BiJdg5V8VQbD4nCIVxAj4r5Rbkmv4J7F1J5
POxbrh3Uq0Ejv1ex1tPcqRDjwgikuLDJ5x08yTQLWkrNi/UODrkDqLC9D3g72Y6n2G6/3BPHxxb+
CbGwr9okMa7wLU2U54vj+lNzdmowhcXd98ALePysTD+yaxxJ27RanGAxsfNqRPh5cfd+Mbfv1c0E
HkDe6KwmzZRSLz5hR3WpBP7/f1RimQC8hSugLODYlFLV4uEy9THYx9xsM+VOsQpwwb12NEJXqzOl
nGaR6JhTWD/5Q4bg0Oha6bkorv7vX55BAEdpk9EHS0Yg6O1PSGpOo8DDLiFXZ8nmVM4dhHHHSF+K
mVixKKaXiLMsgLl9ki+j0Fhl2BAzG386EYYm06KdSP2Qd47b0L6rJly/u5ShaB5ck5/gjdPlmWxO
480AYcWl0oVRvHBTrqh6s3bb8G3LpRiG+ez4KwyTCQAvP2Ee0DRDGTFS03EpRhg+2PZNLFSlT0nD
6FamhTISctGnveo4l21+DuRbMuA/v9NdtGzYkyFB0cl4UahyBPcjodOhGqrzjnAfsyh6HQppv+mx
bzR2rIhozULzQhmggrNjWeAPsDGeYUikLxCCZT+MTUZ5qtqubnmfL7TtMqICOwC4pTw+jOog0n1S
1cjLQtkynVmMhwd4XIx1LjcMS5+F+/DVUjGEpbmU55/6xIu27JGoww5ZRUueIi6SOfFddOssF3cM
AxE+BhQDTEMcRwjbYatZa2eWHGCdDnCtzGkYuXGyv5BDc85KrY6xvhdXF9b38nC9QLyg9q9+edcZ
wLEUZxWYgkkzcVyQ5KSLKEC39ShzVkk6YbooLkacvAfXlm3B7niyGnlz1yX3wTBIHNmqHDQvSQKZ
2c8sVcTlNrdujBMQWKnBX2uAgtpiCZeGDzX1/NBL06qy/sRYC9IxQinelWbneo5tT9gAl8jDMMNE
6UAV8qNqzzU+3AxQq21bh9qX8zKOLO/2rGNnLxPyCqZ2nvmaqXoLK3L6T12x2lZIIoD3KK0XISd5
i3Ff3dQgOIkvWcNNJvu44Ky0+scluQTyELP0RQxWLfo5HAqYPNcIbCenSfO/DtcjHkTjd+Ya3tej
pI5qJirnuZTYZbKwBwttIfrZ9BY+C1b27BgqJJYci1zWDKy+8oxgdHKLJuULVmOds9SZNBAL9rTx
ZHIsFOFPgitVM/X5Y5Bj79JCnT7mdmwnNduepauUdoWB0PM2Cqy0tqYS7LCb6SRH/fQlBWGTn4Og
S6H0aFpmTXGxAV4XB2IBJioiElM32dQHu8G/bpXgOkRMh+GgEUfHKwJAsRlXxrE542PzHXO4k16n
Cb0qY10wYofhgoTGis5KmgewYTWOjI2AAXvWwRaqh/yaSpVvk6Ra69jIarXU7/BpuSebEKGYUAvp
yj3TF2PVDE2mURxzeIvuk95FelYs9xeyM6r/hoQtOxKl5Z46Z5F0xjRd5dTAvJMaf/N+p0zKq9BU
XSK0JWpUkutOsVkMZE1m+ys7om7UsUNGlQa1pk0pqhkF7hY13uGICpzz7bL74B43TCvFd1g3maNC
BG/BlorVXPymXSI3Qjf+9D2RLQJgiGruyVJn4UMamAiX99Jl/hJtlQx7IHhr1Zbf//0gCR5ychcf
9VaJaQaqi0a5Id1E9+cL0BYfeK24RzjJ6ByFCnBqBs8OPj8bXtOtO5xLUxZoqlY4fvcEtdY+UKC6
jMH21H3kfEnAJ8zncse/IuKGl+NTWxNjywy9nz/wn1DLHISfuKED+nHjT+muec+4N9gwhWIVWcTh
G0VfPSDrI4PYhVLSxmhTFJfI+8R+Mxr5X8/3jqBcuGCM4NJB1hA5C0LdS6bFAjwQ3cQXMHl3OOxx
OjL5Vpd5R2EYwHw0wTlwyMXJGLa9100HNNHW40pf0AuHagJOLM75fz4fSQ0iJc8byoozBDHNezC8
sNWw9ZFx3fnYnFLctLpK5suwKcT0Y4QQhpMuAvDZYJBWKHDavosDzduKwIl+hyaVitxQmz26eU+9
ccx/UXpkHNxpFyMYz+O6XeSaLvJawvXqesEz3+ATm+bWDOxRno+4CN7yOr3ejpvGwMNLItMbYaNP
UtiE4jTCWlGRu42gYH+99Dp3/2gWSg46sE0viRzUuYjsXaPJE4z4tyifpb4CUsXpFnPqMcCMMDTQ
FoPuM6T7vp+epz1SY2MY3N61fl1i6yG6Krn/0OOBzqfPx1RbyCFk9AbnRbmC2ah8LT+jHq0zOU68
YuFJsg4ktR7cZbALSaCXChhYxSi8iyjeDWb1T/O6FmFLAkTWhWVTX8SW2P4mcnbqo7oCswpfDvcb
gi4iG69v3Tmxe61yZzZGuiWfogOnPMvOoL7ng7KC2M1mRl0esRsg0whOQgaLlZhr7Y8cdOBVWiFu
FfuW2pWvcUYZBuKZbNv4BsLSMRbuLLtLKSrFMn/4pFjfTvyTGFr2Tksu18qI0n6qHL2PdOWm9pzr
xnWRU19EmS1g22iyLjkBH13Bf1SBLERJzHNP8uSDGsh5dwNZ0xZPFGQFA0zn03jqRH/kkbNOJ83c
lmNXFPbg1mGnRuNqjoaDSKy1BJZmvJiApg9sOXMxWAXmHjY/RjkRMvVIt3zKFHUBRkrGKp+4f+B+
AD2r2dfiK7W93Mc1dT8ZSH4t5xOyU5SRKRp8EPKr4V68CuHPghr19K7u07Qo5jpqg1ZYUCGxCRHs
vcWwctAGupubFQK890cC7eX6VnlNKpPUx73eD+QxG4Z1SdHOrpV7sAmXtnu2sxyL50YHzEL2L7KK
8DVixXwDN7oJv/5zyYpL6vsO4vNAtx41Y5r4gdAFVQmhIsj626xJ7A4pYpI9Ip5FIeD1QtFT+sAr
G2xP/HSko7++2J06mENKRZbOKseILNQL4GJe9Ki0Re3VO92oPZVT00r80THD5yONT9XOTz4Bp9gT
YaHtgJ3WpJwmHWnWvkvTCrjU46rJ/3M8gWpTLjyenObLLW5q/FFYYfY4dADow0DAMpbqD8LoSCUK
KT5V/EuL/0AuEMuqPOLbHnJ61yByh9pHcyMsF7HkHLMBalY2JBA+ksLWEhzfqmX8PLrDf7lzOa4C
5x0D2jI2o14+DlbMPcDRmLfOyTVIAAga2qCENXDDeCHDmjbsU3C3d99dliZ4OKYneUs/s7U0cmmI
amyCT3u+dqjODbj/WPGwha6d70NULHQjgwY2Atjgx9lMvbQaZCkQUIHL0ehp1PfXKlVMrqcihLt0
R8W2ekGRYcN+vJrJ8dg8sQlgdDhEdFHU8SH0t2JhDbatUCIEiRTiJ8Xu/8s5mzo6ebzaKL/g44bq
dwg19VzFZEAob9xaRMf6EL5FMvArl+CpCIAUDX1yvDQhgMXOQaDKnD+TKK/syJW/YPrbrIHdXI+6
sX471Ax0r3mvllYdmYPAT23oEHMvK0tKR2HZhysO9OexIyCxr3+iPPhJvo/cvlag2tAxKBuHE9XR
YkL/o6ZMxZl9/PKyenHIvDBjjyFya41JgHFZ3trBar1tniN2MwR3x5VPQiGPzPPSV+fzaIY+AWyM
9+aBd5QXDQmbG5pLG0s9utX4vZWlzgxgtxBLms+mY0+6/KqkPRA6/aiGaoHypLX81zpfJspc+gtJ
9ZDt5R1ZRgnbHDMAY93l1/f2OC53SUSSs/rehQ3MXYJArXoO6qr5zaSbAb/obvbADVty3Eprjnqz
I/hEmUQkDR7ibprOcXNi3Gtdnsjo1OgEsvtIuEmFoL6DlS1adYZfRNWUnPDyDp3YtodDzbj+1xFt
4UI4fE/SxdaYCQTFJqdXfjxecGvJxI6BdMSJ9mnFxoP841ELIlgbIZUIe4fr5xOyzPFgQgdFpVv7
WW6OXjdXI06AArPnrvHCwi8JZR1IfB/WrE3u6Twr1aWIa57VJ7kv9k5J2d0/08RLQXHBaFQzBiks
4Kp6sIm6DqWlJrhMjTm0WLNsyL5YaK8duYlXkhtPH3/OoWFqPEodAGnImLbKHIZPFyiS6sFhsfiI
uEBrmDlf04wNMHU37y/A3UBk4w1l1ClIVvLqwC9oA0pUvb8fCLTA5pVRUQi+RM0yZ79+LArw0AD0
NtmfIxtVRVyqqVeGgi1vJdVoRHFQO3qYg0AFszEfu6mpVjauhhMXz8lf6W4kRnpFBPRFBIVe63VD
N0wKRHHIEGeKFfOYYCyVnfvNYNjQz9qJDxpRQEZspG1DkyIvfAO9t8jenJdA+KOMOlYkQpFX48Tn
OTuClR9/EHs8eyOQOms0Bbdhg6GPR6lvAhu68Ud+FeqN0PKjLndViNgH4GENuqvYmf1UpisvwOhv
GzV1UrDc+z45yXsyUfi652zm1QaIWA2bMl4B9k9xR0aj5AEnJk2z4AApD559G+JGCTJDdd/3KkQk
BVG2xo76kUZgHSHHm9AEsHwNTJ9ev6rez6hfTkzeobM7/88/qO4o0OCgAumloNqwwDqhtUnXNHs3
ghA2Nxf0aTtj3TjkX2M94/zjyzoX0SRKFLg/68MqV0o+fpKAzqcmQwcgTnMtPHo9SyCRjZBC/eGr
t6RDnmjznFnERBYIkPYmrUc2qFIw0LbTOvB+Q7O/y8OBmyGF1J3QkTbXIzEDf82L0CWEqY68N3a1
dgFbvVfmKGJEbKJg4GFoeaKAJNvDE8a/ItEaDGxhm7R1G3ThZMUqGgBwOMkCz8lJizxPigx8L6p8
Bi5B2vUNpIqgf3Wyz+E7lka0bqduDTsrahxlrsyz825kyVf5ZhHlPYHU9n3X2hw+KtRRhWzAtFTl
npFI/SHqRzKAPShkURG8Yg1nSG3DhF3RNXtsATy4ubyr9QbZWaIoaRxmXScYDVagzKZcPv3KVela
wR9RtLRLhaH+OgjbuJw5/Vr0S01H2v5VTeTZ562nXtk1R7swYoazJMacYZ2+Tk0T7rg5PTy+NJ//
i2NTxMomxM6WwabbSBiPmEAlP3heeJV5+XM0m0v0D+ojiBnhFsnhzTEY1kL8X1oxVCpCBy9qH/iO
ZR9Z0C0g26t4IjnjVkVT44EvtZ5Ofvx6XPkbDoG9aBe/Kqz4KcabO6dn1G5ncuvTDrbQMRwgX466
kCoycmWgft5w+aidiIFfZBSgl6Ps3Sx0n6qmHPJ7hFAyE3332Yh2A6nlhU9JODVghO9D8m0jFNGB
nBfmYEQQlUcbxiErJbNmHJEpXTvTGwtRzskYtFSbHj90YQgkYYuKImCt5YtKz12g8S8uet9Yvh9m
jv+UtF9LnNKGPn4toWR6iSSCguk8vKhoXLMK5RQrdR4cL83FvzCwRixDCpFZJkqHSZckYui8l+iZ
PkXGJ91P/2N8j91cbjebfqkpphW/u81oHGPTOoOZ/idyXuIAkjEuGNoIp+0hFEUOrI1i9iWumd91
BgzTsC1K+lDkiiNW4KY3oDMlEaKlJX1GcYlL8iWo+9roi/2jxjRAMchkO6wlIYfrcMU8XUfP3iJe
s4Dvwm0wyf1ElNAwqJOP0jE5IL+qlIiTK6ZlSLP2B6MTOoC8JasQtJvGlfqL9Ml0N53AegSAYFta
R5NxS+VXz6HwrtC3ijC+qp23nDrWsMgy+zpNpViB6e7cy27R9HLGe56EvnRSYaY3DtB6wi/QtpwK
Fu9aoslguq8RlGGewWFeX6SDGFXSpueSb19LEkSJ0nYw/90nfDzRHAcZqmfoWYgzaz1UcBeaRiqR
xSqoji9f6sTuVCxGTs5uPhBpvW1LGOogdlLnpzHdE22rrmALUVhhxwNBaXTNOsvHgL5SBRsW5dX0
eAs4xPN+rSYAnZg2bSW8D1tSpow277JFPuF2D5bAbXFqrhBT3UP9G0KrN+/IO1ioOtZepuSXdkNU
WVgi6mSHJeBGmoWtaTe6sfs1EY1Wp39NgXoZLGXV9kw8r51LjzDCeoLvxQWBBhx3vFFIV8hesvMi
9AEGLAgSP4nA5dGsbvhmZtVuT760dzc5a/1uHohxHcF/COCymjsQZwG2nUFpmaLWEkNv6rFI/2zO
Lt5kfRJkdYdgF2X2T5SLgb49PAKSGVo/18B7SMuBOCcdByZ4CM/REQAYfpbBbBx8qPKojUn01lMs
kckiU25cxcpEh28PQUIaGLxIthQv8E+TqdDU28vgmxLUNgz6dngzVfnKGl7vU0xPvel0s6/EfxDY
UFP2OFMNTfqJg5kKXInqJA1KhAXdkTm2/yITkaSGDAW89ojO80HRtvUlnxPaMOb4pID6Q1cnpP5Z
SqFqyRqL5PSvHpnCbcA2FfMW3x0MntaKNj5AMtKVpiibGwrh1v0671XjjhoxMtBkfAWHWNxDabok
DzmYzxNM9DSJEl0o4rZoutfB8glNOkpNyfG2vYHFcMvA0+uQOPYjNwog+J80GAfwGur5klEdEhyJ
M7NLee3jaI3ig44de9Koz/Cb0rfnsAcI39qmJyktGs/rcvGBGaEtBRa/Tl2G1A7O34LBU4e721A2
DPpzgoGKts58EW32890Hg9DIFowLe/yWj9jWSxBfO4fHAn7slE9h2SUeUd5BgsggqnIKssji7eUq
pEg2LK/poNAVku6Ig9I/ASvrPoYSsIb3NxZDKipOltQK1ODAp3HmBwGq+4Ktz5YMCijgGTK+zh8v
7dqNNlfyH/nyTew5BPz75mmai/qKwT5PwqUTpeWB/dw9O06a9N4nRy1ZixYC1thLhtqHqjJSZS2g
Pwj0JzIM+uqfN2nb6hacb7Zk9NHIzpOaJwJhbLa8NcdQtgdysPmc1uQ5pcr1YEgFFgLRSMJBOvux
hcTRHuyhUPvL6+JVlsI2cO6DzkmiFTUViFVQ5Lk3WKvZNOSqicTqaz/pCzmGpvNyFxK3AL98/z5Q
KfGpN+galwps2dR1CBfxvVKbAverlUqMnvXFSv3JcQibcAy7LZ2tgEfJjVxSHa861Jr6nJpNHKG6
+oSDUPXHDo8AueoTbW1uPy9G03CtDp0jAr0JNslWg1sDK7QLlD+JAqnQqNWDtuBrNJ/aTcbEQYBw
otPQ2YcvJWjnyhVlZp+NWcpkyAnYcErqO/EMDLqJzaeY3FILQRfOYulDw1LrHareUX1ZLJrOx0ZH
JZDUKtJ+mwAZc8KLas9GJ7/5EVjpGcjpMoYfhz8OB7GXsJl67hEE6WxyO79G3OzQy4oVEb6uEdRO
qUtOOZ4AEXZ16qZ16+GDKkk+atl9y4aBfbCTRpROxwwjhxPkueK6sEPiAK9YA+F9VsBAkplZFOAf
v2ijqN+DrzPkMCIk1LaX7Pz+EvNU4uKQaVs2pIPBQzxpVkdGRuUik348OLeco1ZpA5GmV5/jwHRw
dFIttglUjUny6Bvn8SiNCTszbTiBP6iX++lzFY9ibVm4s8dTUg2T4WKUFtY2XpI308qPWDCtLOsN
WOaUid9fB2HUZdJc+LZb/jLVn27e/ecunafw9EMDJZRz3xuout6wZaRXkMARI4KXOxfYfFdp02d7
t/jUT4YGsJN42UFAgQzAaJUAzHnSGbgH1vg3GFF4SPDOWuXBaq246HR1ZfJvWXrpxj+NgfdUDWx+
GyKA35jeMongr9MOcMSnE0c6SW51AJajUquo30djHzca2TRe1KhbqrGNJoIG+EnW8YWSF1l2RlIZ
Y2MSlG3zrynslm3oulXQh834UMug6mpGbXCDZTjWE8VxAcx5qEgVw64oIQ9QbV2ERgbGJCgquio6
laTdN9CgvymBnIFUKy7ph9sXkTM37Q2haoLhvnOxzT800mGELfHTCeB93WCDDjlYpGuzB/O50zHb
9XEGhBTVGdayAvFmejNg0hXR246JkIzu48rC3qN+nCKogbh2uJl6QS9iNr5iLI3zKHkyYLqPSLRL
Jf/sQLlP7wUeinYmRu6WGXcr34s4W8/lrCBmjwXe8oHx+PUOP1RHbNl6BqjIQKlhnl7y+qTrpmQj
50zCIAWCOXdI1W1PXO34pxC3lIquaqa4DTXGenk8CnfiRlRKh5c1tKUBPGJtqcg0cK3m94NscFB9
VzffuhG77WcWfL11Rt45CHC2Zgyj7bVCi+B4emZSyDzXatuQ8fQcJHACjjWZWzO+St9WISeEd1oL
y3cEaBg8q8O9TCnz3GBrQl1h1oDvHj/xc60f56HUQXef0xzT2fTROWh0IIXMkoluOAUbl0UN4pAR
fX0uHCfeNCE+LUp8xEg0rEeS52tf810++EAeEXpRSQWGm5qX4FfW1J5FR2KFuVysfhTsbzjWDPtW
pv38dsYP6gOgegRbhlgqcVgsTgnnUpunv2fPb1T9RayObHKgC4ATyKpkvkCPGqcKRq4ldUjWyNio
eyVZWhf7q5WHmJSaxk0fJ2pL35t5LPY80lrChHMLSPs1nUDQh3fGJDiyJKVLpqXCOdcqF8eG9AIy
EpamlpmPql9WGPUubNgA73wfDw3YT0CwwrbVUn3GbBytO7ugkZxM4EnMvMakl8xFEMYEZ/WPIzl4
2un6RDZz8xpbB6iDdjUePYCajoJ07/i4xsS8RmKVTbXNtZeTgPnWbGZwEV1R3187cgDydPPTZFKR
BPLPyjb6O30k/ovawSfzwkoVjU2s6WRkkE5UeK5KZmj3nY5cscavGPnfueRB7xaG7+mMpWKjcUQI
5l4C6jTlaXrFs8afyGJbrONXI1FZ3CGPATEfDmnxIjUgIACl6Nc0jg/r4zVXAodI7W0i689DJRMR
Diq086hvuKmnBOjoznlUOSzpTblM8z/HiDb+P8PgOGwysBu8ESg6xjdhzYpzP5/hr2EUCDkM0S5v
ukYU1OTN60+vztDq06Tgwb4qJuSz4x4+nYM/DC2ZUSkaUofcV1BSxDUhfFq4I/Ljvz7Anr5rNQWu
oVTraUp0+k2m45+rIECDH70+0zynXwB1ma4uMNiw9YIIek3Wb1TBzg592CjsJ97e6i595iCPg3u5
EaD5bL1oCtL/qbESETpOJ1v0teatd0lWpj9cIqsycvGB2wYzUr/+U2ll7IhWgy+ffFdB826Of/Pp
SMePUbwWftEoXwTWBom+fB699g918EWVCl60QFZBEAOtF0Y6BIzBczNl4rHwKHbhDpZszls3z4nM
E1j7VhFS4UT5989XtSBb/ooICUWbsXD1kyQL7HEQvM24EOO6mKkmryFq4J7Q5FURV85FNuzIEZWg
GNtADy9tpdqDyRQUpqOLUuJGJ/bEd7ymg3xr2hrVPfVrbnpftZaRpNoRJBG/69GvMTZW9vxQfmH6
YqUAeY1fTaGfVf5kXwECszv64i1j/oxbiozQ35ZeYvr9I0svRW+B1LI0MrIbTXue+8z+kdmw17ua
UjKmkGpK4TSmkJIlU69QyQY9dMhitvkWosPmSJSIl3zRv6T/ZVnWIx3qMJDWRwuJHgKHCPC/Ro2U
emMuYjG0IQUpiDRlWZ6qAt4Bo4szrot0wuwF9AV7JmNlu+oFLBjRAzIp/Ce1ihm7f9yDAT8AqwgY
+5Mogtga2o8nuVNGrJmzynfE9C3OuC9aIHNqnsXn6SzYTirPUF+9RZBYLpgDJRFeXE1SxgmasSwa
6f4N2bLfpQS9cY3T6E6AxLYmX7sv1dtKccDmKroYruAFELv6OuvsmmArvF4ErJ0GJbfT1XIVAMfY
TfTy5sS+8IRJloB+Ed6kVe8Ue63Wi/qYnb/XG9jjIoYargUZWnpZPqZvoM1dD14uvkjkesoVOEIQ
QtwpbDQGrwhLwn3GP8KqAPvjaaVJvnWVUq9JAUnhM7pvlVDONWaA54snBRCmIoVVu2EwTkWMvX1W
qNAIkPw3Fdlyr73Tek7wy2UuAVcaxzoadNtWSgOeRCffkA6v7ojD7BvJPQlo8Jkth9tYfnBn2Hgo
kTPHouvpLHQGUvVbl8hj5lFQOfoSP5//CQnDdHmnZ3lbuBCJ+kxAyKZJMFFj1bcoE1DaI3Rr60bu
SdPcjP8RomioKzndTom3wxe8HdGtxqNJHzUoPWtadi44oH2MKrYOHcGqs6549jPPboEqXtzf/dKd
eOS5U+R1YjlDTZJrxrykMv9qJfor/JE5Q4BgZBMC9lXlP6BET+HPhv4kuXfNZIqQpYYXYfNaZVY4
L9um+3KCDgBRSqczCaRZOibh7LJhTgXtJgShXPJR6eLHJfnuFOxRWcLfPn7go/NM8ilcu+kp9zdT
IFA8EU8x9bl6UqnlCqvQmoTWVn7fWoMZhcDN5eNYOdkNM6MKW7j9FgpahK0cMpI2z+muBHYOIfJL
ex257SV5VtZHfGWwxWUA0fXRwU5wBIS29TN7tIKWp8TlvnFb+yRXgmXp0d6yM5NRdbc6VWM4m+t6
xpyG40CP3XA+fnNHzRuSILBGtEn490ro75r/WSlRN52HiUvwzc0w74FFT7GwleeS8ODpLc+aRMFJ
KL1/gNoU4OcfcC76e/kTaB26VDgEs4XItKVQ3ID/CbjZ2pMhYGLivSJ3w/nO1ZwZPBpj4B9NUlFN
qbG5mM4wNO9ufSJ+oFpI2n7s/gPvgUB8LuIHVEFzJHYdRoj1dwpA5XLUllVw/g/CNnlFuaCrqv0Z
FsK+MNcfH1HkgyQ6N3VN9jsjit2bbz9Hh7DbiuG4hE9UeDYQPYNqQffCmMzgM824m7gKXVhT0Hus
cyDTd2k5yulyD/AXOes04XUudhHxUsjPjNJyYBkwrGI63X8tUQPv6K152yfAClEftxMGc9G45mgK
EIfmKJgXJXle7M+6kKjbK6mS9Qc5/6wsGoWCoyB4XU8jD2JlWTBqI4+9XRbjHQkX/I7lpT+C1Aqb
iddxIVNODWSZEs4I7HtWfOJnE/Voz1zeWZThUF0ocrXwKijuSBeW2xw9x1I0fQu5gfYaHL7V03HO
cM6p1nqxqSHCbUV5Ap/LEo5hDsXlD1bGIVClpxpiWPuz7Bk6u8kRhv3A2nIbgsJocn1Im9DjdXsT
8lqLEJaKaSml4oohVl8gxdPOW6UuVC1/dSuiLZk8swO8xhdtILUulebWfEPSpvjbOSe7WItRmUiH
sQi7Qcu1HQdnIsCeMqM09MwHhhvkRmh5oJQcYiy86+6giPfkXcAh+08dIF1CAlQziHog8RQHDMl3
OYPc83I4e3yZ/1pnZ6hHqWXSAWPrxTSMn6Wcbhl3TO2eTMEa4+UgCLSj3TwkUwtsFAcWe0n5qQgp
ZuUrHH46gM0UANHetcVNpkwS7jhlWBKUX9CxN7769na5gI1+cIBvixmi6BKSt1DcGWpgVL82flJQ
4ibdgoUGGd9CnbPWz3EaDD4raUKYwOZm4rGcKEaRGVngCokQNqKTgnUl3tYYVPpBOkK2mjDIvd7t
U/LtWe58w5cURiZ45j802QUUnibmxU5QjA/s5HIvoqx3m2weQAimXfnQD6fdo6Gl+BVnXZw8LPeI
MPUJlu9QAcpHD4moqgriBY6cbaLGBF/y7f8bHw4qqu134r9zmxtPrOjj9kwZ5MClCecxXDM6YYKD
+8NFvgSMREdz8bbSmRFsbGDRKddadyW8TjeUzfTpB3SVNm7eQpR0i74aiE/LmofZAKdGn1Bw5b7c
g/p2/YvxtDKZvRQpje4UpdXq2cmt059wHJCAP5obUaupOxTmD9rv/UEScjpkZq0Cqf0bujk9r2yn
FbMsJIBPm9y201OGb91fiWEsQbCsrqVr5WfdQa9qKkYEpF7uMo2dmn5+Y4gpQH+z99ALv/tP71mz
IE3Yxo2+e8eZKu7mvPaZd+xWjFKwdWGEfqhpvQkdtJQ7h9XEgkx1n5RmP4sVE2H8gtxiYvoYHzIY
pGBwhRjCQfBtSw/Kvbf7KTGAzD4Ja9FvU3mrsKgaGP1PTpF9BRySzx4fdosdgduLn8tMjBV2utBp
gDLkmeR1g/xTplA6tAHRL2S/aOT0hhLR6Acg9dj/Q06TwiuBs4ezS0TM3Q4gLNBb7CHuI0guw3p/
A8zznx4a8KmOYSo9fm612fqHOK5jFHY/qDOglhe9i1jvmMEN0QTsjcjjcbO08Wrzeka6dR6mUBwG
L5Zg1AGELxaaPk43buh8+VgHh758AuydLM6jabnjtXDAwjgF8Y7J7Bg+6M4qNcga9BjMBxw1o1nH
50OUkw9UP9eCD1wVUUV8CuTxBLN34F9Hw31OSZ1AKp6VHN58nZh1zzgLcR9AvzH2UUH8jJmBrbHG
6RiMoWaIW8opp+9Sevx7CGN36BAy8u819N140qCj4+rAhsTbg6D/paFLbXkNycMtZY8VasDEd1eK
K6JV8pLqpkI6dNWX36fyof+n3Pbb/5//MwcuhRmtI+ELVJra324rPJRc1Ysb4iVjBk3SRgp25GJa
tSqxP8e9QeG6Dbo9OCk5wrZmjEoZ9jQKWfANn9diNh9y9ss1dExVZaNymkckpXuOFcY7W9K87+ga
hhxY05PBXFV2FpZXpQo9qIFKWMeoEZvf8CiTv+qXJzf9z53/l7FyxzFjVW+U5ktuSgRHzJkCDn0f
UsAmjkjpzxxeo4/3AL9867JnDfJlVYeZj49TQI+8npf1eW75H4ZX7YG8CC0EKx+aV2gqrwmsDe1z
zua0/e/nv0O29009SfC4fSL40opBLLVbSt+saViuTMSZ0M001poT8xj9njq/LAW0shmgJeKfsW9v
2YO1Btp0GPP38KGq9VsZU4E7VNfZ1w2JnlVa2wTRpQ7u946bm6Eq9aMtMf9fCGf5hGEC2kMgmDgA
mmQKCAEsuQUkH0z+p4wlsIO+1qY2294qExlq5KfrpDKw4g/zFZeF//HRN3QUp26k/ohFxRqYiYEc
Ma3vOBi0ntxaGexVNGYxyJtO9BIZQIqyH7tPWD/6YADO2uOSdSiPj07lIqvCcqBN9oCqNzwpYgN7
IGvkJTgakpmb3gUQzfv9zP+oSgvvuOu8QFvowawpYJdh/KH3DU1cmpAp6jC3hXhHe1IrJ7uK0IST
pl1JwSTgswxjdlNWnCQ4UtA59AKiiCb5lLV0+wY+vpXJkoMHKQODo734n5WvagNAlnIjlJLaVZQg
x4GVi26y0tjI8j5uxAIFnDnEMpDzx+M9GUQ8z8AXl/J5H+RsX9a37jfEc6KJ4/R7OSCIXBJQB9AD
R2wD6zGJKK+oEK4BN4hNMPzAlvH58aclzawS6TDhkX2gAJKhzBaozdOD2IfVSOx+jChFDum4fyku
ny1wxEMU/6nC0Bh5HG5EBRCJ2u1Z5mc4dNnpIYaF/e2JkGK32wVuOXjxsNJUgCivYUfd1aKR28ZC
bExgE7SOKeJNyjBesPMNJsU4mNBnAZCqIwIWhC5PsVXZIOOCP7RMX2mlBaYEWnMS9G01khRv8Fpp
/rHWu4i7FKwaVNeWdFdxn/8dKnGcNKyokb9XoO8T9BglezV+n7slTA0drzWPwirgoLUNTf2C6wLU
uptJ/acp31GwZbvwjR3tSdeQD2hJ00nUwaxgOujLWfEkQfoFsQX8x76KPDHalXkdwkH68tNY9R1A
VNXZgQU/hzi91MrmYYXjJ9m1uMdYb7xKbDMHs9VbLWQqOhvfeXgUytdKKRP++S1fIKbCsmqsSqBH
ET1XoWkIbCVsY/89+Zooi55Edlv2lK4H+5Pf2aUmNto8rRnDC44PD2uZnaD32EUmDe1pj5uOW03a
E7v7pFHx3qcpQm25K5LgBK1zdVgT3fXjZMN1YQp0RQm0H9IeTaH+lNIpaWSVQ0Spv2v3k3218xZf
3wJ2eOUFMh1iKnQVEwuaYbpy1Cjn5OKtC+dMXilrEqOa9YLATYsNs1vmfT2JE1MaF544SxL4OTxO
PeY78rg94WdwHvgACicFHg9MDnhPtxpGTq/n3CI41wMpdr3uNasp0IF4Jve7v3FlqWM+sMH43s78
MV9Kd4zvhZNt9bduyoENIHG0V/IvAsA38YDYOCR73Wv3KvbYRxiDE3XgkFWvnmyTasUkB0nNmvHX
ezoFp2Y+YYKZiAVsYsx80PM1JcGlWhOQ2OFKvwL2l9SeVRiwqyZ55QeHYBrYPbk7AD3oWIS3UqXT
qtC58N/OEb/o81X5beajm4ea+ITZbrHNTGTJfO5No41w2hn7yGet03KxwvDxmmTzSMup89lpAp4n
jAOLA+K4HRmZ3sK9zSo4YXZoWQa3vOD8QpnInTYIUx6PFejcPTIxmwQ9TDA80SV9it8uHfMFcQBw
682JV27mLljI+i9rRYiSwkHUn1A4s3VHYCpHtUPRIXLXWYzdZ5xfsQFvdd+xp47DeHEh0pNBHRj+
ZIDaxvCdkXzOmhhAnXWS1jgfYeRok7Dn++wBUzrTXEImmYd18f2bplA6V4ogW5f6M4FHuiR/ShDo
uPnZrjROwgDO770ss5K+IfGoKt+qhbjZPd1SzxZkX8cb1JF7VF5h0AIxYeCYMDsih9u3wlc7LtVA
ADTkw4aSl9x8EtEYUHMAxIyQkpAMT7crHUaLGwBAm5+m677JL8gW6t/qwqO88Ey+ZFMlAO8WcnJa
T2uQNqUXa1+bF8MI4cqfMUJ+Vt9+fTuUbbYHP8fj4gjHUplNkeGjoISEMQ7VVsmBAu1HKqm+WK4p
eSHyiqD1T1udHgoywG5U7d4+HQZL2Yxhf2ccMSK/CN+hvuzgP3jfx6Ozgz4qEnEuQpaMuRkS1GRB
GO24YSeKqnahSwHaSY4pUEkLBnG/+AXZkFvEa4AU4dZHFDHt3EmvyNUFPzXDjY3eWJEcsBaEmcwI
fAi9B7b4mi8YXgTenEpX6xa+ClsiM+v0EbGhrAqJrz0Zku5YkPv5n+jwX6dEWQxNmu3XKQ4Agod9
I0woMNON5wJh4Od5IxW137A0SwVsALN/OaJLT2O+e4ian+NraprFCY948EjDR332xi0s/lG5K7/b
bS0rBsHfBvdL8twf+lSVuScW/BnvqGe0VAhuBypT0P53xluy0qUSTwhsGQk6izABt3S+De409Gn3
xOR/ERFc2qu+LXULv2z0KEL3yJWrTxAzlFzHASQxTu/hhbWhqsVxFBg/yz+DgaOG1AZdCRTknnr8
XV/c0YcHWvA5CpPLCdPtbrCRCYlMJ2lrZf5E555CUMJHZbgb9Ah1sI8a7Qo+iDflrlDlTgfbwjcG
c/W9R85SA3kbzrY4p6JuN8sbQVW/ijjcISdAn2dsbEN8Dixg6zRYGL31+TCxiHCRsr/3FL0YcyHF
hPikzm371t3+rPQ2cTv0Qo8pyqBti4mmEFUywwV8HlG2l47LUVnd2/TKdcN8brBTroq4+hiYnHek
BVyHy+NFF88EXiufW2EYHG66IwXnHA3yuIvsIfsnDOWazzjCTSgH/cKVO5wAZPPFFhc9bw2feqnO
mFzgCruQykQiTEJEEMq0NuWZTrHTLfrgW7u20oSr/AE2Aisj7NPT+AUwhMCn1+rWIVQOZsTiq9ue
vVFKBk1aFYOyt4fvwqv5kLibZ24zuUuhtAuAWOG3ihPd3xvjIa/9IF5K/Bcb/skkMRZ40kAZiR2h
ml81xspZCmct0U1WyVt5C4tveh+sVw6u3kK4trD/uUuuMYaK3v/2RgfwfQTGvVlRUO/OFwJRwrCe
tvZ+g6O3fHKwkH3oIH/gjo1kE2Av1H/tpRHaq/1RZ8f5a7IFHkJa/ntK3GdlUBYNie+M5PuYTEMf
WmZn6koCqgZWFV10En1eqCORJ0rqs+WN+zV5hnnsCXL6iLWhA7OxpV2c8XsiHL7JA6TBhMsNdlov
9uXWGHFpCNoCkB/R0mkRUW6YkuI3LWGYs5sjqR6s7Qo6xvdSwkehEjXiJIvIg7EwBPrH9CK/fIvC
aY2LX6tuJQuevHXonoJ+x40lMlJHIdRwVdwFxfmO4P7MmTt7MnQSOry2O3sCfMIWwKNpPTmfxRAm
ZRKKk7IXcvDqOVVAT9klHmRH8Wi2bVAOEU2b6WsKWwzMLx6IwkChOhe55NgsS9JCoasZ3JnWyRQ3
yQuIwMr62Oj5UjXavHqWThZPjrMAwIPLVUsCB7YxslYUNQdR2xik+0hmKsXj9fo7pq1TvjB4NG0x
6oaEiRccO1J5dv6DjaOeUBYcIKQp3u9fhGnVa781aHLz5ZyoE6UPR5yJnfhlOl9pVkd/hX00t26Q
uJW3m3MmLlDa1k9BV4AcUS3zBBRGuStINdkZEIT1JC8DXrgccl7C0Da3qtukVsSC2MUAITKVrYrf
z88iMX0vZY/siPuJ//F4gFibCqUUwF6QvSB0NzlUqPZXsKZKNb/L28Lvyik5hcGRQbwIhuIbKFFf
IQ8ZaueHgSWZ6OAUy1366mqZ3sXMx5smGi6aVLx/GfYAgAkeXMxR6fiL0BzLF5LdwIdocFe0KZVH
ayeqi6XGTltI0qhxYblyVst73lwuJpe88ep23cslFcudfX+i32m+4yEyVUQ8CM7IRAIYEaa1pgO3
1YpSuS1OZjOXEBcjjMZeyBYwadiCAhKkLqvWbhAb8JxbD3gkhoaWd6nhrpqrmL1CpG4eWRN91sv7
qd4t+cElOKzD+0E4kL/XRxmYja9ER1EHqZRJFGm/eQiVt0fM4lQCJA9OwaG2STazLm+enFBlGwWu
w69qH0k+eOK95KQkyT2RnPp87NlOc/BQVk/zmBxZMP0P4zyuDINI0/Alxrii3hMCRsskGMhMsDuU
ehJZum4X2ckBJUnEq+CC83GY2JbmRA5LmHDsOXjNg4kf5y+BqIhGRndJH0DFs67/Nkiw6HIkmrVk
Fnbn3pLZvAV4B1gcZ1KYC1FY/99GiC75ac6oMgiRb3XvduELLl7vqyq7yfAxRFRRcTJPV6mOuBEI
PFWG4UjlbdGIPen+FrGteIG+khmazoHmg1kEbXjtazaMzKvTW80np0TRgFH7Zd+NGW/jYGW195HO
3PtlbaRNCfjUYa1q7rHIz5yqE5Lj7mwBgNPxcdgpjq7qKYJxcr67FSLpWCsbJjZTTUi51xgh+PHL
nrfcFOLv3nEuwE1gHwCAqhO+CXAp7gYJnmByu0lbf4fiMZj6xt18ENmMI49OtMFPy5q2kX4RkC1l
S7T93htJW/eIvz9em0UxMqsEhATvHyxAI7YN9f5cT8GPMdszZd7VOSFWd7sMdU2p5hOAT2D9PLh3
/huOR6BrXwPJjCaJ1U0Es/wwmAfTNxtUL5jZXhLWJjBbgv9SdthGqj3+2+BJeMR2QekpZGyF1wKY
+BGrvRFag/0RF/m9GQUB0UfHHdLy7nJUwxgKW3fJUvImN7+/wCa2PiiFyza+8zw7IHQKCD4bqOQH
M1fhfk+wUv20LcR+L+b+DXF/AJfqNIWy30HuAkLR/lSqZw/wGkJq2ZPZuDlsBoMC3RoD1vRWS0P1
s7a/StPWK8sksj+WzRx32+G6lBieUtYvOvVzoL4eVzUVaIUDZsV9t/eSz53Sqd1Qo0IDieJw7cQM
dVtvr4B4FQD1Tckh7wtsCa3XpEkj+SzSZn8muxcEsbd7I0W8DMmpbAnlTIecnLrKpkrIqVsg/1ot
4tUSuURNUZwAyodb37k89kotuCziPnVhyHx0EHyAOCW7Ev5/DSOqoRd9jKKD1M3tppcG2zxD22Mt
VlA7GYVNQlPnEFA+r4TYk8SEmyWHPZsMtPfzT/Ns/7pIxc/Arz6MS1uthFNZqOC97OUPAPP/tEz3
dMwJP/0MXnVeaX6538DfX3uyyFPvLMdv4e9beT4dMf4UkN84zM7bANBGjuOUbPN/oNAcNKXy2wVD
Wvl+EQDs5VC30LYaE3Teg2QEoJjR/ZA0v0IoJMGRYvV8ZMG2HEAJBCA3rTZmgfMU9dnpw8giPgJm
G/V65ITLTU5Wgv3deZ+SsEzj5lDzDlik/54irRkg70g2GG2F1lXWdXaBkr0knRbMgq6XMwpij32K
PiMbf/b3py2xyyampTWZBYPtDuLzGERB2yZNq44ozieyUW5ulLpZoWvZt3OPzpbAMkKdKmfCHQby
M9DAeG1exXugX2k7orEI1Dnt5b/zZH6aQTHWhFTd15lJfgYLGYKB7wv/zDy1euqJb/fZ2zYQTtkV
gwUz3zwfW3V1f/bgFZlSRnSpr1uhTp74siSm+LivfAXbLoakA5P7T3yDAZ005EhoTQ5nD7yG/KiU
llzCibSyDFOKSJD286aOvK6P93RAeILZ7Z7BRQuK3gOOPUmJ9z4/MmTqGFlZZ5p698G1UHnbZBzf
JpXK0JREaV5cHjfJZNGyDkpdR8aUaavejE8Ut/wTfJrvV35pkabKnafHlLQ5oY4kf64qmXMEnjHi
Nv5MfY/bTpdylgI28Ck1cODSihjrAw9zhFJ+sQXZ5bPkgTPU+SL5DCXLse8RiGishJIiEPV2KfhO
W2PdJm6AT4cK+i+VAv4DQD4eyh0oV9Ggj1ty/GRZWILsQLjrzewvXy5DZBJhiEoEIfGkwDCBosLb
SO5mdIKJO7K7U+rH52b4QMK0IZdvag1DTtdMUJzuEeCy+wtknhN4Bdmtxz00dSxt4zq9M0vHgneq
I+kXTZ+8NdiKkwGdJDccS9tPlPUtQHXux5nV+UBh20QhGxLi/LUD69lRDS/WC9M9E5g9V1uu+a8V
LHZnyNSIDSmq80GgtYEuMWeDLRPcEJXYkyswAmzGFzJDXkQTAeJ0g9qlQgdnkQq5i6e3TdajtxO8
LEgL3Z5cDNf02ipvIDKZMt9ucBKiUnD7RxggWKdszLeSUNaq5Kf7F0ckYyXsWADQVJ4nB8QGzZKt
ViFT7zDBUkb8amD3kIyCZHC+kviTzWMYPIa1czOWDFaebXlV+YLyxL4hwcSPctujJvk6ETzboZIW
BKbFSM32IGpY/yqMi2kIqKdia688ePSgqV49J+2+L0WpZfDOOET/T98sZF/nmnRbbEFRvZRpob/K
akoLLNc1U2XEDI8z+6smnJWjIPNbHz8VbSSK4B+rVbmPq5tlBX4aAZAfNwZPnhHyn11PXsfP2QAG
1eRZClAk121ZBNHf9Tp1uAjeg712qjbVzQ3oumuvY5tnRiVxpC3QPIgKuMcUU3Pn0vCDBPZRQL8J
tLbavtmWB5MUwmX3931QR8d7FclUlz0ZVDlo0wh+m0mMtmvHDhOLtukKRwu6Tl9mnBEF4OpaghAP
2LWJOg6SiPfu2qf4mc3giJG8fDbO55zq90jIfKbSlAA58DT92NZyDsaqeaOB5xrU75A8vgv5sGUZ
vikKom9RKe/RK/p9OkI/QzEyEHH1izpUmrfkDa8uJweIYi8iMJi7i+ZvUA+0ixtyn7dpAGrGhiQm
owocyDU4eDKifMk/Cyj/h68gsMhH2WARxEAvDfgdM+t/2mxfpImW7IHUrjQM0PpYWcCyxR8hLc2x
QkOBxkaingklfQ/eHG6vc8aS/YYSngSSYz7kUyoab0b5Jbu4xwupC3so5ck/kBfmWu853AFEar+g
ye+U9bNXvWapvI7RNjy/WJpDjbbaQ8tsBIR6ZtkAHqtyHdy8fLF4tt2MljFhGbBeK71dVUJZJUGn
bw4ywA0r4lK6AKQEVZJM4en5KfJwZmrF8cOVb3ybd9Jq1BxyqsLySPexXIXcQGl9ALwbzsYPnKs3
3KNHOfKu1HbkidBhSW7IQg0dkCqRvkF+QdnAyEHnK6p92BAzykESfn8CXQGBaYsY/8Z3JhGYYKut
0tDZXibwmxHV/IG1EI2qGHmP/LHoAcV0pHp+EYpEZ8QsiB4QRzkJ0YSOS8v5ifOmqKIeXmNVHdyr
JUUaEw5PdB+2UOh/BdkrmLQFKqzwy8DGSiuar1/ovnmF+QwEHpBQydv6RCMuCexCjIeEdpjaghUT
O0GMwsRou8+8SuB8MZncl2/HKqM5kARr8bd+zWQNWO4CPgB7GirCX2Rx10JFJDJqtCMxIwFQITAU
+A9yAYq5U7QD8zVrasFC2854TbIzeVdd7VmKY2PHLMNjTlXAS0XXjhIQ9RXuN/vmnscrTfjA5bYW
Zp3bIEPKPS+6LwR2npijrpLY16JCbGPFfhBv9Z2EBpsPqKuidirEPgtFQc0J98s5PDMbKQSnCL2s
MYqRKPhwfCeIVHzrF7oUUPOpgIKQB0dgxqvObyhLsYNBOeoGKABbws5MG5vPEOYDj0fp2WBq7enN
2Cb+KxWQKb00JvKvtlysdoxNlY8fF+QV4LvW3SvzTdk4XrjDsYo7sFk4NNK6ed8tZ8MoPHjL4TbS
8gQ2O7lKlBtPT9JG34tJbfzhD9ywrY/a7oTOlvdjgVSDEfc9CYCDITlMZowgcoKZt32J2dsQMLK1
Gk35R7FOhJHzP309HP86/i6cb7bdgaAdLa7/O2Op8PBpTPZt5R11kflGC9/BEPtwuXds489jpuWW
QRPpCDsZ9AsYdlAH4E+DSZT5C+5eeo/Ty8j4+jhNhse3rVojC2wlo5v1ZDJWXRuMq4MfyVfcMQU+
R9xwJb8vQcDxes4iHuN5n9HDWdeRubebr8DT55nJFT6+fUUYQdtmlu7NyUjmMS1deoYvIk+jLuS+
NDaDAySgTY77nkLYykLZQJh5ePvMQUmvlo1j8ZSA31wJqTuQxWjmo9/36eHKfLBfnbUbUROMC0Ft
bp+Lc/FYa2zj33Y0eU45W6Ta+iaISX5zpLpM3tQ4FqoLC82gGA7D8wemy+wtXkDe5lBfx8eXQowC
sL8RC/4uPtVHQkz5aSzoY6OJvl5692KZgXKZB4e1HKYQ73Dce3OX5c2drwbiBmJc83Sy8ypB3mEY
L1Z3Hg2zqTS2NmYk1lMAR+T18yXGUxxwsYwDSyo3xjJrLybN46t6W7zmnWPdqtN9NulvcgP3zS1D
wBZ52skxz330nCPvxqtyscEEUJ/UxK2dRYUd1vXjtB+UqDIhkOap9HsLSFCZOXcM0G2MgXhrdcxM
66jQMgOA+houTxMZevjo5xTjXI4jqeM/6Y+RD7/Dyd8mkN+fM/q7093gJ9RBHg+fcgt3ZbjxqM3U
ARch+JLhx+J5yVmtqZVDidiM8w8k5tzQMaPLng5XBfiOptuf7hDgzmfNMu8Ct7WqOraqJTWs4cSA
UK/gJ5JXWZWdC0B2IQNoHZn2G8GXGUZS7iP9+I2yXnUAzgKmN2AeHAirZG5KEuuMklhwX9oG8VbX
9zzxubCTDdyjuil+KYehIPeiam8V60+dItThm1+yeKl3KK8DONsgrHCv7XPzyG57RWf1z1VEvxw8
Ep7bkDK27g9YIJTUlQ9UKEizP3j1Yw75TYVTjCqJKqLJ5lUU7I3CiWoqqQRume2Ijj3rkS/xK2lH
9c2D100rrTwIC7/Ia8cyEOPF5bHKie5neVd1GG8xKwvEGR38chWmlKiYRSLe3RyH1BHvSKL5ESyO
Kmzxucl1JEFIoFM4+rBe6qY6Yt3YAxBMXqV1J6lZazQi7WLo0ITS0uqa9IRdWBqKLGcvxVtfbQ5f
5vnKAU9ArmX2KjdK50Tvip9xoX9+hZQ0aHcd+p6BXxns5IlyL5Yp/31pU6ngtePmFASTyUOHFA1V
4DGoqrccNcno/SP++IPMRnSOTqgGaT1N+JXW4mgQuMFOuNwAp0/rAWuIunJIi6ShDLsQEbZ5c12K
kyFvdtcyOLJ7dtDTXwLEVmpuUOgxfxHb3cxfhkCbOj0/EWspuap3ieEH0EhHmDf9SrcgELSr/Pvz
N2hW9xnfzAN248ShKquSDXJUW2Czq6nc+8uA7MkHt7kTkPwct2PTfNWQkjdJsgGF5nOhUm4g1ly9
1lDRBMCWxFC9Qazgn7Z4mfREgZOIh+j48Gf3avjPbaLFAs0hmYuQvlnKlA4IbFU+QtE7/VQKlCo7
9J3dv/YthSur+LAx2Y2wHhsf02xa0lCbMA+H0AI6J93KHrF0VtaDoisDYzyEd1IRfdZI6zA0CRs7
ibW7e6OQaP/NfbgZJWMrf/cUCqnRT3K+3a+CktCTBvUyyNqZYCgy8ANBYctWIfHOYSjy2HYVZohJ
46IRaRwnLdlfRRbhNYkcaCeGTvrxjG24hLGAknhhMkX4Gu3g+QfQzszXjjoXOk6aVG9GP/w5nLhf
2vQxhYK7TlORD2S5elrw4mkegoLIoJkJjbWaL5xDzbXbCjsl/mFFk5iiekB1VpCJAtKApYLHgMZG
vkEhhXsu4Imrca3FRfni8h6QgDlmqmKpbSTsUQQy1YtU13pDeUzwYSkc8smLJA8oLbsKXbwlDgpT
YdmA9iRjBzVvnUfifNsI9DofBwsBLqo9R2pQfhiUKbTkYyvpQ4KuISQ1S4oF1uMgl9EGai+sbsIB
fKdYLP/u4wAlxxxOPONS87Wb0YWLPZJaXkI9qjf33F9GmhAFA1bwpNcX7yZYHL+bIzrHNlct9Qsb
pKydyikpav+v/O70+Fx0Ds2sXXNIWxAv3u+H083Av3iKcaiE5it3wlvyUb77LrkhjplYyG+RNg4F
5TwxXV3Anuv2BZ0K1F0SV3ucQIgJskKt+XDp6oqQSX+R4VO54l94ZJNxfDvEF1l5r8FsJiXRHDv+
6qyC1Vnf+ZmWt/5khEnsIaCPvdy1ykSOpR6F261Yv3o+/G06z6yjEK/WnQD1Xl9o7Kbsl2QGrzZn
PuPhN4vWxJdXQQHFNfFXwIYwI3DRmi8dzw8Usktn+GS4ny1mNqCdiaxRb0B6l/R/kl/nlPwltqiM
czFARJE2/orM4sQGXza5/aYPEh2sc1YqTbwVzYL1088nJCRnoooEH8Idlla8Lts/aTM0QorSj1q+
vww1z98mKTLI8JXr3QrP4Z0UmBSX43B1MS39rJcNBYt6GEaEAGFHoh7VkJyADk5h1vGd+0fn4jTq
HNNnl+k91Tg9tKLr325SZcp3NSSyjPHk9YPG9An5Mpuud+UcYvUiFSji+ejYE6yQlHQuwTfPiat3
fc+jph+2VoaQMfiPLepCl6obOlPKTeAXHrrj6q36WVCO1GHlCAXcIi57aIO+yoIfcbl8WKe2NI3g
xJ894n6UrRF8rz/M6lpnLNZhAA7OTD97wvGpJMC2rKMsuqg4rVDwuR7zixWPpkL6KidoF8YG6olj
GyfIPOOcbemZw7NiskSyNjf2KpyipdjBHxxcWrkDIJyTmkB4RoTmdW3APDSSoh3gHY29Id8y3N5k
5jnTv6s0oSZvA6Qqr/xKXIavC7oVvzKzUpdEvtOJgJejMiS0lcD0SbnCJCGtK2hy+cXFffgppG0F
IunYlH9dvC39vt6W4AEoYBgdx3v0UvFt6mTU+8LLIFNYZm3p/7BTSPiEb6a1C3VuLCBGUs4tyAnN
5o7+evdSa3s+EdaIlrh0qXFPNTPx3Uqn5ULviq4KoIpkMJkqqQ+CqsLARA2+9e1AtFUt2zb5N/bI
wHB1T+I1T5Be+VCyocou+2srQkO8YCQhbK7Ukpog1wPNIw11borMYyVMEifhVpw1dCOLQ3FVIS5j
tKk+28du4w9bt5vUNnlTf4LvpY2D/7yjfj9qszT8ZH7SgEifp9KGXns1jpFtGo2r2aCeObPFkkpj
a6uT00yv82TMj4Od9SRsnRfuQTkQEPvjhgxaOW7vi6uM7YF5abyvPcArWrM5bbfhwXkDnF+0n0uj
t4PujXZRR8ELlRFpe3H4+xBDjxH0/DosnbtjtHL1AKiGkufd2CYJnkXPfrRJVTM4djil9AwKEVAQ
OTJa1qOoBvIuT0ef6dWT14rT8qRAQVL0aSVuHJtKoBCWW12fNI6l2KgzMEoLYo+RJ8SRBpB4wAj4
/SXG2tlrsr9dYJa9FUoYs2ctRlor9o/uKXRbf+99DZHiLFM4y17bBVqzgTYtVjR4MZ9Nnj7gsBDt
w2MlbiNDPMVVIh5QOgxDYjs0pSkonOSFHFgRY8TqRmoNW1mFSYvjusAt4X1EKnZ6EyipJdDiIUpB
uqRVSAjGudzf5yu2SPquX3GVzWoWM3WWNl37A3Ice6kIze1x7Huthh8P8RAmNL5ld/HwwsXoNjWh
VM0XGx3YKPhMRbAEwrxrXrttn2gobTXxaFDJfiTo5qJeSqfUs5UiCJsxO5jFyBN0SaZH9I5kflxq
Xj76revzy+7YmT0WZOe4D6/O7niFJ0Ln28aZpocNvuZB2OcEdix3B4Gb3ey4DxRZMsoWdDBs+5WF
+UP6JRD5JZrovDIImktpYC5ZSnVMgu6kOvCaR+JpGWCja2HCG9X2gnLGkm6vfwOlMj6wzonxX681
+z7fJLRofaqG4OPzG43u+GK6Vq3iti+insmeV1K7ywFHfdGZlO7yLQ7UA4iOS2JgnyoP5IpjoK5q
qYKLnVqRJQrolGOqWHf2a5VCmsvjqxVupWOU9brI+LsKMYDDtcDPO5l7+qixf7puoyHndhNhgq5X
6KvAJzqgf9LDsS2aVgUu8DQD1CRBHSOCNR6B3qOx/ad0BZ68PXO9V4ujZ5rUtIIsQT4t2JSpjlzO
XpIe5nEcuk43JB4IGBUjEIEq1m204plXmyvrOpv3UJuoW3KkLGZNvb5zqQKbHAoCkdIEbS7li57m
Mpijlm3yS1K/B4b1KgCAyM/ITTTz3a0v1Qp728hAfrczOD4nGYh0mJpnZyiFFcbNfpJfhFLILmM2
sZ4pdBIf9u3Dl9LSaUue9mbiicWOWzUKlrkU8xiV6P9hRfZwEtjuexFv0IH2KFWUQcW0WKfQ2d1W
aGQbsipWAynMcFrDCIXDs0OqNCIlgZ+Cu3039onY6q7tz5a9kicAHPDFVllkDYTe0Ep1vM8EbJii
Cn55to1/6d5pG7fj+0lqboWjm16wJriAlGyU04NhSQrtXctckARcUVnGOr6361KASAjyvccfqzUu
gNVmQKnB+ZqEw/ssrTGsaha9bpP4JvPAXWzToCJf9jD9Hc54qjVPwAb4gstQevWD6QoPBIRG7ZzO
6a5pwZYfCYTBXdShvS1yQBCDdZgqdlbMk0OQBlSSm4eMeZrWSUMi0MhOFGf013Re5dxn46F3zUcR
IjNbzqQnnj/RSbO45TjJFoonM/qOrKaLGB4SB9TiYx7aZDnQnmW+GROnyQSqLAzQpFfJF7FhSCjg
sjfa0lEfVQZ0FmMOfTHTA4gsyfdcJF8rZ+qoSR6nxlBA4dFVkFUa7W2XLQScT+Pgmw2J37qIoyy+
ODeYhEMJi/5rwQih77Wzr74PkQfSD7OO9geackK5WuGomcc3ANtz3vwFXqUn1M9qbdFUDH0fhPai
R7HhAI0HQ5WnzPDhduzv+tNB+O0Lmn1E0dwOeuirXEHFRk217kFDG2+Hmp/OibWg6rNcj+TDFHQH
ewonxgwSMzlwRx3EvS7RQp7fo9lReWNE29YQJLckVCQkXYNd9xXIUqmZ34JY5dPiTypnOqahNpYY
27d5YM0VeQoqKZ8IMh9Agp6wfrbhXeN4O7/3I4wmIRaAYwK7XGYZHufMPvUkLqC5TQCeyUOFBT59
L9cCOR+3ABcAUKnzap1gKXKHTN7h0zbdfC31vHD3CNgvVQHZOI2+8mbay2zuqjAebUferOO+r3s1
XT5QkYdyVcM7kh2v5dWBzqNyReOOrFSXlY3q6guq0j4dHvSVEObTnSwm98rhCaaD0/s16ltqyK7x
kPrf6Y+kx1M1Cs/2yFSQIxcuo+09j/v0u3wBAcPepGgtU0o5gcwE3zaAFecjYyX8wDUdP+yF92Ju
GzD7pbcvcIT1rI3HAnYvugByH+J5Jeq/vwF2HlyanHRUGWCzl0YP2SdmjPb0klr2TcCyoQPQg2mN
SZL2/F+uQbe+Ynm59QPl+90aqHf218C3ALzLqhbQEYB3Vr8OMmJJul1sl+hOxoL+6d1c01PJFcb2
I5BvcfTAdNipbQO+borC/C3WtVSknB2wfACr1G4sugq5sBAtxuaHoh7/InEuZBN9eZN44UO722Eh
7IwZqe5+NBEKBsZ1gSZjehEYLQ4HSHVdF1i0d79SBDf8kM0SYrUgj+q3kAxNqialquOpJv3nbk7u
pENUYU65xXwXvAJFj3mU57pBoJx6GNd8c9wEOPSXa14b8Ut98DAXn2tCpvoRBFyKAqA1hQcw5gkG
ljV2f+k2egpceiEUcKtJElRTGP2kHnhhQumd/Nl5xgMIiTYheH7b2oIad3DvUi9GROkDbmuPpDv7
b/aBNdp97o3cEVxT/ORWn5gxhsKADuwWSJrHUpU6oNcvoFkNOdG71Fv62VhbFQyv3ytg+KTKNGLI
T6bkmFauics6xA7bsskS399eSjfUQ4PdaLcoIv7d6ryNjXgk6sfesySE4Ka7XRGyf/PDkyjZnjE/
O1rghu0y3oHHHg+JXRFyu5yZVjrX6gxMqAGeK4A5URCKakOjSDYadP3a5JjlraIOWsBOuquNh2/D
zXVbPRBgMMB49CRTrPtmFKWS6Yf5irjlaAfPJMZzYlz7glX5IKeTZXOvxFZmPOrJIQRRbNeLSgdc
D3CUiAqcobvXBryAJTwZvtvhtUHO5MAhM7nQtvxCu324AfayOZkySPGG2PJGWN/TcV5ez6RYA00h
Wkb5FLfIufnUjdrfo3mlpCqYB+xTGyc+0P+uKHErR5Dgmme0Xr/5ufXdyoteXGVo/q6mSdKMJOgx
du0FMiuI0a/RU5TfszxtIdHkcJz4UoTpKYusEQ1kSX2NPPK6CrTfBgtTxcHboQAT70XHdbs12emq
skSBubpPxQGUuzqTVHYGY9l4AQ+Hm993gO0yX8ko3FJ2D+WJ7kbEK0vpF+a856dsHyDj/hube4KR
x4blX3rEKGgtP6jDty497WQnpUDSo1gYpKYnJHcyiyOZwp45raUUcftCPch5lY+Uke0Vd52VF2S5
XlARr4jcW0fQXwFRDQ9/v58UiMQnthm8C9HE7upgANidguxTs0sD6+k54eVYrijLpffrKSHdo5DV
9V2+T7Btk5+w9RTKyiPJwJsy7/+BlitFUOtLoNbA/Yfj3N4hvd7uVHEr6Jj8vr0HT4DnHIpRBQ9j
3T6kyBP4RoNwjGf2gJAgeRCvrs/d2Q+Z7kBd6UeuFPmaiducu2ho4akU79Ch929yTOBFw+rC6dlg
Lz1YzIo5Qe9537KZ5SKpKqlvStC/BbCQK1Mx8PcyuZhE8SBXFYbl7TuHVrY1k83lfxYf0KLxsRIx
eJHRUN0TLZT1RftOLNDSWz3+Ki629CmDy8GOK2TqFyozTVO40gjVT8BdaNjJ2cVikHYXNEylvF4d
cpuxxm+T3ybFS6BJkQ2ZQqZen5O0NGzrXaEWCOONbDfar8t0nHBmn4YSdpQtOW+rIYDTJUqIfjhs
nHN9mMBvQ6F/6GPmQxj/w3b+xe4pFN4IzAPsGpCKX8fEppRfT6NXmVlm+VjRhWzFS1FQ4lsAPERV
gQQl1Qw5bJidRHo7w8xxWQUdKawIqucmMTOFI5VtwqFQt8HizXFgqU6/oSClha7S9gez0QV7tTJo
3Un9BPG3Z3FkBgTEirpGTVY/gXMPJHbMLS9diklTytMX+Zp3sixrl/MzS3fOR646Bb2AlVcFIpAG
2b8LEz8Ldi/8anovFBxirwYPnwdQH2BVjIztArrSsrA9KeQgvFkSZFSUupJ+NnQVDSBXgulK8i4e
oRYRmO+RRqPM3NR26zRaahpBiDZzH2yWE5wkZZvk41fWl5CGKv/PH2QCJLXkWdE5/Oy4R3iVSWrh
oCReQf+g3cMgQy/uq/4FZS6pLEehz0G1gUftv/UF24+Tx6MSNxmjl6Ov8qR9z4tDLZ1yzxQLP4/h
YzlAwpaSkqGtC3qXTV0C67OeNf8F97w1bCpI9A8H3gW6F9M7TjOHDAwwm6uKYRe+TmYebVjYRq+P
koSERNY/dTjnYM6EklnAVwPVrLtTCIgRnf9XG7x4UHorXtg5+Jufxg9A0l6o1hcGMEf+srPcQSdx
aMQpaVdJYZ0zpzyiYpcaVA9v8RuM28CiQqmCxA0ntsNPi913dMOHrIqF7WerF24j8SEJnYaFiFBs
HxmTarfI7YT08yeAwgoWQWX5p/1WfSEZ0UBzAIaOVV0rO+Mmc5r1K2tM7oevBYmmLOZmtJHZiPkh
Tl3GgMWvDc1yVsGjWdLpN0kku4R5E8pgA01aOFaI0ERLnkyOwX2PgqMurRwJvsxV5UQw8Ju80xo0
xfTYUaHjH6g/1wCGq7MP74QkFBWbyvFp2I2oaFDH6hfhQjPf35Zjk0prm9u3Qr+7RjlEuOXBDThd
DP4E7zwpuN0drJAQ4+2480QIEn7Otrvrj5L6Rn6ZQFYRlmQvICRhrN9oaE5B0GnvD7CFolbT90cy
JcFW/RlBlt2WOMupsz9bp85o1NDxXdRYf8nnAkeb1rbUzCU36la2tREpkiQfqm9xZI83mPj7U/m9
Q+p+W99yuZSVnOtTAKF3SoyNI0dUqylrKgKaWg24UYh5RBsloeryrp/yCuAuObo/7Fl2ixKyqUmS
IeSEfbNIEXjScrtkX9tQl/6ZKjjazAm3lljReOf6IkV9VBG/ftTQwLvuMe8jK1wntJpkcTB54xFC
alfdzqeJ7Qg1Kg9F5oWfNwaQ/xKyBoM+7NO4GnkdHe9jQrLyJFBvXN1W6jEU04QjdDuPCPS5oXDh
HwcbWUxnEgrRP06UY5O+C9p9fvqaLutHGqq9BirH4hGPhrf7X0HufOJnsfHiaF8FpiNPQRGfWGZf
vi7QAoV4wdyOGDOSOp6yKghyZIYigyIeEvc5/Ba/Mdj5mmBVFPv7Zq1Urr8wX8dIqxPMvxTRvLG+
/rEHodMMiiu3+ny5QiRmDSA40fqqYKhYhYEcLcdJBOKfrqgJjvBEizpnDx6ig0ZFalUmykFapa0f
uD3FDGxccGsBBYxZxmNmrpjOouBlhEtP1dSVyjk+/mRnksWYyBDysis2nHnankshHPCl/4GRBtjB
qgI4f9Bqg2HZuUE6VnB7C15N+iYhVU8CyoPwGxWoPbo3DUgoFbJhYG579nU6aTyZwZ0qFsdHUbx0
7IUhcCzevuFlDurMK8VXfRlK3GQXPsO1RpDWSKC1TvkOSxOF4n+t+oj9oQV2PLI2qS7eU8xVtoto
+46sSfJjs+Auy0tfihcKx3mtQDLBIJ1UoLUHqZ5pwQnnb0YcM3AythxagsQZ2GFLpR08aIsEzbkO
LOcm9sFRXskeYWSCyGGJLtYMUy2e5G1W0SvHBusH9hrn/74rF72v3p9bdA0EhDk0Jgd2KBWs9zJP
WETZp0url4y2qHGXISOAs8TLlpIamwtHQufe0Oj2aNcsWrMn/FgBNIHolctXXKQyXglqCl8t4vGt
DQvOXlOxYiZ7ZBwsZXYB7Qitw9q0OpPLY3MnyJ8RfpSTHRm2YqphdQ1QATFwWQxmHbUA5rqFkjH1
21uCYDreaPrzSXmGwFdfholpMHvFUH1BdFCyRf+iTp85PhNIw5HtqUUbtrEhdzJjuTjwgcu2IygU
Z7c457sKmWumI3KOBW25GBvPx5r1TsoPNOWK79VpNxJhfRAB7q4+Qu69jLOFFlA2pDgvrhtUOsxw
SnDQMlRASjNNAaG51S8SUK+lDx4aiVXFyxS8NOx3ckeu5Ww4UG3aIqta1RIS6+gmTjaJ9wQH6ka6
eV4kcl/fJXJVj8zWkxVJRCoxVTI0mDr917TqDLGUtPLssHuTaTT0V+JMdny6i3E4rDg3O6I4QnGf
9jGSOMP7o4ETuq7Hdz/Vo1x6k7snkN225F7ceb4jv7e1H4WpnSYz/FTT+qbRqLLh5ROezN126VEP
NnU8XfdU2NYYiJ01cSmG9c58PNVPxOIkhqm/ZBJHY2QrBA+LxqC5oNwm7Z4yTGaW3lk+wNPhAMYI
C9QvMEkxqB9+N9TIHUq3rDrKlbXGCs2DTC4CXQb9XQO0s21vAJip+a0/DboXi/J0/uKikQWWlP6n
K5PWzcML2O/p0covdXc3IrF+BicCPGGdxchF2ViK5efPUTw0hJJ0j3060YgnM3sN4dFAn6iv5Sz/
S89tN7cAg+/LJtC0kjJ6tegZmEb4he6T9KN4UN13VrejxdsejWSjAcS7QyW+AZlrMxuJsk+9GHYO
Ivu7cB/YVHBuYZxKA1cJSQQXQh32YdBPr53UCAY2vhVJ+p8onsW9ugnJsLpQgCG3ygukTnifvgrO
ow2EDFc/7lkHJBFEiUznNpumof6SRabmJpRg0I9axNfSxHdnLem3mhQC1BTWN2avbr0emOP5n0JK
2r/eavtUsG1/8HgBwgpSwnvzBIQqXpGuiIRSs2fQWWO/HA5i0Oin/HQEbr3lmsl9Eec4Z/F3RJOk
reFrRomMhWFHyp7/n+5/fPfPVpRguTdcdiEYdQmxc3xEF63ddJKTpSwR7nFes7+yOsYpygQlrN6T
ZhEVChnBwmEDhB1+RWXUp6MosEGQryjs/Sz0ddh7lA117M6n17D29vCsOfiKzge+XPJaW7pqCP59
iln02dkuOiL3VyTfLcHQjemJ5E8A2ZTN4p+j92IF9sbXYokpMc/Wvjhw6zZRwklv/lX4q7vKdBan
zj/8/1GuZe9vwCCWPHfcD9DnHBlzpCPFYcEpkwtY7XGer9IvfsJYK8LW/EobK15LFBK3Bd7kAiCj
FkR6aiUJo92rQGbhkpwM/9rKzKZatSsWU/7jcziq8pzYckUadqfzrbBxzCafhf/+3CQ2SulY+vdu
7tee0F+vfRbemXjDlhRA2twO+UBjQxEnj53nviyAUbOgr5pPPlpx+2f5iK00Lwi0ee0+nt+v/Nlr
jI8VxQ+C5WCpuraMQzaC1PJhTFiwWpXVCRe6ZXAqYmeOz1IoOLdqAbwkxjb2dk8tawJeP5Y0emey
OtAMsCV+rz+GGpuLXCAwMJtiKxZnBRq+slOTdEFR3K7GgS9BrwJJed8XQfAbs/hU8h4RuEz6riNQ
FtD3FIkev27GX/UhfadESO9PajdP6+AnGXZyxuuf2pdCx366ZHQbM2G3SMK4YmWM9W8UBcRzxiF6
Ac0R+pIGDTClYXeavGbKat3nza/hqNEYYcB+KYFARSVVUx/UIDyvK04xW/0MzglzLwIrwn/9l1gG
AAgWfYa/CZ4SvnIeooYrjyJpa6/NmZGNGlP8H2Bi4DBdsYUwgl2eaR/WDPqK9H2EkI1IOAoRC+Rf
dXHj2BUMcF/lG1CUiEPCVmyDCuOzkHQ25NwPRn/Q8rHuruvJxaxKTgqbalYWkjDVNzA5LS37rE0w
vEt8Xxd9hnSl0bXOkTPy+njELr9xo0qNYsGeThUrD9DdIf65r4bjNAirqF7WuJ+tJ3oX+8ml2dtV
C2P9YaT7iIA8CyCMtgwdSvMzwxVEWlDYqEKCZsc1FLhrj7RSvFSYBhjJJx27Quw38uiBmLc1lz1T
tn4aOTnwvvR4ytJEd1lE14LxQotK6Dk0VJBeKHN2waalQyMJ4G2xJ2aqAQb9ckrCJIy2SdUbkwbw
ARcg2E3oCuEnECLPZ6JrsPBkkKzVhwEWB3FLa2j/uwu88HoTmpML6n25kxItbexsxUPDoe6GvUEl
UBt4p6JDvV4OnJ3npM1vyPJlQBrzUWHC6lIdn1RiLDtv/1vCLQ0yj7Uvp0IT1z8NmfEl2mn7dbhN
MnW4LdUp3p90jBZSnDccrQ3P/MM+3/BrJGSln5Q0zLdyASoAV662EflUQ8VBClo04u6LNt1FssMW
r5l4a4pKIWi/OrjxpUC6Lx/j455SVgFXriwuq42YnFS+RotsmEAHKh6LIWPGKtrLDrMyDIw2NW+u
QIr6hLWhwI0Smv3iM+H5kfj3eYXbVUhhYq9bkbwoDtRXcBsB3zBw1MFjF8P8JmNRn5d88K5+jlid
NiQJmQdq2Zhg4XsuY+FbndwbLtmWX8Y4Bto/nPWQl7DhTavJBQd+AnULTCRYrP92kpmtSyxwnfgV
gEQsxQAHk2QWigoEYOnKWWgy2XDXNucUTOXca/XT4sGZjWPy5+R9sV7ytpiUgqDbIwC2srNHOMuu
geiNMdcFm2yqexrMmgW67Chq761rKRYY+j5NbgozLWlblKy/xaCL46b0WtOWjAfZiv7Sarbgj8au
0FHrpQtnrir9D5Q8exwDW7ecX8gLHaIjytQEShbLmQ9rbKcU6iIuFKJR/y2cFlPzDgScb9WED2X8
W6ZccHMT/zR7OEKLkAADVJwDm6GyCnI3wiJaUtnBdcwt1YWKRhX5ssycaPH0XbcYccqemwww1pku
GkVXmdKZDbzwL6gY0D+W7dOFKuMvglJuRjoOLIX6oh9Po6T6RwxGn5tOo8kUoEGV4KdZn/olIdhw
o7YI09KrLHT68FqVo476kr7DJV5JP/QP9aPReL1kakVllQcZyRAVxPpCXT4b4VSY5szIa/cLp8s8
sGxeeUFSQo4xv43hMtGnIDsI6PP2KUsmIUdbfxMiBcb50trel1r8uZ2QtTEdputpkWzpGGA0D1fF
AZDShdp/8uV+CtHT9TdJvuJn5KmK0kbJRBOd5bOCclz4Ca/KL1uIsB0a+T8du9kbSsF8pZBML+uI
FYfoqnZgjr/vi5S/6XHZMNIOoHUxiLt0/YHy/SjVvJlZZY2kf/sfrPT5One+7q+QGLnSWmnAiBR5
8vDZze4JeBefa2755myhUhFr/cFhcAlGEk2rNfVIKmK1/kN/2Nkgr6ukqrxoy/8OC76uIEz0ZOLH
GMaPnNUdvEgOmPlMgYneZK2d73TvrpGsgbJ2xvI7f/DfCeWqLGMklNfWGs0eSB7D7oTGBd7jCoEp
D1zz+iphpHevjWa2I0Bqs/BGjdMT+E7VqXDo2YyRdEV8iRuG39yWPQmNFzaBFYQXSE/l0EHwMI6r
0K1wvm8oM/OKjaJ0yahuLvHUb4K11yCp0h8FnVoDnp4Bkb2rC+aNyMXSQRj0iF5e8uucsk8Y90Sa
RZ198EVZ2sq5fv494wKSwheLBlpb3N8/+jZIdDR5GcpLpkAL14Zy45z4UgbzdCN0KhInv0O/qlxw
EVpnwWi0+LAzpLNn7t4ID4XjEt0QuSmGt8DSOGzbfbf5yEYcvooLkWhRZ/r6loN1hsKMlssgmkXr
XN7ojsDe3Hbh/wc8qD0O3zC6f6i7M96Nl5viM69h3MFDeV8jVyboPosttVPuIQ/ECS4Drx4Sgw6o
yVZRmPDrN6Tb21Y47U7wCm12s5TbNHOlkD8ytEDGK+bNz6B38aqOjPv/+U79a+xXXBH344LtdGRo
kpf8ONoWnpVwQqY6JzrgG1YT0NfFPC2s6G6WfitIUNgJfcehA6kfAghheYMwGObVw0ofEDuKeX+T
cdWtLsuSLV/b426bBCPmIeQW2SaeK/XINYyca375EY5a6nB1+mKLlSE/YkvIe3RNYrNJoPYA5QgB
3ZV7cwx/PYjT+NUeRP8IgxCour8xx2T1NnQ/RyPi7ll6ez/5JQE0uqHoNpKVNdCk7PJxcNr4T8Vu
txzkFo1CXDN9Gv2mRgwkQlGg3nR6bcgAP5kFEwTRf+5lz+C87ZD+U2IDLSbIVVz9Ngx3X3BMiaKX
nMh1IBlVItR7aX+hm3eI47cw1wD+6YVfHxCFWVwvdlzgkHb5rX/ulNx/RwWjUJsp49TTKWXLm9sl
wTL7D3Ws/fQJ2H5L17K4m7b2wqXFdgOH8VWrqmYEgM9nfDsIr/Nefv6Gq6MaqjBk8nA6U/O2a3v5
cx+2vpjP/gw1TYMSflgydQbm/WYuQ3Y2IIjOwOlR66EVGnewNBj3xH8pJSEjDSW3TUkLdSY4NoTL
asnnqDVzd9RkQmI+J/lQcYJjx6DorntTc8sc28I/yFYq/k91MZ/hzSAlJyoilOIdoeuILbBFT4k3
cqjaJAN5qJisUGGH2w6elyC6em7dh9nNL+2cGr5z3W6dMYw++30dqtOHR50bhPW0WVxTI9AvllUg
yqP5ollhsleVSfKW9CDyCZtKCmmJ18BdtJNkEEJQOnvPwPVda3dUGoRI+P567CjEK/ljHkWyc5P8
zZ98Xzpu3TLO7Hr29dVHRAZW9hdw2gVXjSz0kR7eTxP/r5e8HNvK0+I9WCd6KckWh07M4k4cnsot
cTxq+lckEyhmq645d6KHK2RvIFb/2t5havGDzll4dZOFKyJ4W9podeuTd749FWsyXJRvTEBz1KiP
SqQjml0cpxYNWJL9F8C2tFwtP33Ja63YIeQfPoNYWqmamU0fbk/YAEGlltvdqj5RMeksChUv9b+Q
Sg2x8BjsEKtlhg+GN9FTxD8Fc3GwLh27LY7zDXJLbVbO97gml8iGtwz75o1RMGCWGvWkk/Ogq2qA
gkJinaSmAMTV1duokZSs8ShB8a4h80nLf0Stpm102wERwxwVBEQtcgL1WiyLgtaXkFIGD5TyvtAh
v3JCltvq3+aZWmLW3mz4BKlP43TbxzTNyuBfQOwqTOpXvvbLEsJ3MDWyZ7BFDs29LEz77coZyQdB
zElClVhtK3O0f6unZfh27HQYeM04mJZQEechfJYcO+5KPZGKrmwjFdavF+FHxfVTB9b4BAtJqU5r
cao9JsrpM3TgBSsDao2EBq1QdGBXCnvbEViioCyojhGlpYh8J1jopNG5sZ50N6FewbxPfyxRei/j
bPRhfI7IS2YU7RURow/Epw0f88MFyMfl+WMzG6cy6B60NfwO1OewyFoym3+Nud43z1z5FmHGjAGT
b5W4c3fzibTy81WkoCho215ivhFiL7L7WCH72uMsT4yEdnmv+Cp7HnfsCuMXf7NKNYBFY/8teDDp
+rWQ4HNiANUykCv+8rDtLlwhpqd7yN+DgD7bgSjLgupdvp3pvy/0XTsQ4NLEgRBXwAWUn1nbn8hD
TZunSrnTglyvYyzSd4oeoyfMshfsZHRrmXY80gybnfhjzPD6DZTTYbqVCb1kIePKNRY0YENWOBM7
0UvQyK51myby2zg1ghgdQ0c+Kpii/okerGMwL3Bo8dj0MciCik7BSnfFoQlCkQH4WPeKmSuZGrAr
Z44TFTOuoihNGYo3Wne+hiGU4cE4Aomh2iX0PVwIvDyN8fygEWQLaX4LuclKaZREH1NNPNHRUjhH
/HyIdBO+nXzvjT5gvv6EGyW+Bz45Q7oTXiq5gaHJE5lH6o5A9GIyx0EUlpr1GWwne92WFjmTScDb
NAH6D+/7Fl3PUkxKkQ1ep3VwFBYzHRH4xmskcNl/SFMbQH8lSWMLd+HS/hNw6A9ZhTwOspfP9wKn
TewrDbE6v02U+r2Y5G++X1LnlzknG6JbcBfpb/q1OoKTrrGmerQPRao17KYzK7VAm1ouCAcxjHWL
UOTpy5ZktU1bwhnmb0K8waHNZQlfqvJ1AxZG9M8QccBYilmMEAkWP+oE7+GN3EJCwLfI5xM4RaZO
MP/sbXTlfn/PHbzU1vpinUUyAQQbIR542AYTLo2SbJrPtkPxdMZ8isK/OkLcNj2FjLu/dVYnzgHY
Vv0M7NRBwmfuYychyRxOygjwToTvDS6/ln0NpGn2Hf02p+ewnQDJ0bcMFgjdLrwRfJWok9QSi2zo
D4uLC3RZpCxH6xDcrSlJlIUdos/6D3+DGe1B29mYah9868q+jSw7VmPeuh1Nu/CAOu6VDDX6v3Vz
RTdc9cvh4Yjdd/coi5mlS76SmrmIiQad9FKb1TkcLHwxkHuiA0VSOYvKeN5N4KOIw8auzDr7Un3C
Vn9AKjr5F2PoD0vp9iiPmGHvaOv4d0bk1Lq2prfnNHrTj7Rz82ZLVwpsYAcgoeXAWMA6cSc5itNb
YHy1cqciHcjDCgrgFyEqKzZ6TMHQ9AReurCuDwn01BqshAkf7CJU8dYd3nRd4P0G4GqrPD5AOV8j
M/FgamzTY14s4YUPQ+BrcTvbP6ZjhMj9o3mw/kpceLAtiqJ4PGgl7RIXp2ad1ALu8jicoivcbTtC
WNSlmzd3maJdU65R6zqT5JC2oElWhlS0sq9aqXy6ZKqfnguW43Y6wumf5KM924RR5NX5/Qe5z/R6
+vKx3tGIOxFnU5y6Ez3NbBsoXrQiaTlsJLp5aYJy/Vr1oMyMiODimifZmudCt3TizTLMPzAUGwQ/
2FszGMSiNaSiGudYKlcm3w1BRbq/IW27fddao/ZVsAnhbENsqDx8hNf99XH6U4U8V7KPTlZkQE54
O5kwewg2A86V8ESBCTMcmzH7aZ5q3sJKZnOsTLdppouaHJAjwLAWpvoh1t3TU3N44XKtxygyAk76
yFdx+c3byDlggOXOGp2hImd8izUJceo9NtHd3b8FIzxwpwl8vFRAH3rf627ZAI5rJFl5ZSY+PQBU
oZAjkc7ni7WLLfzAc++13wK4VhYMmJDaDThI+S27yMKKY0dBQppe7daigQ9UJTK0BrBI43XJm9GV
g1o5xg5eVYEndcDOzV0pgW0fkj+8f0oLlwX7/belRTugjz/EgMLi0oVChQbz+my2+eBnYQO5zvUo
qXquXhiBu5U1ReIOcakUocogKILr+Gn5UU1/iEAEgiqBKx01D5f538QnnFaCBjmtTgbU87uR7bRE
jSooy0FBOl0rbrypuTjRsPXXHwWxPBW8IFiJxE2AZRIef6E415hXJ01HBzM0w9Silwic3WXVtVE3
284bmp92iimdE6IKEWQtK+O79fYcUINPvIjWQSXxIVDKyytqQwE4P63XziS6hjezIbwVgAjuebvv
0v2fH5xYxRioXm/INCK7xg8N2pcIPEd997Pih+JQ7JPwSPX+K9izjOXFrPOzLMzOzH5Cc+wDf7pA
UtwcJA8h44fQsXsip3m02k5ecaHJoqpJ1GMdkWuttM5V9+13aq40R1bkZyxkll1zotEwg2Ac3ecs
PWis3hzR5N+Tm1ApvulDlnywZ3VgLtvmHPsmU4uyKsiq7F5XR9EymzxxIcQ/uoJcIp1DJh1YFlwP
GnRu3CCYZj7wVas5zkEYZbOIIKkqWMM061crVsK9S1spCCo1CavGpmNnff4N8pxO39qrCD/L+aId
ItL7gDNiK4EkUAZkRzgrOP4omp03b9JL+VLqBVYHlhuX3XkwX+94dhAcJRXPmakYXu0lUaAMcLvj
UvAsF2W6Fn5plLcxnpgC7V3G+G3QpOzvg90f7RAULGO88b5gUHW44CwzceJbXAxmlPhqMVFvwg4+
baFSt2VBJSpuRzL8rIBJWXF2nZOB3o0DRf8uPnO0jO4MYLnYJeqIjj6DJ+dk/gW6AmzGvA4L6Z1G
1gBFtci8eiM+b3Ku1feN1rQn09ljeFezrtIqfjLxbZvQWC7nOBfHng9BkFJekhLiNwpX7A6DvlVy
2B0bXvzP9yt31fLkYHrDkAIzyVU7G4vYPwkZdSQ8adPg2XqDJNX5l87eKTePCVrjnHNdex4NOZEJ
ny4BjF5HXNZs4K+Z5zNe13Ib9hI/e5QLMnxlyJRf9mCtfHUL2a4q5YvkEQDd7KgSdkg6zJroOrVl
Jjt7Ws2qTCHDjIc8uPzF5gZ1o7Fp2bUqEjw1zL3GuZ+YXbpbCRaEcDxDg03oEErmsKTEtUdntzGH
0vkeVG7fO/CouWagboaaDab+i5T0nCZUIPtHKPlBKLzfQIBPo61g3xhEHgcI+yzuU+VbXYj9E9pu
7zVEm1VsglLL+6RoBfMQ2ms3JFkdxIV02VV4MVhxABGg9UurWFh+I3Sdu56K8Yt2s4mbmCHwp6dR
b1h6ZNz5CTtOiXNnepRpHPaWACzUKNlZwTLycn8X/pglzz/UKmqoNcwQZ9xbdgW4K3xEofNaTO9N
oDc4MBOUB7D+ZGmOXWqNPX9d9A1jwcv5uT72Wv0JitZ4YrhOozudG+fDm7RpxeNfNDOYrSU9dF6u
MDnsMYhoragJoFqxWTQCRLVp99jzUiDfRdD7W8we3lNEJ/riNwPKRRRnUXaAeM0Z/5S3nFglVG1L
ifPS5TEhAPhAEOlVowOvwPm2W/biIh1SmJHbKTIFgA2byyprATCQ7j7ZV6xhggI2BeIjF3TueGMJ
fd1YbMC28IcULZUByAyGdiDFuvXaeNC1+/SBbjgqIM6dGqBqkLVGRBtipb5AjiOb/j93+CxE6aSb
3HtRaIju2SJgxY3Bwe8GGX87JfSq/iFZ6dNRjexcQyJdZSSjbHubCSz7r/iTD5qVI8wtidHALC1Q
GHA2EZADpxIuGWpvpfL+kVWrkdh3SXR0YXqv6mtWAIHvIc7q5bzWsRQQaeKSwhUKorvJSnUVUh13
awzRKAgnGb60/83FFWJFrIb6eWjidaoA83cwa/oTsmMIlW9h9CN/02jbqeL3HQor6+nGok9Ss0UE
45st8GSa7CxYPO/lFJm3vqe1GqKVmWDDlmXHpW5y1TDYojVIRN8OZUUeLtoL6ZZMT7IvCpiCZacB
XfuTmdC9ppmMKOlGtNTUvkbXvSLf2UNETN0eAkc86ZJTh3IlHrnPAf9KNAL8owjI+r9vYmXNn2F/
gxyCfK0i7yqHhz/XHzMnUkpoOoGEciyqrX0FaVLjiy3NP5zoxTjpmjht0T8CafRKXmHK4SUqkWnN
Dt2lxLjf7GA57nZHzmeknrI1VeBlBF1A46SS53YoxBRknh8FAXFZxD421j99Bp5SgbdvifAn1ICz
Y2pTdScKgNXRF/dzNQ01MAimJSQeghjFpQAOenulwnfykT+r0S6pbrGgIbe8qtSFBUt5twkHBama
NG8mnVts7ED3OZk2CTf07CiM0dUmaAM0r9Xk1tINVAy5QLEMGjvT1Zn3CtZuPdvKyeZdLuaqf+D7
iovSEM8ByPuT1K96/2jBvJd6GmIAkh/ReYKD0VIX2ufQK/Fax83GeQVY7F7HRp8sj/o8qjEY1UY8
ZeUNGAi1OXOCPjODiPAYtmPUL70xSnPrvVTWMQB+imtgFW0rC7Yg4mcRWjFWCCO0ltOvombuJoqE
OCFnWEblYpj17KJpIuP29bdKBlULmmi44wD6zk8PVW/9kyXH7xCBOqbuRy+rWAsXTeWTqpvG7sUA
EcDXb9GTQT4u2PXOqPJ/hcJFSKGjijfJRHlosnqe4srjYA9zPkpzKnF1AC4VcJYbx6kVaa0g9VXO
srnR5r7OLbdCPvKXejbcDobO9qvWI2ZPrC9J32rw+sNns9vdQ1V5TO1pj15BtwqulTq5HY3uj8m1
TJp0vhkCvD2q6MU3IrwaDPsSPX+o4oX/nF9BbI2QFyZbOHjsdRqF1myiA29pg+ad7Ze27wKcoaeP
1NiLHChY8Lbvlc+5gsCRtP1Mrifelm0AvT4jzbFODFugJ25aMtbeGXuQwu0CxMFSZkvyq77mFwL5
PWEbOFQ5SujqqsQWQ0Yq2F2TXLpGAtt94mCXAqmDyDiq5rCujwRtC73qdfMFoEbYV2zOo9hkt5vU
cVBSYyc2eh8+TbsAwrtdki/QdV2406VZF6219HWv1bLIWCnYmTIDKLBXoVqevzDPzC0NP2pl5QhL
BJd3DPnMUdkvqCPVEghpwwOmo71uIuL7xfmV9yQbUPvU2O2rt293Mek4dr71BOznAnQ7KiZz5KMq
yaibnz3Aoyg8PKHt/No3C1WmyCVA3t3yZyEWnZ6e9XMOArS71GFcN8Ys5KpUjWCC48C7A+LfZtoT
oHP3ZV2Gg5ZMtx+Xt47Y27d0L6e8p/Axy4CBvHAHJU6yB7ofUvaaU96od4NW98OJIrbd0BOxQ94S
+C4b24Z0PaQY/3JrXLTAUEgwVLQNXcbsGBrSycH6cJzOcCE97VqpJcN8h+rDwwWUZnzX/PiVo86A
ubcQHb5/qbQ/nqmy/SOKN7ocGJVaRnEz3HI+A68AY/qFPeahpboVmj89ggQTUvuhm927lirWoSIS
55Tc9ZD6QvTj1oW0lEq+24ZYWX+2/zyYtXgUB2+Yng2i1K7wE92YZuoIx7AC+aOUP+OoiBQyZcOs
mrcA+m6qjK1HR8fYeA7q+EDsI3mY1tV95GKPDgeO2qRG8AYTMb/ideMxYKZdVdwC34ju5gHzAcSQ
B19C8fcTfNer4eFEJBVkML3sfQk+/7k+znnB2bNJs4EEpLZIkcD8Dhd+4LryysWnOmWXn5avFVa0
9jeSalF3NJvhkGMcC+vmsn8LWrcguKTC9VZV9NH8Xysy1UWg2nEG3T+rh2On4ovc4Q0bjZ2zVIXe
avK73Wq/IV5biTu44AOW9QbVDimK6GDyWC7PV5S1kIolTzdw8Dicj8U4+0ishXAZdHsvH/jHE/dC
Tm8T3byQXq7xoFkJryWB3WcNQlAvBUJwF5FWdqEP8HkfoWP5lVxte0MklrAq7bOb1lUI/Lm1zCRc
q4t6c0+HbiYZMQ5QMkkK3ZfUAD0+ko6Hfq0dz1GfO1nSletLiaXlq/ulEhLU/Os6LsV+lwZu+U4p
Ky1Vprt+9JNmNr/+o8iBx0JpZ553zwLIwYvgHh6ScQxsmkbgfq4/bO/4xV0IV4IceNa6fW3IBHAk
U94S3odk2Gghz94FB7cI3w8o1JeDKd+cXmGTEQUShwdZSWGUqcBKjIsSd1F6+9n0kn2Eoy3Qd3lU
p6y/CSw42NXcYxivcxef2ACt4xDWe/JgnLDkAFnh2z/VImakQIYgIUvhE9JC4423y9SdCxhkRo22
WpwpHTVcEm5ft7cpvN7Eftenc3SKEsJfJxpPcHSZihPHNiI34aUQ5Z2CCHFVjXhtmy9KVDtoFigB
De5OmPaTlCh+DE88vEl8DwATK4AKN3Kj2HqD/WJn6vFUUJGENFQwPHx4HgtB1L1ZXoBZcohH8poh
yItAbGQLhMWBa5sIq2loYAJ7NOv5UHf8jhN786pqUquxlWaV+WweWPd4sPYBZ2gFnEx8+VNIJ6Cq
8bume20AVSeFvJ7BOJZ2TGipp+CygQa4TiCz5Q9xkynabeu5MkqKJWldKR188wchmuHL4LE6QDci
egGgD30CH6xaJAQcVojkaw4wiyJsz/RrSffXcCYZLIyLjJgSeZpd+7qbzErgHZMLb1ly2+f+Mvuu
betzOxzP7cn6YSomShOsclgXLOKF54TX1EIlQRbJC1+xTgcrQitZyG+OXVGwSiNzr0QnF2CzpUC4
1ONbBxQxofhzncTpjB/gcbWDuyHvFvXW9aD2Sf56SDtxIp1aVZ0YwhY7XLFLeAed+DUanfZKfAvk
KFTHwm/XzwmVxs4mwhzdk2oXdK8MHGtxb4JdZxfs77msfLRl1kqf69K5gO3jOA6Rz7ZES4bSzB2Y
GnQFREvqz4XAwxvA7ASGkSiQiozJ2GtXUENlJpCoHpfHJi3SCX+3EVklh7IbazX38PXIv7E5NeZ9
9NeE4XGf+lZgQ8MYuEe1XZsjVFx8z4KF3zyDveiTF4LGlThC/UnJtQxxJ7GuDMT6TUt/yDYigJtH
RK360gq5lm3f+fcZdXvHHTu+rwV1Gp/85L+hAtMs9q6LNW//y7zE2Oixrw+FZ0YGuHFz38KeIr4o
1zrlcF2TxCNEt55Dht8PVgAGNZUBHLNFPnTcIrirZD5jitG5AFbQzU/fvHm7bdawxz2LHb+p+TKA
F0sxHvV+j3HCK8TYaVu/3wyojbPUT6dY7Qyrn8tCSR61/w9IHhBxIKYELTYwm6vJm5+Wwiy3TLP+
zXicfEETvraWIMlOp6XZ6ICWy8Y1fUtVYeoNQeEGiSPyAEc7KhxyC7LBBb0KWwBdlka3g9+fbrAP
ev47ZhnYDeVWIv9QDtg93V55rcq45AYEjhn8bFr8En9e676zZ0H0u+aX2Lb32q4b3kd8R8p4CcTr
iCf4fIynNq94SNYkJQ257BqZzsUH7Ej0MlYmda6XiyDZfTR5b8BL7dkDOVl/omT3HiI/0yPdzpmr
djnMmhvcDInUJdwCQJFEjZ8Nkir0qaNlOTRoZzFumpJFNy9k8CBk9eQgguwtE1kq3BuMCtq1n08K
KiKOU8QqoVQ1WluRzoJ/N7eB6ccZfTXE4LuNIBKlaDul007V/4xTiur/TcTah06EKFkfdCViUCjd
z26vstIJZ2ghJMMSwVnAPC5cEl8LcG8AUvM9cepioHv0I7Wqic3zJMksG6byVWoAH9sFlzQYKE/e
UKiVmK/idUd4VNjbEGDoof/3BeYVb5bo9L7BJcwFiv6IRyrxeIOiFYc3F1fS2PrenOaOqsMSFNdf
VQkBfFwbYtSysiHIBvt4xaP3FgXHp4LXPXVAAB5GRqIcYAtR3aEWpSAqpRcoAmmgA/GJ3YJSYt+K
NrW8Wt3XdOo93fWlriS70gjlrYGGUOP52mlZ2RhDmnvvdRQ/8a+n0Kg19xh6QjnnmS+1wQXt3nqC
tE3nR8aPmXRlAwcxG3beqxcNHJVPMhQgEugeMBYoYIOaQsiSX6JaUHD4/Yi/ZoFhb7K9Q2elusIP
bQQ0X9zoDUzxdWqDVnDRmtUXxfuwoHIGat39mZ/8AqQ68BzAo1atnz8xM0o2K1JShuz3KA9/LNiP
TRLcun1VBcSJ0b7t3DRx2z5y1AOTfl9Qdxha4Hm4olWMUxhlgLXnzfdQOuy7hAF0o+APkwRwYxPJ
rQQElBMPxr7S8oQPIPrDWhLuQy4YVpnsdau8SAwT14p8BaP5ZMIwHf9/DVabSdQbQymmdCTf6MCQ
kU0DlvWCdUAlGxxbGNojjmEGzvzNhKYrlvKYXapIHLR21wRM9tfY+tU3QVFdN+GJrOHZE6cTx3OS
PlZAM9j3uqleKz/rmy611oMYC9C/o5EuIv5KajH8y2ZbO3EJBFSDey1VpoWEI/Q32eGyQTKilD0s
2ulOUGORCbVC1j3uJ1eoFANoV9NcC+KPBvinjdrUGedb1vya3s5XJAlvjs9/rnTttr/Y9IlzK565
TOdoyLflkmP6iAAoHgx9pp15eKNhFrLN0ObiIRGcKGl2ywe+yDzTOex2t/RrZX1PCQyTSESAIdt0
qrf8fVdZmfSfBso/Fi7FXYesFfejXOOViE4/bnlkiBSdp4vYzxx3xlIawD4Jvw882H7f6nYm9rU9
W1db0oUu5/38cM/HPPEDV2UlewP2LZonfG4TXwoHvf7Yicx2dGvPw6Ssj5ffrh1sD71IfKSWWwTJ
7Va1Uek9NtMdCxKiANOiamAcvWx8xLCoQf59kJyOTNclwRc/GdX4hl2YAOhU5ylPWLZ+fX3dUmBI
Z0DgUxmXyMFa4s3rnmOUZie/FB19dQaQHvjqyr1fACMncc52BDxvdynjW1jOlUKgGbOVpkeiiVnA
HVRX+5jAdY0DNUL3DVsLrS92WyJBzaSxXRqJJwAOLaJaHCaFyZzqqfjtOJ0li87rVdFadYBLYj4Y
8yxfdt2hF7+T8BcU5wPdzXFpAwBdD5vUxPDNn/ZMfF4qJQIV56bO1l1QJ9VWE0F0nRpSXXv818Yb
Qn2XYV+fdrXvrWEltevlsHK6MzRVLsT0Rb16XqFAAmy7MGSKzyRH7Y5ewsuBbE8ZSjOHh+/74fKI
7T/9pmMcesGEgTd03yPC3SMCHXl+ZVNfuTPub8OnEfy4EJvE0Sal84qpxY7PyFq59TTJ+OFDV0NM
1XIzCp9z7Zxun7GqSfoZ6oC7nx5lSwDPwLIru2sf5jrBGp01eYbOMFL9e0eLm4dCuZzcepG/j50O
TkHi23hn5WLbM+nvHs1NSZ06PkixgWMTOBFeEvqPXqwuFYIQQeTv9ESriZCgTM+fmwbOWA0KLI3X
ZHavpTL3CdfopGCpWjmSoXGFptEaBn1d46jvNQ9kTUfDgqb6xyRz5ayC3lJy9aZh0XN9vmIuV6Sb
Bb7k+QkGlSYPuFEeIdLt209/VD1qVA7l0lwi7ElPDTL9qlH6CCZ/Ztj1UjBR9MAiKNj1W3/eyyDr
C03I4c8EsGELyxB2inE1Tj16ffwJGsRrU5Sj5EjqkkXOZAfRKY6HhtNeH3yohm15UTQhnHa/nNyE
OTgN4F4tdHFkeK6m5ltRFpUpHuHKHYVMTcxUUMsf4COzMYE4e2mcZaAC86A+foR0qd42k7r6fIYm
vX5T7yQQWxjHOLW+EXCmgm0td7mixYj2Bxftd4ssgfPXdlSMrHX+T518/knRUDC7Zl8O5DalkYkv
MSJ3QSrKqXXhrMRSQQofhk9DODofUJMqizmNnv9wis/7eEL93YBlwF+BKouI40IQE/7VOKmewHjn
/lRAr5klhvfve4TX2HxugaAL16tXeCShlzbpvekwLZHtKrSMy28U5Zvbl75o37bzlFdfC/dg++I4
1l7RF4f1nbFs/XjK7YS513lgbRLwzhDHzC9XAPyaPJC2xo9WzEG6phBF2MiutHZ3uTXgr0PmHz7y
vQ5Jk/sQNqMXbDEtqVgV52YMyyUbc1KqFewo8vCKaX0nsdRwq6YKvpx1w/INztQLV2CveydSMJFU
Q/xfVRWFCYgI/ZRxiQcn9pcDvr0c4ZJgLw6m/Z0OWAuVQlm2jGvEWqU9IAA0slbWH4oidTEhcv8w
pNDY4Nx3NoE7nstZKxHBhJ8lJtKYdbr/L3EQIc8xoORODbltSp3cSK78Ceb2P62rar72hzVlXJur
cqiFibiyZav//RLVfnzkpz9HyjZKs792qHcqsCUf69W7x+sbKKutdpIHC5NZ913S9QgtVYg8JHg7
agcdiTkMGuKosQqRxEJBi3YbgOK3fQ4sqfzeOhthTHrgkQKwIk+cHVRXSY5ZPaloFLm3oPa3hn9Y
7U/TfQt0rrnuufBUQVtryYTsTNPT/M4YgR8hxcKfXokn9CgBCtXllni4kloqgh5INcu/XsXSFHor
7fQ+Y2O3IJGp2Y8TfwDZYrfGJ83Yj9En7UwEoRJLDgZDs1zYoIt8NIZ5gJUlgelcXBmb1b/1fvsr
f2lmyPgySdNv8xL9mHN1LLm/fyPNbBnNb1nlb75iwL0/Lh05aOgmFn0wahyrrbqCmWyyfduetliG
YrzAaIS/G+eV0ofCd7fZ48U1Dc5Px/xeBZnTUK75fLk/33kzh+SwB5xz0d+HrLaNOoie53IWEqb0
sJ7giry4wZnnR7ZTWWP2rHwjqHB8RS1iVA9kAe919WuID0VSuRiW7joykN1OZZE1fLj0B0lZ/wle
ecoqCuRDqTAiSE6eWIz7dtmvaLKhBgI5mzSti81Vece/u1Pz1Y5IDRFrAsSJvF94VIgwObC3s/Bs
Xpm21+6jQoE0/IiT7MHIQ71i0BTkxaemWXYYcuxHKCu+7nBCiUxek9AmlSuMFuApt5UJTl+amBIn
WXYc5AjyhZVfiHPLqYDQbidfVmOjEM7iAOYC4u6dZJRWxmWHRyDwMHDH60PO4EelU9IbtlM2wzcV
NFQlRTD/xLP0iV1Cwd2MS23FPRdFq7Xrx1CwRTrH3z77eJnUmsqwKAyVUg9KKJHXLg0IzSDSFZrc
jOQRt/0/kZshKnMG4NDN9iDZAztDe+h20oVqV2LpTwwEunrp65A3fgAAmOY1/tF3iURQpfk1xx4Y
At8vplCup6j6PKGNSn9yvpNyndd8m9QYyBVk2/1DI0rYE6jTsOczGo+yygzQ1w2IPjVlLG+j5stg
xdm33bLStMTmJvrGEqb3tJvuMX1BqhcSbswDmRqy8ciFAZIg+1I6ikFrSe4Esty77HtMGCKt0+oo
sy7UzLCvAVS3OYDHAqTFdQstCAMxM5oapCQZa/WWSkAGeCvxLaXEXwJ7cWu+WcbZC7cENmflYWMi
rHmjdZvl7poW+uBlMzsT1Tle4QnH0KALYZlAHwmQCAVw9hj/na/TJNWbIioKdInmahin2pa3MK9S
wtQppbOzYIsLhZ3rJLQTOs63QaKwP6Y1ab1YtgAlC9fpLIVTQ4Q2VSwrdBCJbY3L5CJJOSJjwdd2
CinQ5FxVK9Ma0NIZnNDfsYrrW0eX/T8W7OzmAJGm6G2tJFbjOrwey9M9C1NY4lvV0yyoPIxKhC2v
4E0mlqaUJeOYGw5b36NCjavXkjtQubwS4VMKbIP0SXwYJjFM5HSAlQi9f634wQKYpG4Slm8MqDCS
ehxPcenkcax9pefbhPplf42vpmgmTfhuaVcn9J6ZNKM0cG46Ap3JATqqMj7R9SDgsScwITgDxvKs
+i8Hnman+k3wHAnRSMunmU2CWNZm5sH76M77W1cQ2bfHWJ2ZqmpZHP4GygG9+sKvH0073l4Z+gU0
I3/OZHUaaxn0U4KCXE0RYRipx/tIwxOgZ2ymg6RwXTXREp4WbouonAV9Yc0mEneN4TcNGUR3Ps4f
b0wlPZq8ZO26nqnJTVqIVhjiLGQzj6GJ3+GK2Nr/BuODpJzxbvTNq1LYU7QP6j8vOm46ES+L7kCO
t/1Q03ll1y1Jyp8ggdS9wc6kFPZyOoDU3yNlf6gvs/9NT7wTX/W9JEef4FD4e8VxVfAKETg8ixvu
BPVmG6SZGWVQS4DZTmSiEUp1sc4DvgKCdMwQurt7FSslOyEvavPt+r6X+tWomTnnv0Bh6v6g3mEK
tKBk8HwnyoSZmljLucHEU1lLepQkYYJDV8LybMmoQ8qOhN6sdBev58apMM2jOPNEiS46nKvYozUw
zXgcRx2fi31hiuzopusLl+2mtB2h/0Lni5X3vt6x1k6Mv2PEQ0ZytSFjROSHWp71+O9whaAcXNtN
J3H4mNC0sw31Knvo+Y4lUMJH8bH6SKhgbjWIsqzWuspnqja5oxg+V6jHPB8kNOFVa/QCVWZulZBb
5bAK6KJTvMYWsYS4qdwMmBNolbT3CZ6KnwDl2CO5RI1FnMT3qNI2QhQlJnXvC56Vql/MIe3OMZOI
RJaJMf3TIHXmzlfIqXN/tqF6VTDPPnhkuLOqv8j48Wjs21E5SjIKwFYJkBrcuXRuR/25yAqv6BqE
4I9p8EP3qGcy38ziOQ0Qy9Sjr+nm4Q0xXHKGUEik753PpAEgt4mTu6uz5cWE5iXsMYTXH4TypZ1l
K466jMkhUWwqmH8WIVI95w51XdLxfuqYpWBYNK710kmL+ORalmgRmjRtP+F8AZLg/eijSQdtZi8i
LWONeRYKnKbHn2IC8e2g/zBeYlga91oDHcxiA6VETqT5e5WO6yJbrpi+4Q2a0ddYGYhCeZXTPSjo
8hxrUtIyoZkYw5XwUMaqTDs+jlQwoAJlye2QmZcCiAYgGml2fknUCpYanTn2jLkxkB2YFtASyOPN
mfNfiofR0zi3Pq7NuJcFGegiB47yacOI/wJ4l2Wodrlq/x32Atv3bXXFRfhJG0cVZ6TPikAv7PHC
ubAhNEGDod7WcGQUGSGKw7qfxJgx337oMaa4F3BvK3/1mn6YQ4XZ2jSccC3980XttgJZbhbTH6w8
kOEtBPZla539VRBFnp+MRKol42VROGYHIzx8SqRVaSzlUVQPNqX7gHVzuvKsS5dNVP6cNIHbVbTL
dUK+KVJiDQfeMi3iM8/mQpCetAgRjVTCY2qh3aFQJqnWU/05xxBktdbv1oHhPooAI+QlhX18ftK8
1RpZw/xwBaGyBXc0e9547K9fBf+8pU3RMa5fOErNCawfYvluHgV1LJ4FOWzm0qsnSFiT2kfBYiB4
uZx0dlG3VMvlKjQYqR+L0iEU+p2hxcm5fzv5u7/BB7RiWQUF3Qo0GZa2+EAl2rz5V6rMQp28xGDl
Wh3Iv185QkIHSSPh4GmD7IDWuB3IAnnPub1My2k4nt0Q1L5jCvY6YXu9G73ieAQOpgE7eI9jv9Ed
wnrfjdBUBo2xtm4I+2Mq2xu/N/It0TO6MC/D9z2bfAbc+DmHFKtCGxsHYY+fD1Al1IC5p4efF70V
q9/rguUnQSIEXPYFFM9wFbaXw/hff5vXlyrKJP3D5tJcz6Vs4UUY61kW1JMAtk6M2cCoQJYzCorr
DgNTigMMmitOXdiafbtAPM0Q73qpHLuaaVTt9hma8VvOSWdOu8UlWGqjaoz6NVUQ55MIgnCtC+dU
1DjriAaXKIIGoQ1BEdOyN6m/pV1J+odV97CPPYgU079npKv1PSRhMijcQ2xKfso+947bFFjjW3Pa
EKmPBGRsUN9O3yjTuIca123QfyFJQKQ5p0BRKfBqJ4yIuJSzXbWJ9P7YpBhWAK5ywyLSQm/XxnwS
Y3BbJGPYsIRn/NYBzEiyMEN3mWyoEutI/XoMkSfxDeJ+0gKIcS9rI+3s7X+rNVbArhihr2jfmFZ4
WunqYywdv0FOQnUuUTSwUCTg/01+q3xWSXGc224Ic1fW8YU+ccZoiwadMWhaDFWCUj/g2iKEb4mW
eE+wXxBRl00rtP4ZOYJctQZcE4frQGppGJ6duOy0xzYFaCS63IDAZAOb3BpTx4fJga9GRIr5uODQ
XdEiwA/qJS4NHHteAOfphqQGo7mUlqsfejRDtpyEAXAekKISgScnPM+rA4dWBDJJAFQohHEQopik
UjAtccr713VkpHN4ruLEkZTmQw2Lnhw/ps1XkL2Z0cGsHvYuNAwlYJQYLVMNje6tO9kBuvdvGpzc
d/mf8G5dZU/sx70vHSwt6dbL1vewmT6FM1ho5nPfYO+Z0W1YSc8r9A2vDENdiJbLHcLyJXgGOwv8
jytv2VZkVpMK8Cq5xSIILh93KiVegM1L144hCASto4JeuHSREPq0ULDP6/eISF1i/cwU+Oin06Ks
JzteGd4LTJt1puD/hJPsSFPRVnY7SHH2tdeNeXLaTYpNrkTDnIsivebWmKWE0cyHjzkR58x8f3gH
BVE3oiYvhS6tj4q0Qnc9tQM5B4M7mxqV9zRlD6tCiKxfx4SLY6C0vdg6zVK6Ap4bSKJZpuJeZZkz
Cd1YlhXnCJWIL/t0SCFTBHOLUgvo+z1tM2eFhaBwnsyg68Vnn0cX8FC8APcaqKWgKCOGxkmHxRLL
/V5KxEBfN59Ql5Hbcd/uSFGbZY7zJ8GzJBw6mntLQJJZaMdCU0zr/utYbPVA2fRTj6IBR5hT5yBc
AWSjKfCzpJats+rc60fMI35PYiAvUxEEKmM6vPqc7hH6YI3jO1Plo1JqiK9gqOWYG51Z4qvMWUiw
HeC13onKkEm5ntxXmS/6BMu9GSvryPHsHQyk/o4YE4ulMOjvbOPluSamBQ+puAzqhosXtlk60xMk
SUX86E+UjpUI+0/0fcsJ2uhwaRxfT21E0uCIcMVPNvXdyuqkRCIm2/CGEDqjb59V1h8LDRvN9x7F
FtXpRIuxxyhVKyOXw1YQvlZun/UBCsXjwG9Vdl2dLtE46T5tDnAWePUcXpQC/lHzJz3ZMxgmZZNY
wWpUke+ZJnOfFJqYhkAXukr2MkPk0mXZ825PXFe1ykQUl1dGD60sY2Avre0p0odNdRnpnEN6mFH3
LNACKlIbQ/gLXLxdqtD82YQJcg3c9j31RLk7MT2Oy6Xf4i9spWMO+JOKWeLdAOfcJJRwBOcZPlet
a7EK/do5174CyfaJt7wHIp6t8XtlqqsSFQjYKJeNq9EucGv/9WzP+p7FQsdRO+YJCWgH5uR7gGHa
8dIa+dIfYoS58Z4z1sEMLrO8PA9OV9Cw9DSZFFnehAdYeA/slIrCcCht0+NHR6o+MpqeqPffVVgl
BtMmIC3INDLtYCvuI7zSFKiuUD4Ouvm0C20cEX48CjGwFFjbfxQh8AgQjySqbnKP9/u7Ev1Q8Ve/
slRtBOmFr/qisUETbQ5fUjp95/jsiB7f93LdJgY4vs7tcq6M5DIZg5mSlC1v3qFLwdP109mcUURu
1hqknrnfr3P6b9BhafvynEy/Sw/vJW84LNvJEJ9xbwgwwGKU2wX87a0cuQkhgjMkM2Ahd5A/zUdl
+b+PJUglleXU3E7MPCe+8c7pGwSsNgfykz62HyZMySF7rJTWVtR2vQndvo6AZ5b74dRClxbOG61T
SYKzsruIK7WSZgVDSTST9F8X7RsWa3yJkApPhIq6QwskX4hIjM1DFAxUWTweBvofeNY86EK92XNQ
D0weFwUusYl69ng4ro/rYWDWQYW+Bk3zFXkPo8QKcSnQbJpOoNKdEvocq5jfQoTCXHQ8MNlRxHf3
4+70A4jWMYYcYQfzA/HV4+FRg+gHbt1I+MzeRvurqR9zx1SPlhllvfFGq5e/03rAXtnxa/65M+oE
H5L0J57x3d45DsWcscip+xbl6TUHoARvBK+jLqYA5pVfccMwmUi7X74n+3+MAJ0uXj14lSjtq7J+
q4C3BSRlb93N7Q+JO9Jw8QeurYHcqlHD3oSdQYCBvCqiWkGLRbMIq7XJX8Rw+YNUfvWv1LOgN8fT
4HyGSzACJlTz+5T83M8Ajwvf4AHMnXsqjX8Yfzuak2mdfIF+hae5xXrY3tSxUagth1MSVBXRq3qI
jQYwrIB+feAtwamfXQgSAnMYpcgooySdC8lAlUtRv7nE9/E11JNLpPUY0jnHSAy+K3ZMWGiEA6co
FM3Daux0xO94iUxM/dAalSezypQO0+TTQQn7Nvp0+I3EPgf07McN07gExqSAQOhAXX9qr2DbMPxZ
2WWWAb5kkkF7m5Kg/TmKuYKZZZxmgnjHpeo9LFL9rRmSs5H+n+PDzjPKI+nYD9aghKe9N9a7jwT3
q9T0IWnepurbr8fmQAczOVXKCl2aI7l+s/eSc231DbS4NHAWS9CHD8SyTcFRXtCS87Oj+/26iTOE
e9oVXcxbTgLLB00Qk1bzhXt83IW41sqZN2ghxKfRXpkC3FWv75F4UpruuRqDT5kwkhwp6EJNg/TP
925fmilhAn2BAocVQpJgkAd9+m7Yw/gwWMp1JA2v6dOcvUENFmcN1KHk4hWVkBb6tM9GmFOqSgn2
AcfpoEoKXS8xRdOTjH/QVmtjqOSxSHLfZUF7z0HAJvb/5oyXPcPgzcE7ckO4fwp8gA5DQCOpp7mu
a7fgK5KhzANya5SJ8AnlDe42TJ2cDLxpStmPS+CD9sJdtOCEkjAt6MA0KIUElzayo7AEA3S1ba6M
kEOs3McQlGPJDYYCpsWK7Hti9xYHX4xbURh4BDADMr5v+Ami1eBDW40TXpLWMlVjCj7828Rni+bV
XX3ATy1+iszE+fRgcFn2hhSTao43nPXN0P2XlJSsifT/s3aSf3thKm3hi460drwm/PS5p41cdoaq
qwyaLKhxXzHGMu96B7TSLOxVzJQmL8XwsOir/ekWQ9g0cGLwxUawEDRHbe/kXacPzncKB7hM9ALa
VE+q6+J77j5KGS/4nEs5W7x9y6++ZxVFinOeVPxs0yNSXkVsMF6skDZvsQZOJ16YJAxymGjWpLZT
yf6aoJOIaroiSEa2L8OGTKomDK7l7xkv2jpxUMHomg4q7b1ew2D/nrimsRmrc0HsRI1dGaCJvDq3
94FC/GNLERVUM80tT3BLYDKJrSQ1se3ahTEewMDJu7CCCqWPf0P8cmYnfmemwZidFSRA9of4CrWA
xj5OEldeP9gdaFhe1vbmQSdaLUWt76/XRvL4Ma4VjARh4HD5xtVE6tEP97OTPl/7vPYHRJjpVs2w
80m/CJ8vMmYyGc+oAm33HaaJU0j3FSAVpIH5sdqBJC3Rp4QQRGp0DofGwh36qqPm81lZMD/b56Dv
LmuJyZSvVGlpF6E4BYGte/EipVwMJBiGxyzJkpZe3gWVHItKD6Vf5mr1RIm6BnmLCtXnCOrh5m9M
VAJStCvmBKRnLULBq46Ea5zhwWKt8UpeyvOztusWawA1zGsmnJGCG1s+AMU76fB6uIuu7wqmA+10
2oFIJ07SFZy8h/CEZVFME/ONMQau58lb/Pcv4oDmvHS7nU48rmi3ULW255rnIdAY0G8fJXe7rXRC
cB2s5V4wEFX/ZyRh1PppCA8ZmXVJI/a1R037r5+khYcD2JCFgDLSyS+j6nLaSqSxgk+InrAcHANT
xtULtDOppSmRF+lbI19/5X5BPAQ+JBP4lv8Ljl4f6//zZBAQ0KnO0vxImzFJ6JfTVkoGthEt7V7B
7mYxsF9W4kwGWxZXt1d94HEzoGVbu6BHQu646OrzGwnzo31dCjKzlwJN7kwIb2cs9jPl8ww2ptSq
9aQ5YqNwIyo9yCGLVYJYkkO/yPSvENNLTx8bFy37XrnJGkkWiRS99UZtaIOQNFW6kPMVg1AMb5dn
y/u7rmxS2c8cNudJvxjBXbvqvtjC41qy2WFz8Swuk93wyVVd/039SeD/5N5yTfdAmWy2n66OXVms
QAzLiYqKxPUw/tkfHuo3/UjjXVelW4rjwq3S3QlCj5uQdLSQxkZJ0D7XPM1P74QzaWvNH2Zzjh9R
Cf5kuBvfNS9TomKatqt8YdgCTWeCYFYzcg43hMfTIj4tsWBfMYot2w2A/NBFypj81wYzo+Ph3Gug
6meiNBowszHA/HX1QTIKDsY6pCb5hDMtcJEmoxHHyLfjCUyyNHNdDTQPyxA4WvyRD8MI1g2Q1sxy
n4UfCL0dly9ZKuY84VOJW4u679qMZEwz3WlCNGqdUo6CfQiF9x71bNmkgWA4hEWz93GUvwQe5Tyn
zxods+CyxXinhIllTy3J41gDlqRKqsAM8D9o/DKOoDwPiyafoh3gKId9gxzXgl/el2DukjYiAavj
34vRgBfw01ZLEJHXoJYUqkupg4Q3qWLKV1R8rI5dH21sUAR7ambpAF1diEMVm5jxPZzraVcqkXGH
5uaRBn8w+ukTZU+39OAS1vsdgvGrmyb+5qGa8LyrvDD6v4hFwC40iZUu+4+Q0HceKYdHJaikBmRF
1N5Fo4ICDzj7Zl/v27AQPWeIoV4VfgoJ2svoVO1lRIktaAkjb1jyH55rcWyc5w0lPnHiy3iekM/+
Y5NFFSt6KGUvYpyXM2QH1Oep9b3CtmRAZyIyJdFB9tTxFzuhzYBIYrmGm4krXS/Gg/PsIracBd9M
ydxP/az6FrGdQ7N05jFpMkpohXcxRDLGSFt4PPMqxUthTh9INVc7iZZW+w8g2LevRKHmEGjpPb8d
n0w+bRWufkNxIr2LmfK9CtAd8nap7/OGncLb7iEWTJzD1vR5vZ52ReZUNuLsrXbOKCDNo5ytX+7x
OdtURPBxslXR/PYM0f/R/+nFVOjc6wsE+bPbuVi4aZhKSpra1sjZ281XqwEYDAANl/g8f28zEe2z
qNyWvQY579plehlYvREvBnnrc13NHNsD0Ptw/c1j9Dw9czfyV+0pyVopD2X7IncZSh1qsWm+leuG
5QT0w4wO9LOYfw72ueuvl8G/IhGsq73IkHJy6C8iKbn15SebIX3bzQH2pCL7veKlqq87/kOG01k8
fIMSbtL1rG4Xa1wCBOGfwFQB6ZMCxbnxLnI433IcYXBhC/6hdb5gb4ukZH6x+IkQnzJDVdcc+KdW
sP/n4pn/NBr7lrJbm2uCNllQHiMrt12+9Ysc1o4Q2ajZszUDG6g3qjosKgspx9D2DpokknIsBpwP
noQJtuute1VDk+c7EWHZfaTyvkTaXKbWEdZhm/sZBmIPs71niPwrn4izdiCspWE87Vo04RBvqle4
KvwXHaLnhgyQ+KFZ7suiKaCSCxVMHVf3qcftlqE+eikYtrdJdNIX0P/Q3azSL/FCPyYe+7mkwYzn
BMWTEX/uLukwjFdu+Au2SfIX7aH5+LTJKITWTCEidChOMiFqn2azUBoSJkyuJUHx71wgEFGYQGqm
hIXilMKNKW/CJvXBNI+RJTQLwCj15COPhm5PI3SNAcANjaGbM9/qYnT2EW/sQNJ0jqFM+BXa9UGr
aebI/uVtJWhdbyUDOEWoPKPDU8bqBXZqS7qH7f8kj1gz3FWvasNzSeMNxf9iwld/7rFnvT6sXf4u
hafe2UrMBOP1t+jgJt663Yd1BSBsPslmeWqmPzntgK5KcyHb53gI/Dz/HwVm07znYAVem94n6dSa
n5EerlYZDY93kCbAT6hUOm4HCd/Q6jewTbN22nqF7zErSj4gE4VkBh0U1nFGfEv9uR0a2KRu1fCZ
xSwc1ydQII4ksOXz9Wn0OwgL7dECU36JN2b8t4eRHApwR8C1BpVpj0p4X2syyeUSWu5fFczM4hj5
PLcDHtUJ+QFraFvhTZYQUu+PPn8oTGzbBUCH2qsFjaW5a6tMw9iqPk74bdZVHN0upiUL1/F9W48l
qbKId0iL2VEspsspxxC7ZISt0/CAueTq1NWbo/0jTIVVYfkb9MgvtvhXHTZwINquEWkCLy6U2J3j
1NeImTUnT0dQxi9C6q3kfJ11VbarLKxEWV2LMWz84Y6lkevkxBn73Q257fd4pFnxCmaKWBhfks7j
Ic6NbqnLZhNrZupIXIq0HfxBZgNHxXhxq5OS9qkj+D60TU3wY5cDiD1xSClTBqIon/qYut4ey/mS
pFGmpl9Dr2nARVjn6Ry1Zpu0nKsHKXFSQFSVHUZIlPH+36uT0r4WKh71HyGl7zWbcFecp2ZQmYAW
GdyoXhPUP4sC++via8AlQnSllbQTPkRkiVAFHNAdvRPd4o12L35koLgg5ehzIpdkTWJ8qCPQ4wae
lgXMmG/sdbetHSOlDRWN/QzTwcio7GaNLZ+QuYuYqdAQdEsA5AurOGh5S3Nfq1fOXMn7h5Gpaf5e
DMSEw+53T26ms4Ugea2c7BKwDdXfciRM8TrrwkAWVcc1DSgld+XNXNGSCtLSy9Q8vvJ155HIUrKN
36/ZrlO8Ws1U4XfAfP0wdkWnt62Fn4OvirHD6I5uVtp7VowUgBQ2y/PIvxO1u35J5ARlksICqb3F
XjktWRuBzDs2TCaguE9ghGgSabk3mEHtj1R2Hsyyxm+YPj/IcCy7hRyujnOvqH91hLtSocP+Ozlz
xJKGIT7ju1kSToeMRvWLs3Rann3vwZ/kkoRxri0nl695Y2aPHS+DmApqf0f25n0MnrRPQjiJQ4iA
OeEXzmWYKJCAurLVBhXf/BTICVat8bPq/kBmKX0NzxHgXkkMZ1m4XhYpGxF3SqzDNOri5olncavM
6vB3gs3y8vW8I0jLpLGB7dWLB/CU+SRuBoQl2AxVZk2s/3G1SPlVY7n2VfapcVCi8NKJoMb2Gi8F
sGzuOru5YE64wRrPjmjao+VWI8JW9oSyG6iQZsskBOwHhgyBSp19uHIz9+7wUO5BRgal3zSXXu7C
K99IJH5krQ9TwvqELKYqe2GWQkHn0w54u35s5oLRp1UUm6PmDbcaQwohpjmJhZT89M6wtpKwLLpj
OTOHdLkc03sMgYPNVQU/llLzc1x7Qfbn8zJbaR9yjdCAHIVoOVItIEDjeCHEY00l1/2Fs1WXmv9M
yOqJQ3Z5LDztx8HmiEN2qEITqGzjatX7ueNdmz3P2F9wQ3U5r6TI8l68w0hZoNFvaDkMseSHnItc
TMOm5hlVF4GBgtQcHGqxWIR8BYFXGHi9SFLwsyKTypZI02aID0Q9KhGJ6XbRfyqV2LnHPm4cH8Cz
RV5pxMi+b/JOye3mOgEIThwW+xr0ZpPBCOH/z4s9iFz5vFzIIO386RDq007srrNPD3eA2ou9xyfy
Oz7vj6yUcFnHrZoj861vRppwtbUcBRzAg5LNyBcI97kppB/3o1sNvs8q/XDDQAmkpYmy4bOD9xWw
3qe2pO2nvMxRHUKPOQAqjSITqx5ZTw2/xIkGeAJiU+/pEadGfrop1XBaUWTcolnw6aMrqn31E298
jIBQlVvZ6hi1KWpEiNKQCpD7M+Ppukzujn/9nFRzG5DgJPIJe7zEMv6J191MseTI7ZsW93yptGQh
KSETZvipNP5pBfstX9O37s8SEAIrICQ4DxzxlhLw/VkE0C9oYpOZAxl785T3D9C2PAZXcPbG480H
W00Irrm5VSmUp782Kr6yrs43JcY/MT+CH0zS7HxmcW+PrDu8zYk/hcNrR/cz6xMw+nF9y/mtk0WC
i76/pfbEtvmOKcG3eXNsDG795LxrjC+PPl8KYGeHYkChv2xARHml2ke52a6zQqDvZDwJTKKwrdUd
EmeVN0XZoRLGh+f9ZEJPv7FdSQXJJgBbmOBw1pAQrvG1O+xs49f280EgQkUUNX0jkoTuQZBwvZsW
/N7w3zhcp1fPAC+KdQptx6tsVkC9iERIkfztHx/ROQgzb4nZIwvd1FPtdyllwF6VzLnpC6anBDDn
3sHXyhjQCwpj7XsnPCY39akT2HnFJ+ipblsQfnD9HwUKXW3vzFBheoqJgCJa8+q1sfR49UjoREe3
knVmtC5UN6cR9ZrC6w913Idcajbr0poTpn7w7fwXrL2jMQh7i6fxyVtp63CyAFJ1S7/kCDwwgYF0
wbnMkC4yHf6me6McQbCNuIoMqu3FUKyPOzVL/kkwZfkUd1K2E3iRhrmCfMpJk26159OQbE5Pqe5v
TDEkD69XhysfPi1eSI79355hn3vsOvP3b4GIY1iBUnKXPTc4+WCiD8heMIgxGNe7IJ7THoRjGvSf
n/ZXN9sdcNGqZBOerQxWPL7qJ0ExsoOS75is0Ml6cDwrs2pVsf/lvvL8A8j5ztcNTQnUpe9BgcvA
1e6uMwPWy129KGLOzBwqoGbrikqrsiE+h2uwHWHJODm+Af0VOvBPdzSIftUcGtnsXrHLu1Rfqgki
Tu2PIktlOz6Y9vHrGV08L0wwjth0mi7Y3CWCFt4Bniffdwg3D+dt8HoA5rovpkNSEeY4Y5q2YvYj
pGaWSWbXlMIVLYD9Ty+qrRE+woqHhfpiTGFDVB+jrXTJBHmBJc1dHcft47TZcuwRiGq6jxdfQ+ES
HYUM9JYkQcAKxHo+Sk94OPfdsLMM+L8DFSWx4FuAFtj3HseDqUNJMS+9/xSMLspUYimsjBwV8JMR
xyUG9qLyrg17MuHxk8bdM4OxuSySgNM3Y1oGCkRD2+KND4Ga8igkE48ln9X9yvZxFzxAs1YhudTt
Ic7IWUr+1zSZa/x6oTJaAZ6CjfCmbsMvQ322WpnGGeg9vluYychY65wh0HS00Gmu2PF1JZehCLQh
my144Xpgq7gi4A8GwJH5mRui5VtxkND6CqXongQhuWpcLerGnbzPTaVGZfeFuWcxOCRx3rk7/fFJ
eI8xuhGc7r4rRqBUORvj7mdI1LK0XZjLixgWwbhmZPm0ff3gPMAWDrgkzVxPsjKrUtkaoTexvcW9
H1zkEtE1Ey7epAQ2U2VUb+fY/ih6E14DgUcDSTEv+WwqDjC67v2ZJVFniu0ZELPQ/1qk735h3kb5
FCPiUghxUDd/J5Vxuv2mCetZP2upObvJiNYlIl0T0fWtkix6LcuVHkVqD5hLEoErcAEeuL7efVum
f5AU/rsVh/nxCYHKWIQLBch4HuQyEGfC2Ia288dHGSf8m7nmCMrN1XctAE68DFeiczcY//aDAVTJ
jDwUOFs6k35SwUtyHEKyM2KfOSg0qCoqKKq8akN1GrdY34oLzKsELFdoh3UhZx/HwEh2Sd5sG4oi
knNofhkH7DnjCzV2sxUwCkZuBHTzcDe2tNhHfp+hsIws54I++7JbHpO5SINLlZW0CXesa7N+A5pT
BX4sKEjEeRa6mrZteEhyTb9Lc7Y3yoS0wriBCDlPE+BPx09y7jGHEaDDErs/3tAiwSvs5fR3f/Oy
wZKTq3bPZMN28JTc5lespAJWwJaxB8ngDQAcJf5Gy9O83UWhqQvORjmsoHa+B8ND94LMEE3anCOd
DfkRh0Ops3yNLBxqa29+RUkbyDnrmv6+ZCdGeKAtLxE0dTb+ak2a/Y3s4rWhVhY4kwqIZHm8alCO
bss9kaSKGgJuQ+J9QdrmSM6OOn1cj5cJGKjOcdf7FVwQqkF6pGG/BJSfwYDw3wMfN5Nt2wIWTEqE
HZK6xCJeDozLKvwsXTY/QKHO2ZoXpOFAIMt7giIh65mSPTRTZYODZNDXwh3Ate81GA8j0HOVEZrB
M9MlK9FJf+E2crpT9dZPctigIYSDCNiMJJiv7bh9pVluWwU7/SrE6M1Li8PB+ylm53dtTVeM2BIy
xGpjr1RHHTsWZfpClT6t+kPdXlB/eb99rEVQb8rWuOih0ulE4TEtB8noAONauXjN4EbIftPmZNPc
eyXWX5qbRoFUeLEo4w7Vm52aSwmaFEf9TOL3Ct1w4JG7jLZWs7hbYYa6O5tsbqRNrpSaLGqStCaJ
My0p4k5n5KLUsmWWLxoxQ1be0iOkcc7FiDumtoMBNbE5ZtORX9HWI+AFZNt53ALdPwNBpnvygenm
POowi3ZK5rxL22FrtGV80hw12preCpLv+e9w6eqp+9nXXcDjzHnBWwgC1SxX9XMNElWt6LhKwMcE
4qyghG6kt/ZyBifPSb8cQ9uHk34t/fBVzPmULourofigOs+ODXz8iFkBzHwPz7UQSHOILT4F4BqS
A71b9XS3MfgJlDJzjzbrU5TAuczgfC+G15lmRkUUtneRPcRpIrr1VXKLCUljb4Zt2PowvLhn7p50
EFScpdNJJSf7gjYSmxD5NIAUuj4atduFmxL5CSAUmqFQdsJtTDMvtdyJZTLxJCRVUBoQlpYAMJ4l
wL1sD2l+vMN/+M4pqf7nQF2xvniz3tAT5DD+uazs+DFexF+++MghPEbQcbaiIOt8fz2mOIdUrGZp
Kaq7Sjg9ftpAG1kFWIRE/WcViYfFUeFi1vR/Xi2gQjToQzdLqnMm6Udg4rYT4FPUcckEwylHYJVo
57ERyCsKrRTn+YO6/dV4SN3KBZ2fIDDQLVx4TUNRFGicUVF2ffSuBdtdxm/+YQ2qeTUGqhmoQVo9
I5j3X7AoCqiWVKoQNtl/h4vHLi4LXM4iOxAo3jvtCkP9sgaC9cxw/d9z2xhqyJcfkO4JFPyxAQM2
pXIq0+WQCWt6bOq40f7vf5O/4TqGgFLjy8T3zb/Ty1BzmkwI8XxMCIfvsXW9Vava8dMmI8A7t0s7
rFH1mNGQAKht6gQDHLO98AT0oT7ZzBTTZZRDgbVrRCdLGF9luSgJ6ePbGzNoQbP0bjeIy1/eKpne
imtu13xb7nyA60IxJp0T2qH6/14UQQuidNrPdOOOktjpHPi6ZH2wbcOQzbBMs6eswbSm0WAMdl+B
tj8MecU4GxpeeV6YySUhYtrbqjTREfLF+qoFpj3sX4BeTizgNtwATytxkM+Zn0FAk0qyJaAdbmBi
cS+UchyG3lLpAI/vGj3thQcRkqR2fVrbHRQ+vQ0wsbYL3h/Siek2fkl47N//HNWfrXjzWWb7OKFI
0jD/oAqhoqDLQ1DiAZZPAShyG1ecrVp4VhiYgDhdhFiSMiNCNuDa/ZAjaj303gILTQ50++CS1acU
SQZxP6TkJilmMcN8D8uusFlezoJQQAH377kPmxRSfTV2/HkX4/6KZ/x2SBnpWm6vKOUv+7dbTp4z
UxomjmQ8Scu1qSbiWCQDNd/nmbePtvxaPue9leFe3USphGZLnDm4g8eUjDOc5OF88gfzSJMlUpdT
69Go8CHDly8HITp7tkXpuI8g3XTdTu++elthmpyzIXx4MmvGwLPYrYnVb2bDoNROtYLm5iSw0wMs
a1LAdqsnn54pKYlJCLPZxNOAyxeJvOlLFvz66alZEqP9HlMNm6Ui1oHKhFxbbkAznmX3objlJTwW
2Zljk/3z605RCZZJ8CRGZX0qq/eC4ZkExYyVc2t7KdAtTXXdrL7wDx9quw5Lkf4rR5hPCo1e8ku4
EwImc+4wPTrDyUs78uiYxA4SeFpEmvHbsipq9sI/0ELiR7A9Ffuz/IAd3ruzXK+NT1vHoEHncv9V
Wc/WcCN6KH4//2uzQoC5x1lodDdKHGoccMlgBxxrckSGjBfMxlLtlA8vjehtRzAuGyFqquVGe30L
lE74vV1pEh/SHLXL1XdINiJ0BUgE4bnCZNv7a2f874hnoC/9BteKfEd5HWX7ezViCu11IrRA1wKs
glgaYvqry40cI/EPBEln5m41aFV7m3Uzlp/Q17CK4plbwvp49ZmLPzDJzQPpUrbLMXp089xC7d7g
Yvii9RdHGXQcJ1SYwX5mv6EwNJkuuApN+BHAmBmPFnwswedLxjSIIw7OUiFaOdMwteOrFmYZ3zmL
M+lcMaVlAZu+3jQPwysUFsrw1p9g/mJCq4rZgy0vzxgMTqA5zZ5mhtuCpVMUDDc16ruumpT9S9oh
iE4QsPGj2f5x1I5FbFCKwI0fphuJ0rKFIqnGgDutOTCAYFyz/tK36j83eT9j2irLfecEKTFrBy1x
ESvR61L8i/0H+WPGYouFhTKlpdT/WN669EyUf8WXr54IbDb0ERCZfqTidYqjJX0LUhjc1PaC0iYD
jew++oHSnOcjSX+zA8BP1XGoGIVUtTSb1up965mkfX6iiWEGrxDldn84bSwJhfsQxqu3Zt11eJUm
rw2Bjq3Mg+Ja/WH09wIRdGT/E9ZAjMXeD5QxhC4TBKiF04JyVIACyDdviwIRWHs5Tmj64fsgxp1N
JFo+zVSA6C9R2J35x0j47erl//RlhUn8PkGd2lIxqGsl0uvf9rawa4pIK4pAuuDnTZeWX1LFMiaJ
X3UrCnejHjn2J+7/UTxmqBWmNfqrcujQONOalVRImejlwtjwyVInJIMlph3OG795WVm2C+naXfDr
yfQ01QgoSQLqbxS+ULImTum5JjAQ8aQ8xR4kezyO+HqfJ628JAoZzQafHuS92gRkk5Lyx6qLuoKa
w4uJ/sLZJWS8zIFK0Ouog9MeT60o9abrP4bmxOvkWNecc/xWfzMtxjSqnBAvYG9L9oESDyUKYqeE
pj+nZOKvkl0shLK9st7xL/pKnme911BmbM1J0V45+v9AGyYltdaWQ906jo9T+opjDwSx6MHDkfeX
IOCmXl2NruQZarPQrLXAdElmI4JwliG38vCq/n7pxX2fT6L5pnoHr4354Gg4goWkgpDyTtE/YeJs
83FiyAWwzYksFFhbjMAJX7kLV5bI3DIr1TlaEPA+cWQZalkoA6jHNd5LEdKvmPzOfUueeNH++ziE
9rk1qvlCi/54gjGUY7+dGSosb7Uecdsk87/i8mjAtH+W7gUOU+EB2Jq2K4xTry4k8+QkVX/r2l5K
Uy5VY4tbYVQXH1REjje/dfTyvIP5W0CZcnBpauvHDw62W3uPSYiooKPmUxdoXgRuH4kMW6d1C5FV
gnruy21NJ0sI0+cl6owv+AFB8IjUv9uWnc7fJcgFynWfno946cC0EDcaXDqdPaT/BjvJk+Vv60I5
t/1CpT7cXNO/S0UW41bDkv6AeHcRCye38WAW4sqq9oKjZbRpmm4uIkSbK7/foyAuCRr4kze1996P
lbL/AZcQ46Tk9fUO733EYBRiqjFAyh0qugjOQctz6eLZ4LTjKZxuJ57bayjkHKGNhPZ4SuMZ9ZOZ
hqC8nq0hjnxmJ2uwDagl22a+wSVgByF0+2ATJrITbq4PZssdxKf2zUHjxBr9kVvDo3Es1xQ771Ng
6saHW5/hr4z4aKQAXGhsp1UwYnFSAF/h7NZxwLOhuzllS+dnmwDUwlwu+hHsrBEFME2HTGvHDwZO
LrYEd8PjFRVHFap72V7NSnyGhWeHnSv/yhORSNbKB12CKPNmjlhsBvyNQb1DUqoR8JkTEvsJyZmy
rMZwI4BPGyAlPv+Bhfc59eBzPvWY0kv/lUVqObnxX+FsaCbFqx5jM8tDGbQDWKMRh7N1VjmUQNaK
8dYmShxjdFLXW9cxCp2dc98nok46KivBvV69fPuZM2q6VwjRe2ZAn5EHoBc9AjebxgggGZPQl+Uj
+WEnQ2ofLKrDaqRkEgG12PmpCRTyJGepcZr1CtTK/sYVocg4dkmSThSr89MXS9ytwt3ZCdbZ9uGB
luqTG1hi0s20plcXcB+jXkBMwS8yZWtFn6URdtazuTwf4UJzlqdyrJHBbkkVQ//a3LnBMEz4BNYN
NNfe1x/h1g+mUwb8yB46zxyBl48RZOXBdQwy/kOJDpfNbYIS5Iy4JFBpjy88SCklms4SKkLsJPD5
RDxcpuW7EM1wPPb0OiVgoDYd5sEb6DNWB6fIw2kaGmC+bbZX4M5le1YyzmYddSD0PF22pvcSNBhX
D5BEZMTm6TfKANNHlChii/eC+DpoN6zOychgvwGLGn4WuT8HYR6Jz4w+JnY4rbawZAWCscR7/E/n
mzgeY9oL1R7MDYiPIsSOTKYu/g59Z2iPivaIopWV97vG38dtifs/IcVqnEDDoC3bOci9C/i3uXke
8IipH5TjHIxK8oH4Nnobgu5SFHy8FCnrqG+MIa/1f21F/2r1SzPrchmHiNytk1xZPRVkvRY0cDy+
V27QTbbgbz0ZtgDDkzvdnfJ+/jdY9RNe6P0DN7Ek/7jnFTx+mgt0ICAYlyp8gEP5sA5BSxUP2mSE
u2DxE8FW+4ahG7Q4IUzFCjKlSnJsoa0Hjiucp4K+P7kyzwMeT9cUxelEMosJl090vk9uFRTCKhVZ
4K3pEwOPGj6FXLcgn2nTy+V/kzZvQW1ilTKTqTUw4g7lrpQyAYaugBijFDVNScc1BQlZ4Ycmpftu
4rbYThr3iIGtFoZD/QkEbU03tQrOkUtqjQ+qmq/mmfnwj1/RremL/fv3aM6JGmI8CMbWM1UI2IT7
9aRovsmrlRuVlODs4m8pUhPrh6/Rj2BnTVqA0cvTWdZc86zTyPebdZXRlPyRenLnHtjFORs/3fMH
7crFjYvtG3GadaHrkdX43OuDdgbZj6tZqWpC5dB3yTPqmoAyUoL/odabOJuqAxoo1p9+OTR6bI5b
5/iUr6sq6HOGKlAS5bmZJi7kzMx2AASfmXo/tYhDt8R+gu9Vvmx1tAmfZf0BRu9WVsCKFjE6CFIy
t1hlcaUXyoH27C1HInDQkzimujDCq403Mrt9ph3Cg9Vjd0LIVYfFCN9S4ZjB+e/VuPg2A18ox32W
MPWKUL2HhoKWCCg9hGBxmpT3X1Rj3phKUuWKNvapzno15RfoST49keCCPgmAUzVR/f4TMa0KOWFV
QKJ1uZJqF4C2DdmjgxoMR5SOU1ZpmH2nGf6JJvVNy4702gIpSXu3gdNtuyr037jH0aWkd2wsqUHq
UqQiXlNrTJe7OFnCR81eImqw0tCEVqYandwLULkWS9mbOHFXo2xVPLxtYOz81PyaZQtjibH50KdF
XpwNpPagNohPwkN4RPjY+OBPPYeIoBIYzQ6CGkuhy21+jqwsbRWgDqeCdc1nkCcL3SymhkC/Cvn9
0S3bzHe/SVZIaBdFdEYd9LsmzcE6OM2qnDp5H/RSx2WJEsIiRknTCB21eoVXdEz3Oc5Lon9i98Ux
gUyplkSIBwk1dEzd335mWQeA7MvjqsNIqED6txqDgSuqrqXkQJMIoPiO0E6f3OF6L80DGSs/MG8c
UUYd5LQDeJc4YIoMLsGi9QYNbXNn1R7GQ2nkpzp+iUK/zOqNCcJ8y91Bk6Zd3x5mnf/0OMLxZt1i
7RRFw9iOXjC9hBR8v/VQ3uWMMVavTu+Z3dWlz81x64gr13FV9ZEz4QFKtgkrp8cz1guyIehwXmTy
osvy04LapHePZld9PvWk2UUBlcRauKaehkWIx1sxuAgQWX3hly6CJccF1rIZv3ONh2AqXjyDR8v6
91ODbq11Yhl8LDBCKjlytYOf9LclSXv/61HqHKjKufJEow3rZXrYGmzlWNU+AomAxV3j5JbdvbY7
C+Gj1YqLRcgIqX8oLL/HPXx2BBOO1dXyr5m9/Ui908Lop1JFkcHAqinh3KqXDuUxcCGlRgXRE2vE
Mu5LYEmRnk8hh6fgChQhxMae4yh6m/zlkjnxQSRvKdVgTAHy/AE8DNEiO8lnufnONmpuSKu6q8Td
N/IQQvvdFEbCNOVz1+4tjtFdBQ2Q+52SnTm/JQfjaMYeoSGbF61NnEQnTV6wj+wHQkpoK4ZXuGcn
YAZQrO92RHSZrT5U2yZCJLDqGqRl3dX3OHVfrPQsJ+/JjJ9Yy6cui+CUOP6FbMInoxpp3Erydl+r
oWpPz/csRiGwS5K9lBBwl0DBLSmB9IvRGr0Vmq43cqrSfUKIl8epc9KX0SPdw336ajh7cuHeC38A
SOC+ZMvPEP3GF8mKI2V7PAEonFkE1K6jS2gAxa5MvavtAZ1awT4FPMPmFEK2XOOwKr5A2InzCzH1
f984H8Tkt/WVufN/+fCgHR3dIOZTorrnqNR3pfjJWRxAn8RmjysvoL/rz+gcnzIo3FlIsOypFReb
hIf+GimBInIf30nGUJDqk5SesQFsmj2lSbr2p8hK7590aklxTNY0/Ev4zc6H709zrJfTGJUohJ1y
jwTgO6XOFIXgSFGHV/HCpTF+6UIOTE73uOyXhgB7ZpQ6fjym0RI3uPJm7VtejWTxEUTZfOeu//xf
JC+HDgDgBXINXZr5E/jf+RlT+ClAdjr3muvVpxrz5p8nANnFezUEPF+N3t9B89Nwf73cO8iyLzXC
sRH+OdSkWnCc7punXeUt9h1ZaBWboiGCFKBxgi9a87rhLoUa9cZxYFt2o+MlFywSzk/KhSGDamZv
43ksnPeK/KyW6XIytJND+OQbo/WX0q1DnXmyg/q0WgV/rwzksejogUQQARFR04bJ45d2oHmiR651
jLJqGta9xQuYDHLXIcNFuIpA0RlRE108TU2LQRdsjApWNp3JmevOJrduLqUQxSb+wKSpDXlsiEet
sEVFw34Z2hfGffUALLhZzpS6Jl6xRJIHNF1FQEYdVHvqMTSeb/H6BUjPlTatoOYUIorCeyhSPOlX
128pLAE0f1EiviDUzqUz80POKhfaj7gE9wCbzPl/wdI4xcT2WezATShHA4TkqVwgwyQKmNJ5Us5w
wCHR2+cYR5rbFVKHhzCr8r2D7xpUVHYd3qB6bBGBNf69aIG9ip6UR5bJrWm0BBhq+nv2wUpd17P1
XjS0UbmMyZJzLhkNIFJKCklVRPJ8MKzXYqs2kR4yT0YqUc+xhZFjwJIxxp/zV/NQazmml3unGLHw
Nnl4aaOc6Qry/heKFUMT/CXfE21Co2hGsJ5t/mj6mn7eXvQCx/A9ezsz79UwyfqHm7jQrBXK8qaS
/1mEohjrIZuPOw6Ec2XXlsiE7lzz+l7AqrF1K6K1SV9hOE7rt2TRqZ64HQb5jGSFrNgRp94t5eWV
6UKM7umit32++rqDwjQ6C9b73K6nP10iyEcTWnixB41bGulmZCgNcucrWXIlv/K1HcnuGLL7ak0Q
cmi4N05lsFJzoBt0KfFem3MaSbLieBKZrtMZxTRk9cvJ+Z3/9Wjn3vHO5Jo2pyZ2iNSNgjKrnAp/
+fxkdGRhyiGr5Zq6CpV3bEJyJyw2yhfI43jnIa64btyDwMgI9TEXxMho8115TpDBNeu9s9J91eYV
jtR+PIBXNWe4cKQRUwexQhCXCm2QfNKq3fy0Lwo3sT2/yOMXO6ifBUlvMBH3ZVHDzLDIicxMAAXy
992gMkwuxhKiflYs4cXV/b25EWHvqzLAzIg+lSvYXJtHA50/MI7QVjU3EX1W5ZkLZX7FDAb+2x2g
+ZDN5XUbSTVlxd76/qZQHsGwU1/oYsqLq6jhJzA4UiDpus//zlKpdr0DKHcEMlKyidurC7PBsP/U
QyOE4DlCBznk2b5yIzpF61gxgUi89nwgLB8lEj8S7mN6lB62as/Oj6lQtWss9zSxguMdC0pOOM3x
HT1tMR7cjH4KXOhd1Ijl60Ci47gnFFC5kzFPFEV6iDIoe2Rj6QgORWyrDGM2VZcM89NVvMGNfbI2
ZDmAanT8DREvTRwUyyoxEjkEJTB6lBxBl6oebzQh8jNWHhJAlB4mnsEnD+ZU98OJ9eknvVpz79eo
+mpZ705vw6CDwQRs5Erf/2yDJNBzaPPendC8q5Zxp0R/CcNZ15DRjrK8cAumnlu4Q33gz6WFP5ap
hf7QUwrdQNnj71IPtL2nUMk5ovyZ2tVxKv8kpqN0S3ZHkQRhAKE6yi59+FunzA/SLAkSRjrECzf2
zd73s2arUENi5778PoRmt1ttu+ilr+DAD1Dqk0Yswk/H71uorCLnQjonUY75Dw1ksZVTG5BNfR7h
UmLd+FEKImmOmjMk+eJ30IYnEl0/3k1UtvzkgFFK7/1bnPjqz7Lb5e4rSGTgQADRUB4x5LPsPIxo
T2fsON/iCh4y+gyqkeLEpKwJcPCml+VM8YHzabtokj9KL0JSyKejnYElpV0ecUjRGzfkeKrkZYp1
G5fElCd1zLsEP8HA/aC4yF4hHaQIO3c06CWJo0ZCek+HAI67vLwiWEVRuNuzp7vZOzNWQTV98n4a
ZA1VDMzlfV5sCm61+wkGdSssgah4yawndNUXa3Rdjc3dykD+g6jtzRkko0C+WUer9BXfRf18/jRz
ARcW2ucpnpgNbiZRZB2uYPVSqMwiwATmoGoBMpQdN7NIqJS5su5CQ9rlXVTJYm2h8syiezYmJtEy
3K+ZHzkaNduddGvn0GfVChNqFFGWNkrt4yYS4Yu4THbHhMnwCff19VN5vwYiI1Yh5G3fP8xiJEi3
YrMD5RURjCONrpReOb+8nR8w30FwDgLApUeVORUeyZlJWwxK/L0A6POCr1/0YmD5ulB2BXffJIIG
w2JCnmmqa7wgANT1Bk6j1/KOiE7Bg4pL/Zxw7mnwduLJUr6Ohy33i2Uz2fDvkBmkRRbhBV0p0x7V
nmsNu1UbniO8epycwo8/xmYde5rXj8cDYrHAaYVpmBzil/2R5f0PNaGJqmdDs3zp4EOLWcti50BY
STMbzFG7hKGO7mcY/TT+eGOjzAdKCRjxG3ZRYVjecWxfTG5nPPUhhXeh1xvWDOcVtFH0IQZCP7kL
HLi21ijIXUSIjnuwZyxNNzWaGfcDrZw8v4QJ2XfPs0QQYz7LJtCFQqwQCwUGTLLDL2hJdGiLajCH
AFHy54Tts05UZ1V+QCSgHRUdKKmEUuC3ja68bDUCqWIJWumMhSJMH5myAKqJ42EH2ZvBZrKB1TRY
ng36/O/N3mNFz5IXg6bfgc5dOiKboVRFFbyJAjKPFlNLS7o1zmRdPcJ9arAfAX7jsm21qVoplQ0z
It7yk9me849+hXBq0B+UrR2KKrE7W380qlOIL9BPRn6eCcl2kZ38vuxsWwoTpB9LKHtRa2YSuk2k
eHn0khmAtE4CfV+mLaQ9UPpRav4W0RF4GOE5Byx0FaesnGyhShtZ5y27G5gyrq0T0rezHq5CbhUT
+Ky3go1rUZWFfwgX71wcMnLe+9c3Jz7rFh4h+W86VzlBez4gqwIuG78fSUNd1sN37kdE04uJDnF5
0BfI10ImXXlmCtkY9x5ZQzeFod9kkTtVFf9Kl5bQaUCKmqiVUrA5ftRGxB4tTJaK8JUcMg7JWp0x
P43x5LHUWXki0DsQuqRKF4WCiehuRTZ7Cf72oa6kph2gUBzX7AWKupsCcL+5gvUeq+Sk/P31Nm3c
9n3J5QMzBRpCO0IJOm0BWTWA06eEWXA/eWPOm1M//6t6pZNx2dp5yd6B+bwkyTWdLnvGf3lpH5Ua
YUqp8UwXW6PwnWvwpoimeFyNJt6GV/0Z10jxo6kD9trzAEBnz0wK8kbrvBmF+DgjE36aKKRFbUxv
k+il9AzvhcwZM+ASBNqvs5NMlgrp07o+ruCvoQfj0w0T3UoPwJBJCPeXcdjNJ33pMPhqf7bZeymS
zMRRSOhI9IjfuKdFJBj/eeGViDE51S7LOLc5EZkGVPf6Gu3wAIQIGlc6+pjB76KjLnZ2vYo/lEkZ
hvm7HKsYOOskIBKRh9das6gluizBkZIGfnF6maVSksmXgk7YJFg483m+KhwOqQbIdhe+BulYxBSQ
zVpBP1+uP3uwLYtdHbnh/jw6+x/sjyGaqyxYm59EtbSeShhlqQ1o3P7s/gj4tEOTA4lp4KkOX3uv
cg925klbb6UtctPJWJ12MWp9eoGbybhNh8d1+ZVo2tedc42HnwqeOZwwg/13PDqhs2lHyIacRciN
xbJqd+LzwXGNjjHqIXxBJPKRXliB8Tito+/kR+ilXobW9k5CJ4rSnsrT5yc+924yW+ShTSqu/o8f
Jue56tkUdS2I9qMKSL0i0jXmqxpXWYuNi1VbW8fAgCXhPG4kUFa84NxrhI9Cl1VFhGnkAWO0uVzA
VZ2s4rwPNf4N6dEmyG/3hwFG7cSebChpqTDGTf+QSWjP+zDSW/QpzZu8Gal6b0t9JuliEyntsjp8
ltLQ3N6+dc62RJrUzT7EDPJMAfESz5+gyg8Xrv9Ha7SZ5KOyvVI6MWgsUu4UQNMZ4urxlPNf2w8X
PQdX6KRK+pyhfWNAxyhOzmeFwlQ9ev1sr++0SVHoAQ648b24yYLk8MG4qYj8oQeXHLbJmX4Co3Iq
HmiJxNz99f0v7JSHFTz7LY+cCRi2r1ay4ZlQfHEPbq/pgr+zWFiNZoZruyIAaAxXVjSiezwo28oR
Xx55i+J39c1XxE4ed1L8nhkQcS2QNN6WZuk9PoTYqJNiyKddtEhuCGy+81fcKP/X9s2QdzYJAPjY
ons/kSurGaacisN1E1/ASthqVVztPmJWXYfC9BHy+lzUdfZZt3uXBjdNo2+x2s42kSgR07hTp5bB
FlFpH8D749IzlA65EDWDS3QrTd997MO0dKpcFBacBdmkSPU0bzVIwpPgDkau4m2vbL66MsfnJ4v4
xHMqfXBOQfeL/nJdmCgM3ItBrs76DscOEgqU1a+GBtb2ACKwFjeQY2GoeMe1vcYVEezIb5a/xLh9
tCSEMCWkcV1pmVk1P2BbRFgWCFudE7n0/wH/XY8ZBAvv4UAYCZa482j/b5BfKCSeoAdp9S17Xynn
YpES3MW2QGPVj54QM6DGSJwWCKGuVC+O8OqRP/ecIFlA/NSmS7+TDf4/ZgB3WrmM024GPla+y6oV
dNUrfK7URdxf8FJQD3WrGcTZI2an29O8K0/TfN4QUXOYtF9jNjV4AUNByBYAWngt5G4fUiWrTGA4
Z3R0WGayfRYvnlnRXKpG6XVOrIQ/JNJsI0HGTE8qPu0C/pUx9iYykkEhOeBs0WwTso/EKF6M54sH
2Ubjmqi5GzdS2NtjcjVfdesA3/blLu7BqOM7F+k7KK7dmofLrIJ+qeb8iPB6V41ojdAXzbJ82V1F
r0gD3Uvr4BXsBN+qpHyS1PZNPKrRMq23fv3jJe5iw0HID5jBFe6HT1Mr6r4+0WkDi5qqJXVVPafB
CXX8mgNwyD3X7QtEstCyL6oOCNemqVnywiA4eIz2C0a+if7HVeKYVxbSmheUjdouL3xc8Vn0nJFp
Ghydw5eOtW6yaGgfP5tw7JY3wdZvZclrXiA8lSufELJpcwBnDRxxyrXxfI7r+8axwKYYHV/pR+V6
l8UNil9mLIwh4fVVdB9wMhmERZk2lH1iqFjH/PHTeZx0d60Un5enb+FHOdV57+VhsVoRI+XW87n3
rFehC2mgV0JXXqrxokwZ89HErN5TTsGuP56Wq/ulPV7c1nN3B8NowD8CUY34HCKcb7khpZxpD0rM
aZ7ytfLUowQ4lkot6gRMM1J/jExGMKg26t4T19Bz8TA1VtbCBHoPj4v48Briv5/3t50p1IGxXsHF
7EQnaqCkUeVba4iSbQ/SyaoXPucpjfVxBtvkvU638673RGM6+cG1rG/1Jr+nES2xBK8birYhtN5h
D6g0gsPjCs0yNCe2rGhyMyAxd2AbfCoKfxAj8kqgHZkeCvyf2Y557Zz6vG6kGWfjRUpVtHRZVPwv
hE+BybYDVNzMeYGkKK9BWtNM0h1QNpPxyNz3lrBM12XWnhxN37E8eVVpXVwPTzPn/iJtZiEXDMcS
xRUyXiMb92hoAWA1dCVSnAfqTQFRhmSCYuq/ruR7YiCu9/IyUBsTgriSmQMDbyDOB7ZNzFh+GxGS
SNqVg4dqxqafRtPfi4Fsb2XuScfI0IkDMfbI2GrWqsdAG+ScfShz6SWIuCgP3wrHtxyC6VALkFgk
weaNwtewyY4OaG21WMrglHcPEFHmDhgSiKC9yfzMx8hzF2EBsjIACS2UT/xyyCxOJmio6xWO0CGy
d7GQjpKHHn68LdlhqyRLTO3mpdt5gW2JiVHmdDKBpwWh3f7wUScrnFe8BgX/VtujjuBD3uoFsmrb
qBz4IhXfaRgEQYwp7xPY2IEbRj2QrMuuNJ8na3Ml9zPk+2GPf77pijN2LKYVH+/r1qFJ8FD/M0Q1
wqTNUn20/dK0FN4m6e5iHQjMTsIogJAJsTvzHC0xAYtp+0cp7FK2+7EIa2DDJqrQ5XtxhBRr+x/s
Y7KF8ClHDaC8LT69Y2KjfaU/bfzuCxFvKKJUDs+QeIU9iObrPmyojml7/qyXex/mACjKt19rwuNd
oazPixdW/s3pQN5KGGdYEb444B9VPdwBY0hMcmu3OlLOMyd6tWgMA0WigslBvXQ64ccbDFH+du7v
8+l8LG7PNoR3AC19ohrkqXgTaSE2WqLq1VuUfZX37+XK+Fg0dHqYVwhzy0vlnTn9MOoRiWY2myAt
GQXFlco2Uh/FuiS9JOt/pA6ua4aNC12VgtyZKQHYCmNSLTLS8JurY588kd37CYSw6L7VZdSq7arb
XuQ3majW4w9mz9zaGeejVWKC2cXR2/IkV4jXCMbQA1FGk1mqvQN61MXJUOZW8LgvShy8mIZya4bx
kGyLhrC4DfI2Q/M/QjYXzYB934pbV2oqv9wCotcLyU2dtKDudHWMDuD0IHiQqYlcDSr4MXcT058r
xEvU9RK1Tty27TYICiN283BXhhaXyMlxIPJCic6JTsEfwTGTJfrzgbk/NMcy5+6PC8YyMNCwGFDo
GdU2U2mFR0Q2HVwnTavdKfYpEDd6esEVDSMnVeor7NXudIfiXTo/P7NmIzLL1HTrjq3NJ1tzf78Y
/+bzKLqQfCUtm3NehpgYbo7/LB0ae3aRrrw1L93q5asBQVvyWc51oWum/xBhqzaqs3/xiwnC4CD/
Knti4IWA1DNC9/332/6fkwKVWg768Iidt7P65ZNdCVT+mt3ts0EMaP8LFZsVjQQ0zMMt9w2VRC9B
01CQ/54ovvGZWRZJy01f/bHrjWh+3g6UIF/TmyEm9HTCDxyYUV0Kab7z2DWm/ggTJc5ynxYMowNQ
clXI43nrcjg6rd3sPiskhnCq7FWbzujY7mudCjV3mqm5t3ry0LZ1Db1VrP2EfRMFF6YWvr9p4gLr
pN5MdkWk6lpPj41TJFs5Ol+sZZGTrttQ23L8oXMN87CZEOrEGNl5YXoHekDwf8OPSku2/khKluQ9
m/yKLz3r79im5QlcTl8/qvBKrSaI5y/7XDj04Kg+4LauZGb5TEPiqxt7cwkJccY4ZioJ6Ux1FC8t
vKcL/2/VvT3d+6yDVRdrZV2QYPF2MEhnaGxx4Ekag5CJ2kLBJ4+YrfTfyVpksmcxcmYtgE2PELSS
xwdXylDvRz1DGhKIi1Ct1bA/IGYk6Bk8KfjihqYDwQrchNGNtEn9hy4KXKvjQ6XENkeOP8cGjtHy
jwNWUQK7dyYx4jnaT9DqfWzxllXSPxMj3Z1Au4NhoWvTalFYuo4SzfxIEW3Y3+Mu7m1M+PsQlZWM
lUFI3eN8jQZxO/8jzz0wAGIJ3mbebZ3RM/lw9VSoe5vq8OngRD9pU84O7iEeRNoeHMshkOwKsb51
To65Pkh0F/Q0lXhQEItwQfrWhFhHqYdLCMxtqA2nu0HrHXJChNMZLvM/yU0Fk64lmnirIC7lcFaD
Ywebhn8CNWIKpgBXIHLJI5FZmuwTutYi2NAXKAKUmJ116v5kH9jPTGFEGpUCpr4EZCPiTpssrCSM
Hu0Vbz3B8tIg2qXSLfVQftzMxQVhXz7kMfzfNw9fbpHIECyhoxVVeERrsUcn0kSDvHZVQJpY/r6k
FJbHJg0urLhIfu21QI+e8q1URZROuvdOseCmDlo85H3OAuPNHFA70kdwdIIFcNcgpAIQZRSH6UqQ
Cq02gPT/yBqqYOVsO51Dys0Bgzw4KWIDt7jRIPBhNQVqmauPmaGcUgQg80bTNYnGdbRPmcmf3AXm
YzY+ie4873iXeZLDtPW+TfUNatO5Z5Q+lf6ZjJnJfTXLwK9P+z5ii902zfI6YQuO4Jc807TXniL7
NgANhGiYL/sqVnFqTf6zV+nMpm6p2jtBJldF1F5Y/s+qrSm6gBbu3aDWFN0gIohLcu7W3BBtxQxj
QCVa6wVqGWF/rqq8d6w5NVke2UOMkk3z+/Tte5SDuvyOkjvYCA9SDp6Uv3g4U+u/dAFFSjPSmIPy
WM5pZqVyvcf6he7wf/47HPxuhiX3l1FCvr967r4GxEeew92k/QflwhZdPPIZILzhpFjCMTU0i0oJ
VDyrivuXxvsafBJJi3BNwb9gTCtaapDb3qYQigFDXdF7E+Dk+HwSrtJk3Q79vSehtv9SDj9RP8ik
AYXrvbf4VrFacNNeIrSJPTbaSmJq8EmpudyGmK4NxhnD7ngoaTcD/KSK99tXtje2kmhxaUYeCjP+
5YLG41UHMF2rWTN+yBGzmxhHKZKuPbTylIG57Bmh73qBAv58Mlg9kPHXKBR4NFLHWY5DwU8yArkV
LWLdBpi71ENBAn3FyXbCph41xchklRDTY9puzaVgglsxBNY9h5Pi0CO/Lh7VHbFR+Z+52idlULPI
FpEsmj80DxIeqxGhl/2fVpPH2Kc6MXfZ1/MbwYLLm/oKqjqVPPppHy7QC2OiLDdA7+xjXNHm5KDc
pX127JI7KdMx1psTrgO1b+qSm2oy4pwdlJDlvErGHTUHzv/x0oJyk7AS53BzCIWyVR+x6sF+nywB
hPR9JefNFIR1fbPvyi4vWwl+r9zSNPzqhVLcKmlwlO0AQcqdDwcmN9F4FO9xnO84YK+A7VdSUYDZ
BxO4CTc5QiiTOp0mkO+YjSVdr743OY9p1Zw89F2CXYkRIdvbXMaWkGwHjPbA2/gyIt/YJZicmOBi
ax8ABpGzZFzZzSlYxxRVBm/i7vBwgiOROm1pbbdM+htpXAnKtw9QnBdqQRiiyvoxVaj2BrS2Nlwr
08tM5CKG9nVFZ2QCej6fuGpptyYp+17zwHq19PUBYx/ToNe8QW3I2kzxD5KJBIJB6w5bTlitOFFy
SQZDDXBmn+c4+sClWP3pMSwDLwq4tPb03Yo/RtLP+u5qQxxFRXX7Jb6WXh9P14gFTxZDF+ynLI5g
nGcNoKIovjiXscRXemmPalqh7/ZpqQb+YyI7XUVLYg8VfIdDVXl6mPxIXkf21qx6VxheAqrNAbi9
hH5WQwicf9fidhQ+RHeMhSgyWSQ+cOovMKlSRQBSwdQ5vv0QxrBqwGGuOMbiZN6uIARTz79qVPmE
CAOLOTtKlJSrj1CBMhjic6BXQtzBREOlInIBykwKEM7Y5bI2yTqmfCL1QOh6v6/fPBxk3bI/dLUP
uSMXeeCnKKy3KD7uD342qp0VZrLH09Qj/BhSb4pq1o9rxdS64X82+Q5Tcc20yJkV7mC2l9TAuANQ
SQ1XL7Co0NmxDm9c+TPM6LCMDD4+BxwUo+QB8fq5Azhk81jiGkqDGceoAefOH5qrGzLi1sj5j13A
4JuCVK7H4AwFQlUCCCSc/eTaoip5oFETzcxbkgfToW0SnC0wWPkHS/8Gua4N8IgjQ2FS/y7+r8qy
kFZG1GPgQ8LFWhXIoHPxj4s8PrA2WeAVclq6k3WebbzRFA2Nw1lHGGHJNzPyUo/7D0FAfCAw4IwL
Fsg+ANtLR65Y3kEd+SVjDPZUpbs15i4qPj0APBMBDHhrJq1JU4g+OftTUwg0Rgvva/CiUpWAuKwc
HNVn/mCE6vGZDchjjqaFUGfUeUFdot/VtZ0kDxMxxX7OlhkFEVM2G2ga85eisbv8ycC2O0EdiCAs
bI++dpYfBTQ5BJZ+RA62DdiCKpl4QjFI8eWGlnI4KHt/tHs7BBALeSWl/NICOJLKyOCbKPwNNOVk
Z/QOem2EaO6L7CtFpQJ1D5oKy1k9xMi2uiA2yxn5voPv6ODzQ+OOE8yzy+rXX/kFx7uHkq5GIbX/
Yyfqc+dJToJlAMA0RdGaoaDm7diFH1yP6AXo/PU7YmS7N1kNGHLBzTPyzw/MxLXQE2KCbK0TL+V6
LCzBedkmeNNQVaqmOWiL9HortYcSTTb2jb3hAXYApmCK22xMzjKiJXSaIgGiDkA2VzICV6xn6mTm
hvgV3r2hsDXU7ghyY3SnIxKxCwBlZwSNWXTvknEpyTx41wAPF8WKe/vFxmVBzob7ylVlxZxyXqpG
p54ODugwSAKn5CSKk6W++Er+kPYWGWVHwwfmiY+GM2NlNy49uDydoqrl2jRQFXb6EjYD80boMvzS
DabAZa68A5OofnEbSNDf3764GnzEiy3qgCssgtad7YH/ysCaVZaxAp9/nVb8MmrOPbyuWXQXXT+z
uhPccCCHyRCxOpeKJVfUn6t20zsZoQUOfNM58LwmefPYqNsnzD1t4l+fq7c74Wk5qX40VPFtWz3D
fC2N+e4FbrKYqX+uu8gkSVlhvq2sND5LRo7bFM+0owMB9Q8Shy1hSmWTrN08Tmf6XijjAwlOunA2
hVvJdWS8qpeJtNUQhlj9YqcmWSAJ8DBgqSlIcaIjohUYYM5uK2HPID8ZfhkY1j1G9Lfs5SeHpbL6
i602XDwAJyblbmYqdcXg15dkttiBqxyGIaF9JhX4xygnFZuQQ8hceyPp+Y3Cx4pPMPRcsWduPwF6
DMn/YCuiaW1NWyH9H+VWUIsZC9mMcxS9tX8RRLnrANWSRkA4cV1kv4B4bPkBbgtO1GuWqIvO+N4U
FRZviICu7kgf4HYxX3lajnI40LYX89oQn/yl4hvMd0WWes/jzk5olVpL01X8p69/ftxl+nzk31rG
KHSv/ZaJgtUIe98w2eUYbZSMSq/bEzAHXwJ/7RwguTbT/MQ7HjZg9KPMqp3OKvduuyN4jB/yHRz4
R2PRPa7XaCg+ioiV61WlEgU399dDUhHc7CD9d7AvVDX9JpRMHW5w+cN19Ly15Z5M2EPmkjKguOCN
nIqFVVXESHnMJaiFRtqz6KGtdnxuMNGhf9e0u77uyfBuhbJ64SHQLduLZ2zxnWlo48JLMyDMdAwR
L8PVl53cOf++538L9o2Xnh0JNRgJQFvxowej6aqcO76+g4ZYbdumXqTEMLtFT+z0ATjhg2jAX3ht
EScp8xrXcWEv1ArsAYbJEd4GY9R4VSsOVNImkCf4eIlbCb3h0Hh3vmwg70K+jpfgn+NuVb7TJV0y
oMZodlqLSKnlKwf45XoqXfjxSRS0jQ4gc4Igf5ycpS6jBMV6PXmy5oASpN6EunAbTRSj50euNfGl
qHrNZxYxTN9tVzqvtmWqKd9Ea4MXhXg1PS/Q4BSMy+NpCgaXu8E0fTybYeO84uxZvaSZk+s8TCXJ
pyFHce6rvJS6Gqm5rSA0ebwWAiA4etv5BXm40nKn7HS2XM44ofcVTWTMiF8h4sHyVrl+fkutqwI2
yYt+JdT8pdM5m6F3GxbBzFqr+l+oRQuxGHcvwr9WMNhflT65vCQ3q0qxnZOjmxlHWYk+a5oJPxSm
Rfj9/Z9zj7kyL+roimCPmvhiKOjVzjIaUyBkWLm8yv2xSS1pt/rAoY2vuKjsdM9+JE0r0+ay9clw
awXDMbUp296HXhur6UzEVogvwewtL9W1l5RRizKjlr/55nZMpDpN5O05LrJ9blyXMSLjftr/AbX3
SiiL9P6675SjrxWGosLi/a+rOdAR6W8v8J753oQB+ZHENvIpGn1cVlq5t4zNB3/S/ovm2E6E58Nx
PQaLcytGIhM0vonqDfQDNIEd3E2b7K2ZzTpTNN4DoYUu/OPj3h0HhFVjjd/DgoTyYzV0gGrImv93
2G5vMVdNtZcLCqChrHl3DDxwLamJrAt93+bou4jPKQF730r+dlILJzrXH5YDIoVOkHfzcbybgKed
uq94fBohjNSXcQPU2A1Tt79CJFarJvehXi/dOaSbB738oCb2k4iEGzzOyowY10SAlZg2BeQq1MS6
L+GrkJYLUByJSEMaPgUskDDge7csNcqIxQhvytbstMd7T6O/QVBKjKoN0nLEiWlO+H8++6joISd0
S6fCuIRdsbn86tC223eznGGeSGZiUfVennj7VwLaowW6RfbCSYeH56AEE/nfepdXCO4Y8mmJSHI4
gpfQPqPyG0m+0SBBWaHA+230AazmqDNq9kqr17RrO6s8PDGMiui+5DdoVESH+dbppiSqISqnaDGt
QSU7XETNHHFBc3dy5oeizW9qcjbLXJOxtQic+wMPFIPGZzj6teGj+Q74La6bWy6kNW0lBohayJXh
vFC/7hAW/GPtMT7jPmCkwZ/F6QyF9wqasyDvl10LXo4cgBewwgim3h2CsYRvIDseqT3rP+M41W7G
eIE5189p2s27s+P2GYzDCsbR6BFdgEm0N0LQSdjMEzZzEqxGUe09BGwSqaE1pr4EXHyA2YIzjNED
5J9uumKC/owWi2ansjT/B0w+BJwcoJKMk+bSDiKxHWbPv9a2tS8tGkoq4zFXUbiht2E7ove2Lc5f
0HgUF2jSOV7TkfKdxVc5WsDjLhM92SWJRVMUiHKORudcwsgnr7ObJbc5+QNcOec0Pjiq3wRwoky9
VtLtX7YmoiS+ooKG0/dwXZ6KzY3bvnSEK0cjrpssxbRsBH30c6wrnFmf8Vpzix/dGoa6L2WRlOab
yFtwjyFtjhL+b/tQQwiTeNFLep0lkMcDUPkCXxKKGfUnyuj9FAvO9Gys2xqrcntsUI99Awe/wKHO
jL49adzZl85Md2HAkX37V86O0MjUVXvGNLTV4Wumq+8nmyhV6d7Ri0edydyMs9c1SdGMpawW3h7x
UirdWdjmLxk2UJmk9r+ppVJ0vLNl5MWpa8YTx+2qJJAzyDqKDpwv9kGX8+n7l0C2CGmDpf3Dtr4R
SSOpXikcpGhCYW3ArH3CEXNjl4WaUCceFJtPPnFIxL/MVWRXfbdktIFHYmCqNo584fk624mFHDbA
nuInSDolsRxyYycsf1u0XFyb/gZUOLZOwHRRPOTIZblREcya3XTEG3PmMX/WMWel6X+rlxSbwFF4
z7HUv/RjQEiOEPUsjiQlLKyLhxEveAO5UxF3PLt4sDWHiA1c+zbc/OPoE4pnb+EZW/K//io1e6Xb
jpXYgD0MoK46B1pq6gfJIPO2egn7enqrNq4Oe0QmGHyuaV8ga4uCxnDvS+MjNkHXF8xaKxXXFAge
lVQBAO2iOWReOjJunlL/Uvz8xmefqM9rU0Ob/JlVwdGisZlxvMWXA9nd5GGuYnmUPl+41b2M+qn7
SdQv1z446Oik6NTqrw5jt14eu7lXcwN9eZaYyVsBifALhbCTSvokJmuqImDQGcaAXocxmPyPFSto
SwfvbpKggznJbyoH61BI2QMIuvxn6jPMU578k5B8h4+Z35D8+4J28ispMvGh/OiecmA/DVP0yylF
pYetn4ZWmj4eswloSLORtu/CPRWykxh00CxttU3TNLU13gFmUIbSQHUG9vQRwOIay7ADAUOyxdlJ
e/m7ZfqRW4tJAqRhpBkdrvy1BizWI8MEV1KNE71SsRRe0FO4ben7XlM2j21aPijyYUcTHnN+R19G
Av0+OJGNUB5PUbsVz7sowoiEc+CAW3f513lfDH0dENTxy1Q00wbWJeDC1zgoIcAaptNBUkUBkxg0
3Kfu7AyEJPaMIP3A2EJompvThaBVCMaeImQT1ur8KlGri7qsb62xVV6CAp7HYZZLR+yOmjWPaRF6
jcE/0t+B0Shrv4DjyKj/Rm0gae3uglcASHcSeo/+oAhB04LWK4U8hb6gSVNoNUCLptAxJ79eDz/k
hyowGhXkC5LgoRorDBtxojmA2bovmWdsa37gdDGZB7knNxsydAWkCgUI7bNKplHpVlopH1ycD8eS
l1n36XTfIR0+9JmO/1tx+l1mV7ND42lV4MIXhDabMU2qx+7rTDJELFR3VUwKT1ViZzEsSGQT0/br
1taL1BO8rZlocPkwEjozvUkzaT0Vby192qbpyUQPvW/gccpKMD6hyefhECHT0dLttkU4ubkHrmUI
TxAY81MRKDLHFGcC98t/lbbIq8bwYls56d5tnXSardVTUSFA6D2vVk+1QTfgx8a4Z3hnmzuWhcym
86BSf8/bp/2zyd/MLFW2urcy9Hm0neyMtNcgQvTUKROoyqS6CdBhvCi1H/8xa6qwLhW3XACoHDLQ
XzH/aiHwHfblDBNX2Qv2c8X6lG3856STukYLybva9R6I43YFPo1mheu+gPPe+UfVhOC2GfDPk4qs
xUZGJ/dFWAmO3cmsi2/jLXpdR9DIDDZV7JOWWmv6GyoKuQaaiZtUG7qigmfREo/vQ7kaYIRxoII4
tzi/lulJZmup1k9K8be6pXm4cyb+rBptJm1ol5+v1irQR5x4gtGaZ+wawHXb3dQPTnE4pmCAsXRR
okUfFNDO+1ChlIl1SJMM2f/CKKOayZH/FlwVsIIDpHkMkcIaoFV8y49ZfwzGgD3OUaPKff8edoe8
4ZCIrYteL0jI6V4J05VJ7vfY+zI3Tweta+aqd3c+oEiBIYxFRhYa6o4IG+ubjnr2ktJDDcdmYlZP
jjpjkd5udf2NLR1GWVE4FgX1O/iZFwhqPKCGowbpcmaiJX09BfmEQKK6MJX59fOllwPUJdMQHcBO
VFzKujnvh+JS0B9Xxn4PzBtzDKFoijh8siYvn+1ljvOCcU8TlgtMVdFIH4EYrVCLaqlIgxgjh2+P
f/5Q2ia+UbloLwnBB3zY921DFE21CVaxTfMRUSJhKpxACHg1NBUH7uhD3vTCAde9IOtewwb08rK0
BUYsltTrclPYbUX9FlqMPpFPOfo0tIakLeD7U8tNVmAvPlvwXDElLXBo4nEEwehx1p3Y5ZecE0a+
HMYQdwg4vhfptnjO8QfNdVxELFhxsMSpwuBWIsmxRZkU1fERWGlJAdcT8BHWme5Gi9hkkwt9cvyL
m+bm+O1AfE+n9RhjNE1k1Hh7xEkWRlLrle2xjna1voMYpsJfeuhuXArbFMAVesHt5+4At0lIz+dl
SgYkssHN9LiFBRGzvdPNpGci8IrNi5iD4eW+jEr2MzVdMfZbmJDv+K4tMbr5Ymg63CTevBOykuaV
lT6n+41O8CYE0UO2FS6T4+wvUzTxsvds2U4acVKMWNVEZUCPdMx0/nrVrtM6D19sNwGX+ccLeqBs
YDQmtnnsCLfNMWPunH5g7H4rZLVNr6Ti5lu3H3QzvmMeUNRLivi/hyEjLim7DDPzUBQXji2g/fbr
zPE9vvLJU9mZPc5AaCn9l7lUgf1mhSpftI6Yowda4JrRL0XiRuBI5xyk+fu1JMjqPpBYwZ0SIee1
SMDZtsPjBwzoQlweQcTgTBcsFU6HkgpYPoDa2fBunViXaLZhEQliPVKkOE7WcswWgTw3telHDIJm
cVqkejr9pZd6eLtX3qpdTsz2CtVKJ8l/XTkpreLuhERG8LRckqwh8ZHBfc9VeerXKOvo+OGZs/qV
Ihz5AEhjP6V7C4sDadC3/Rips5wpV3GQVh17IyVex7zN3XXAImTVoU/bwx917f9fUJF59F5s1lXr
3Vpyi5+r6abap8o2q3P2RBkq5vdz2VilNDWxydEGW5+h/iph5hEpCeDkipxGSDwYD5Wl/jS27r7s
tGKw6G3+MmSAKIJqG2ktXhfbsLICqy3vJRUoLtpzmstig2gSK2+5rFTd0eD+s+u2s1/mvJgpbVsI
250RQ+HvGYENtl776Y8c1rYoowuJEHZ6YrRc2rSRZG2l5f55fSI7ovW7utR358AlW7f4TGAG1G5z
5zgVmkAb8pIGvizx27uCjJ7N1ZTpmT9+QPuXMQMMamc9He8sApU+O9i9trKQpvW2GfZVDjh747G3
JeUYTT6Cl+2N4SBLbdX5KxqMegNoaCK6VVaJJF/iiaO1zshUY6hhP4ZWVB73BmN8t28E886rqps+
Gg0HCD1JXr5P+dWjlV92qO5sc/tH5YASyAQwFhHnqhPEJgD2mAPPQv3hWmAnwZjnsxG3tnVQ564q
SZYVVBh58tJHcgor5iz8bkLXceK1nxl63lCcAlkQ5KXhrykEFTi7sCXshELqjCnXPpXSE3fhjCSH
5CZ64BZVAIqFLo3bMTpAG/aMANm0wN33dVIgorzfi2LlJj2QgFKqONISoqkF0XxImuZv6k3B9JZF
DEemODKI3wjWA6/jX11aJfEMM2hafSSbMtfPiqJ0A7izM3I0gE5ELnDvRkx++o4i3EQzBCUEqome
GlHAZdC8ibAdDQ/Uqe0G5zCPINUkEUbQLC8ypk0Frj9PjITZYFGXGJah/HNSkw2adWIbgHoUiKJr
y/fjoHIE5motgfRhRVMjkxeehaJeh6R7oOMEDhP8Os/YR7a5lcKS8RXA0/bYq/Cw2q22lBuR3Vgv
if+dt6XiPDws3WQ+/S8Ik3vsPvwTUqnni4nOyZY42MtAiN4vB012pjY7ogoi0cmIjujycjophGGK
crUh7a/tjZLu8WU0lLYHSc+Tr0jDg2rrf1c/csoBHz4eTykvsyJ6YPU/p1BXnN+L6RP2Iti2ypxG
48NazBPxFYrbW32cFBynY4OLKm0UdsrJ4ZoGLTfGVxtkwa4axAFFF+7Cu16Cxl9/sgthborfuzpo
k2ohP8h6xBFs7H+e1OpOFnfZw7Tkeb45sbAahvgJjEgNUWGRRbGhT5NA1Mv8cA2MZ8WJ3T8Jt/v6
gfJPCUuUrS9T/tptmsyXIrEPNHSxpCnUsPxv/y7lHtYI4KzakJ/IXKU1dBHW6qKan1r5wCxi/EAb
LPI49l2m7CUgWfwCAkcpwrVBXDfbjC9cV8UZStf8ROzAWtBnrOwSaUCbNvPfr4Jg9mVFN9Ka9DKk
6u+snfG86usM6SqnTM3nXvmSe0KLaOHRVHwrOCYxdYY1+82r2ssyGlATm8u1UkDOiaQ0jZl6TLUF
TOCjm43E+pr1VsmV4Z2py3AqDipchRO6krIlbOBP2/j7jQkst/lL6Hp9lUYLQVfSmETzDkJ3YzS8
7qKrfqnfoi2gMO/J4OGMkjfE71umXSB/lCR3AcCa8xbvylmzmEWHfQeWuB6zCIy03UGr2TYsbMtf
wzGr2nJyuFUMSrMkQxcoQ9pLfB7+4zagWFW2oKZZ9Culpib4tvAl/8HslhvtV10tOAkP4hB8RHbu
kLSgwcdlXRrBH+tnsKZVrAJ3CUQ8NnRaGm1tyfifM5PohJWoxRwUcXg1Kzh4dgjR9FMtO4XfP7P7
tnB2u/0aXVe52GgfBGXIiM+20iq7ymtEy+G0LJRsfDknai/5kuiVJ8VT5EdgBMG13oyvDQDSbKkh
P2r54198EKiy4kjCHI8NaD6cPhNusOpv9YFQqwJEp+QHeVNlNNhzwp/orJuCRVfOEqvW2eRf/Qv0
+3q+YoFiggrHi4fLejcjUlRABXIenSPFPIYuA4zdr5itivdzl3bxNywpeHErqgW8r00AeD3RvsvF
EU6igq47OU/xi6/G76h5jH7BWU5Y77grfCeID/dWudZDLScAkP+DPTF0+JThyCJ3wp+dkgiviDnf
z+nbka+0JHIPfDUcLj8EadzxxbH+wt1wmDaBZs4G9JvKA1oCGNEBzgCI6riCy3aNiF+aCrYbQbF4
RU4ZL5hjLYy59dlEfFuRSRFKZ0gT9IMkTTun3tT7JDyeU2x7oZ39siDta7iAghUJ5MqXdlLmgQBg
aKbmvxG7lS1+HxOyJ9cLzx3kal5vLWEk1myUkwNM2C1Ob5Pyt3+/bpHxidTuM+XbJrXVbfAVh/Sd
ZNtEw1M0rqfuV+wE4xxKoZm0ni3W5z+TlwRV+dLmhdE797Pza6xuC+dClZyUUFRwbOodDAmBYmvx
TamtPUtJ6x2FewSZNznh5IWkmnqCLIS2R07MtRjqDIf/GEEGtQjRoBuP9HpV3SgKHLt+Zd7nqdqd
2CDeu4e4nWURiaJN9tK3F2EkuGZ4xkOjFb/uuVgwNMQ6y73Qk03OuwYXfD/11zV49vxtnHDb0iFH
Ire2ieyxDx46oPJbV2Hr2Pprev9DAB8F9JNrU377rqNbjmp6D/gvva9mZF/L40GXFT/9PSs3twuh
4inklCsHxkrCwa6Ka9M9ELAsw3g/MIAEmfpWxb6RDmCPxF4rKUFodmGPsHV5nmcve+fZ/Td21kl+
3+4AWZ3/9pxfrOMjq+J/3NdT6PnGsDXiJeAZLPEI9VO5nXqbPgTVhfngOSHXcldXvGcQ/gLMQ0r/
wA+E3/i9aysl/Zdk4Da03qVvShyxg96c3uGyeFuREc8YvUbabgo0AQS5zHSWIAFDjyCZjU05c1Mr
uq+RgCMnAvP41DL5rD30KQJEBG21LWBotPsrPfloAKh0W93NyjtSv/rKHpqnQICkWyO1F6/GC+HV
IHt3p+uFXbtzDfeP2A0O5lqhwDXxHHI5cuItdqaC1vryYnB7v9SVgK8AgEyn1MvfryeE0mQH2Acp
rRC2vdO9bXoIIT3zX2l4U5Lm3nXxBgOG8CuNiybVplPbXlvimtp23twscB24vdJew6kS1P3uRch2
JMNRNu0HtQnZCQuUI/Morn6efBFUSrNWYnEVKWqNIPLs9moi2AT5AXsQ/i6sVOgs6P73k2zB7RE/
VwY8gf/wYRj6IcSonvVwOgxrvSe5P1LVLYvJfZ6na3A+CpIfx/N+T8IThFMQVmNws/UrXqjRAS6E
WRP1u/BlzAIapdfDRZfYQIQywMSldCOM2lahfBpHluBlzY+4e8X9qbE3Vnt5aH5pyAouFNOcq5LH
Ve2ar8QsVB31xtjxLrLXj52a54lGhTliVnno/YLDqeZu59jB/Fr2itomdr0N2puZ6vJLskOMAN/5
aNjq6rcZxHd9s5XkRyIxD879dCzp0PU2LDh+Lq4ksWGrJrIEO4rcdS1E/B4uHK/OuV1oQI5ZBYkf
59Sx/tYjOaX4BpgbtyWSAm/qz3bb4WpJYU64LvToC+mXT+ZlIj7glcSi44OC4lBQ3TXZWBXf5v6V
RrU7GUQ9pJixvQl2IFmqcrdZkRJsf6VG7gXeNKBobS4dJ7xOLLMCBjEoIjDitjA4GGnR/LYqL5kH
l28Kwbo3q0JX9Ow9P4B5IptTpxdye9LtNZoiBVQ3xxgj9BEC9dJtmKy7LMmMCRZ9OsAwY/N+mF2y
wgNi75JfEtIZssZm7O7s+EHpHF9TjRH+TjEuvTRfwUCHiR8FIig5M4eZUJVWOTrtePUeT0I7OlnX
SeGcLw07l9u4M1q+AfLQnH5NpBjOuy35wcoAF21IXd6AS0x0UJpX3pQBIgvEef0NxUMtd8XQU+Z+
K0nwGjqqUfZgY4t54lyuhkPj5XA/xOfdkSUJ4kg7mLK4rxoPo3FhIdyxKl+8/pkgDza32VqguTPE
Zu/9gvot96Ob0PoaLqT4YfTz902wjDPW5KiCednFVpNSXzIc8g0/2+B9PZGBbkJM3h6F2Hk9C6uP
agud0X9d+Z3T1vcnJ4CF6GQYH7cTZ6bdtkrQYNbtk47b9k1b0CJBQ5HItMErlW5mJe33jYOKq8cT
FgVFpUxovp0PrfhXG1zioZph758OryJwKFbEBL9IpWNiz66mAC7l56fK5KG8aiFdLh9ooQQsMdjh
0CnAxziTJ/tMyjQqeXWbabomccj8HnPEWQ/3mSEHryuvsjAlthnjZ2a/0Gvtk84ExL6CbvhID44F
ijjqqQZtjmFOFbyAKyNXRcuHepSGXkD+RZz0yLEP6TaojDYPpDPQo+E7auT2SxUYT8JPRnzZcbg/
v+lFGdr24ZvI+Ab8dA022QnGYb5mTqHOPd1M72h9H+IhPSUS+tWvOOukkdKtSlSiDvjGVUQJ3KGB
5nYoDwcjdVAwmEZKqCmCqyZ51D/MjR0z0NeS904N24JtrL3uOi/Q1eUFyBExold4iQYBSoe2YKDZ
yAxJQmIo5UyqDzmDbEdu6KnTU3DbbNJJ60zvQvZ3UvB4YqtaN97DF55RosJwA930kXoibSbAMqVX
3+CjZ8k/BfsaIijQiB01KMjxmnwNX8rShqJLZrsWFrvEyDEnybVYhjG0Ir8XTZ1+WiNfagr6KCj8
ygfXB7Pnj9zfVKHwCaXhlav5afKEdE4RBjVxOZD0DGm8apsedG5eMvtzna7Ki8Jud98ldTEhlzhG
YOieR0ZztEe5vD97YKbomYoGT4Lw0fsL3HqdaR1hjUBewxir/e2WMe6/2GsGtWleNUcfqA1vhiLx
HyHXhU9dpfRmP9h8fvb1gfM+hwC2kSidR8MacoTGNTobXx90r6k8Gin7/qbrOGM0ZMA9B+bF6e64
5Gt+TpQKy6Bzc/4jSu8WMQ19TF3pJZ7g+jU3rdPZiakQ5j7PXcpZGUBKV7SU+jPmdjTwEUeXqIY3
qhn7wm+VPc7o76iroiPRAmnTSMijbToadMScZ70egM1CfAYKnj3En5ZRMORfwId0uKaQrcJbhjmt
Ip8Mqzw/96HvdxcTBuMgnjyWEixQoBXp337TGh4Sg/RjycHCosUsZPCWkrP34FaI+Zl+hj9hUmT2
UDtK6szQIvjeYrJtqVXmP9rIxUaBTtlq4tYjwWRJotQ+OWVRQjTE51AaapgmCFooCnWAVfRpgTW0
s/CXzOiUjZOAtFINXP+O8t/CpZc6+8EMSs6W/qx6Ixjond5ELRo3PgVCpm96cGnxsk/ZpNLcbGfq
emKS5vuqZWaeBtJHzbr88Gwu1Tm2CbHxtBAG36Wx+Ld1Bg9JAURKbQy/e2OLioKWw1jKmTIhSwIr
xUAFWDQG1TAbbez2VUVShM/tuiyujiEMpEJUwMXGrdwd2n/G6mb4O+qgFK9P2yD2r6yMI6zUETtt
aQBsxGj9j0eCHvsjsQUw8hO5bD2g/9YOwlgbrdTYOR3OGKyEYSA+jIvPfcL02MhI1g4w/zAM+ArQ
fgUR3WvD+eVGjqbcXFeu3FftdWwuWydhwN1n7LTeFMiEEfVCBzpVsFkIR84dvRN41PzzDk2pX17Z
j6mPRwvR3mAKHKBf0dHjAaw9nqklMw7lm14dsDSSxBo3o6gvpZ3nvv1ZHMy1CnnfsqYOfzfS0Vbt
15Kz9NBc81TCHgErpmGiz4PnBBd9oBks11BQdPAh0VDWsag3eaxZGlS8LxboguPT17cMRRoJlE8z
WOLpPKVIx7Z7HW93Y0LGuzcq+FRhKkSCzK+EpRnLo0O5x81O5BYv3F2b6H2+oz7LQ+IHPUMH91nx
jX4zdq+EJr02mHwYjGdOvhpElr/wXDhtG+jUSHQxHHp+2zszGEyZVVqBQBs5y4yRrIEMfYNKFQo1
rIfZC3mWKJj9FaHlkSl2Wdo28sjrkqK28YGpzirn612sA7GyCDzKvUtTwv2A+EuXvWbCRXOFNRB9
QitSWZu9j6Tm16oIAkyltktlmPQIh3vBtlgv9SRb5dlTkCjJeDs/tnFikNfd336ldsP3JtjkfFxQ
luavTqlgOm1Gkxtfq5ixNHdmVddG2cybP4n92iW2ryOoT/1cE50MQCwAn4rkHS1DGJd6bR1HMIFz
le+xCesVefRIVA+t2OWgRsxTP24Lj6PvoNHZMCrvaHogrZiX1A2vdUWw7kUquT23RkkWIDcsfW3r
jUDZlvGntnmAAMGbaEr+zYpjeSiHNkENk4mi0N6l+TcKAI5oX92uq+B3YXg5evvlggOEtBcKCr2O
f6Ey5eiS3qa4tY92yiEhsTWujHygoh9gfJ5biVTWndvJLjLJkTclnNG/eNCUfOUVWKM8nQTDpq00
CMU2UnAKa2ti6BdyAZSDgRX9sYn7LfpL4xUreoW5hIIgkihj+5m8q+uy8ENINNucrgiHqAkqaa6+
/dSAgl2zxGSxevqzJcd5UMOXkzXiErt2mzLyZDbMOTJ6ZxP1sdtb+QnojgFmtnD+Mm91sZTjW/0+
hqOq9wPG8UTsGICjCLYm7RIiYTr2Jx44shC+LExpxXFJazXW+CphqCZ5WBo/XGWkJ29IA4HJQzQe
36xLp7nGRoDIkgiOQe/xscYHh+6UjxNLaUqCbUfJ68IWUtE+uLYzlndmCK9yd7UX3HMhUFWIHWWC
PaOPWNe0KZgpIeS2Kz7xeEBLmCSVluL5mDCI68HVcanizso1/csr/bq0mThr7S+3QaYBu1EutaWE
hqNoLUm8r1YjA8vHBu8tb2B7adIJIzwWbAeJxFrcGgmuXCtjJmX89UxarXmoHa2VM0sKO21yr/0s
9Rkte+wbXgnBJDwOSv2WsL8dlSQWRITUGBDok2IM7M3FiJQUYJwcLcfxl76wwPQlLnYwrKdvUVk/
e1hO4lHkNGpDpMN4d05zAYOnta398SvyVkOmRVqbl48ssllxI8q60Zf+SJjGbGU1Qr5QSUXUKy35
TPKbPA0l1sa1L4CtsmZJvUFlHa20cM9jmerPoJljloxB/LeS7T7f2byzWPxzepqxTU5eQQVGHOLh
T7oSzeD8FS3F4gJN3I5mCfV7Arev1Ho5ZDKvj6PGP1mIRVEd2gfIv2mzSz0Dp+Aq27JfnzI2hO7u
f5AY2/weUSgZIAecHWXK2HfNoCD/JCl/OVHIu9/nvJ14kvykcT2VV9h/98sn9Y4n/TitWihy/59i
yzcDE2138XFFCdnKrr7rzFuTc0KlpuZRkDVTTV1PXmIitRBdnseGFxa3qodg0bAfvkFYGi6I4STV
7d2kH751N7MzPjbzQAQ1xRq94lrVgHVmFvs9ufxe6BkZ4mahr3zBqIQql1I8KX99QO2DagCn7p0M
bSJ+WeTT/6qcnGiSZf+6wEbwbmhIHqF717QOswHJLYHInEQwXVPzFN5pmlmN9r/oZDrFPpebBum6
kBeyu5FTRZAGIsUnz2+ACDUUt8KyArQVV1w0o5bPn/okcHGFPkQbOpZIUXweiPB4YXB62li0iySy
mShMlowmmVxvRBXAm74vDZ6MVbf1MizlPUEpQU1CADM5B3HSsLQzToZYvO7FCDDQoiWXv+nBc5lD
Yf6s3H0riF2zP8SNqs9388wdN/XLqq3FQqu3rJW5/dKwjFhtInaxlCrBUK0atIyw9UgoPbCdaNii
uj9udU4aCqG9DZQh2uYOY9kPCmr5YUvktx4IXLrD5f7P6SoHP1U3IERD4NAh07SArMFQxIF2b53y
Go7830uu69tsb/tlNM7u412qd7MU3F2VOfFeFbfTQ4GwQINsW9qgty017rWTK1Cda6piSa5cflsJ
uQO3xP8AbyAVAdjptTwEIMtfPZp7Ewxgp7/CfkvSUCF83tRgpjDemoCaxjwAq8ejs9tu6zATdaR0
PVGqDtt4dukBcYNgU2SBOt4ubwdcy+gxXZ+yVhc6dwtfflCeHNmMuqsw3iNNMC2dKQnSW9PfqbdF
/eXC0eJTfrFp498FC4cNT+j3HhCLbVX13Jn2ta5tn0Qk0J0dC9Ph4EneZuDSkam/AHCNyLz7bJla
CBrfs0jvRxQMCyhhgx6DqgHjb7+gpXhlhwFZ0FE8zIL6/oYyQPVvl0MMJU5A8V7hHlpVWgCUYcuU
XbvUXiomOGxnFD6KHwl4/9KHRswH1+cUnFVI7FL0yE887gpJ25ueA4VlOFcR6NTADymsTt7ZxDz2
fSpLibRvHoOnmX8qP2j88bgIhHRqnmZjqS65vbyxY9/7P0vAw1f5oRCpgU6J3HywwutC/wFAUyo5
9aef7CX/zRzdkm5Z/BBTDGSKE46cNds+txLNkbFvjtKLCCrRbX+WDJjK8EWJFeq+fbv+zor/kZH3
1qBE5WSmvj/hfAM9GsoCgNfgj3yU6GkISQo6mb+Yna/gOfJdyA7GUeHyMBllVY3lGFguztj1WN3J
DHQIHLncC8WsAJic9MqJv0xAqRFN3ho53dL9WjZg1s4tmZ+h9AeLMTE/jBxsSxU7Gcezq8U4+U0Z
SqdzFSun0bKJ4BoFd7GqsI0ajJULxMYkRZ1lBZgvqt9trZU0NRBokWNU9r/50TxSDak3QGqa8wxd
6OEYvry7v7I+myryYrZq2jQtL/AyDRv7i5rZN6aqdCL0swrWdNIFq6htYYNMiG2Fs5BPGXUlHeah
TcAn7NoiDf4plu4rYdOSEbPNpDK4w2+HiJiTLNCkkw7O5liVQRiKnLUFSDWDkIz4HQE1PM1jtnI3
oiHfV67tiQwzlhAFK3TWuRToHtcTkDROi5mbf4LG693uaqdKh4L94uCxHrJOMcUg9RgnAMsqfC5J
0dbcQlTaIoI5zyY7zvwYQPiS8jRzmCOg//DGylFC1EvDE1xaoJv+em+sWRv1vYhTbmYeA3ywKWGD
DAA3O0xZ3mIAXSXODUKhPrYfmo4Ft+idr4Bx2tuc5OlC4QkdPADAXY3RObk2sZh4hCJwWozzFi88
AAMkgROabsBYxXbjAz7f/DummZbdwkkmL5OU5XHCece5rzN12Mc2AcwkscL/KT23QGS4x/TcnRvw
4mu41U68qwHnNbjBtRF/66/LSZHY4Fz3nT83Ogj0/wsAYEUUYoTA3oSwSyypJ18tnV0Vuzme+hWu
dz/ss+epihLT/uvuSYFTdo/cK1QC2IKu828o9tnxeFb3Isf5PV4i5iDefkKGEUT8g46wulTw6MOW
VPAaQw8FEGYpHRBcW2IrMAtXuzTUa9u2QGsFnSKeU12mQwZmGvjGFVRISXzYjbFj98dIL8WtSaIf
P3or1bfl26Mpk6HX8jMSWSDGviNyHUvtXovyw7i+UJHvQOo9eVP34+WTx5f8kd3BjMEqULCb2Zss
ZTFhs/esN24ddf9MZsmPpqHgGGMtOsCNVZkFSGCkiBSp3dcd1Cl1DBFyTUKtY1ODlZz/tOnaUAqM
4kmc5CifJZb5GFnIEsrszF5QJfNkIw9HzrkvpAa1ukkVHObuij6PclTt9BVi1VSH9kZY+pLnrAkj
eXfl/yOEJa8zaqy+//kH2cEEe4rPmHyKM413/mEVzbDngRcIZKTs6P0853hz8P+JlYRh7d45VcO9
rxhQDM/WAD5Qj9dZME7371an8FC4hk7aoHWqHl4h7FR0L7c4WP6GAWe9RBaMNtapz/Apm4HEGji8
PLJeQbT81+6/e0WxbDy7n7rW7rMhPfvz8y/xhd/RkQ8dwLB6eCWZKaQAPEs6YKmEZCSN/cQvx3Px
RK5CkUTnYlzNneiXHeuO+f5CTg5gBYLf8YBcT49TgJD4Bn/CEjh3rforgjxDiRrBu8W1+7N70+Es
Os2u5iZoAlOyZMSrEBPRqEq+bcUkakl+P24z5MYLAYyW6sdsW1sd7yZVdfPrO0MUvc594pl0KJjA
JgaD51zBeGsw1k5ZjPdNMK+aGJ7333w1+5Kdf3p73hKvWKDQaJnhF5ZtT/fNAECSdNDsotcwY9g6
+kkp+aJu9m7uYxSbPocCxy4dit1RYgvG1FpKNMUwtcivoLpUS4ORgP7caGZ9Zw9vlTMN4HFNmV+4
UWj2oHnvoJpn6vqc9bpgIRhHgxxT8CHOyzBQ7lp6jE22iXB+HlXz8EfMChenFPLp/05l0DiZEG5P
/KYGMUZBUec3kSluhiHUH62kzoWda3mXqwHlb3ZKQARnjcKdm6bp0GYPgaZ8rf4weTJYzAGaue1X
076L//X73a3EXfKPonRA8fuGwMjk5/czXuy2+YsYL7ENvZQA4aUemN2bNgLlq0N6j3qmPcI/YOsY
q4nDGCm3ba0g5S2KhmyBynGeEcEa9nmxzu7l/xYX6t4dOwAeI9b/tXHqTyCaTmFTGwP9VK5sjKxf
h6ldKWS5EPDx71ZuLXgJe8m8TcUbODqu/sN8o7grevOfJhNXhGxXFc7ujKijpXrWIHtdHz2KXKOA
z+pHT4MkHVCVzhtfHWuiVbNSoF2bT5XGueoFbkQm0kEY95CrVg1wB9+jeRnFPkEPEJoX1YGdGDyq
BBHV5WEqwSXfMVzZvBPsq6oJ1m3Yes2og0tsKy6Aq9axX3WGm97l+Svc58l/OFOW3JPCQ80K4G8K
5glrVjEYvR/cJaPtiujbRL+IzT+JFmgpMWmr1B2/Eq1Alm1aYwYRS7q0tWZvhQV3Ugy0Dy2Y0vAx
ck9++AG22ZxulIfaIGBxanrw3YITTPx9sJNC4iLzSki8CLrpj6/I1Ny9cuyckaG7tx4/Zx5+Vx+x
qiTatXOcNMthINjSBpP9pSDHUkoqh191Dwye2Ik7+N+4Ky1G9krc1zz2RF+6+bVWw7OI2vQpN2CJ
buYgGodvUNtmwHYE+K6x5X8GxhgO21NLjiQFrsh1MY2+EYO6p8nYU5yT+Bt9QjmN+d09szDH3LMT
vH6Csqa8zy1qgZ4FlnIDhEF0RMjYRCJAguZhiHC20xStXOMpS+k0tUctz8xuWy6thcucMOjMP9my
5m6lus0cGeHzofsedv+Uk1rHbVQKKwNZZkuLfnD4f7zPhObRfETiKpESL8WKMi2TtzZqafglGvD6
GdTkAyS5geLleIdlWbUqoymq5/AzEX7xNKzcPF6amhpJ53LLPtatKSC8B0IUgLkZvGxcU/0MjHTP
GN1ZaRGz3Am9gMA5usO8y7FJb9OvNCYQv7FUe/6xbPArEFmwy0+46ipg9HFXNUChFK3jrz+d4MpE
2cuMRXjTtdyevN0HDTFcRhmwJgiqAy/9lRuedesikb9YYXqMMJwhxXV9KlHpXC/YabOG7V1cCTM3
muNxIsX00mNS0XlwGctTNvU922q3FQmduUTnmIr0DwPkAmPc7aWuSflwopLWTm+SAQpcUIesmDja
hEXxUORkwins1hkl/EQVtEAD4RpnITYs+U1GK9uhbDf+nglAXeZG03j112TZvLuSiCH8gDeBO/kM
sDn4NYjEa5lG/x7Ct+Ajc4sP3WpoVO4iC8X9n0h+zsPtPbNXqDeqKrAYZjgaeJfzq0y/fxcZxrSk
XsRwNyeqZNVGwy4kSq/S8rX+6CGHghQiBYSnSHT/uClAB4ncK5RsVP8ThTtLOFbJ02ijFtjKEIlu
DQANYVBzVq8G/YIIk2oCKHv0oILstRWC5nWMRuiJej3DVUTfEPmw9eU1D8nuBw/EwXd3qWn5ncGo
bkmozSEOwWkqvyf2+7lNJOt0EJRLm15zLYOa46KrsUOafqGIjYfCAhE8po8ZHEECCbPBYI0UJF4h
v/8UjHLjFwazWazb8cC4mxdQEVJEdfaL//bz5gn6skXc6l+9N+hLYTspWML20h14vAxWfW6UecSK
r75Dlkytc1iIiTFs4FKPYv0ymYW+J7kI8GaU4rJX2iLNveBcWNh9GCxTwi5FN8fl83Te0UC+f8Zj
aGZ9IEoxEI1ulb3S8Oj0dTG147O7tgSis3pYlK0ZhFY/3TQQt2K3+0vRjJlyHWK2RgiUcqszWPwi
jLg9YnKuYJdPZkEYzHtxWluwR0FOP/bz5BPpC7A/KP5+aebUUyvmdvEOTCwaLGTNTcZQqthlwRuo
zQBSG/jh7TXjADZP/lCjyazPu6nNkT5N9pLfnq9YzHOZfqN8Nsimek9tVHpzCORdG/NpDMJkasoJ
DxCXJbSHJG2nCyXT4VysLMM5WF1dVimPCjVqMSo5YYYchCqlIBqMxkU1IZOdgSwHQONeWkPu04J+
Kb2xuTMDpi4mvck3E7rk8g4hzJOxIUigK6Z/B9+uUFua9PwX3ZN0TNm7NO493xuQ259XcIbOPwtY
IaVpO+4QsZItcajxtLMLZRCA2KGQPBT+zpq/VtNtfU6f3HiOAtI9wTu3OIbyYyYroyLiPlTPaKqR
lejpZSb0NxTbZ20MKxsYaMgIee+wye1RFdIqCJakmEfN9rLIq4KdVlQNnb+L8ZJR/rK2/ley2bQ9
hmRUZgP/uhDPOUx3N3c6qtW+Esp4ugEwFsVHE3s6Htwqlj7szaa2HZA3Jg+BdUK07rGqhjv/y+HC
9O+5wClbszzkYATgH9X282zws+1KiHf0mFWcwtlddsQphVi5RFo1dpHqcAk35BMPzkV1Z1eT+xO/
kTetmP8IsZl6CjdO9MC7t8Fu71xDNOsKuJhh3zcTD1nrHtla5VmbTJ+8Z57krwQKp+5rUcxW1VJ3
V2boWwsCH8+tez1kne6uffvchFQ/h2coQdgXrl+5s7L/kc9+ZGH6t1cCtfv4/7MWOKuJqyHc2+Uf
xz8R/9eY9JptRrsi+oT/+QcHXtHH/wCkWA8bVP202MpoFDqAi6pz/tU4qq/qO1NnaCKQGOtFOs/p
xGbQAjP62SnkHw2ZF/uAAm3TzTDj6nmj241fJa25bJ8p/mvXhC6nObIPerELciDf8xecHx2o53DW
3nBvv8yGjPD33HqoSE9OUU+v6tfrtx6lQvxMy+feI9Armk0DfT/HrdzLUBzJAFjO63bnm+Q9y8UD
okSRN8VuQkZt/0ne18WcyD65LT/Ab4TyBNB5FK2kWBVY+pZpqZZCVI5BG5fsUGHKWpEJ6SVuJlRD
e7cy3Rm6fFjXV1kfWikG3B2QxnY4Pv8G8++8ELC2BZpEb3/WWT68NnVZsxV6D5ycNgEVzkSRSDzF
BSi9qAMImnSH8Vk2KE+zKAieSOcQseTE8F5VERByPx7k6qKPONhFFUiUcWyLbW4NvMnc1/Q1Lc0N
oboBGmAuGbh9wOW/Uk3guzrjgadOx7F6hYrm4JBFQ/6EsG3mviK9O9aNqiBaq4bxipC/WPmAUeiY
eTTWFMoOAdNnLDECPRd7hOlSJPzFJX+muNFLFD7Ipxm1RB2B5oWnAeJw/Fpnd1NVLZYFbBQ8xj9z
GMfYFahaEtrx4oNF19MjUmacqF2H+p8IbEhLMb555nvmVY94e1Zgs/BuY2rZ8zQ4rRfRusAWOJhf
jObk5nZNcegKcnHauMkEGgkCVJFsg44fBqtekYcRIIsSBKF6PAPCZTmU1ArK+y7d2dgyPLyoqfV8
HqJQ+KTd5KBt6OGjJWCnJ/xagt6ARRtNk8YjacD+0pRNLa7/OraZxRwE5F0Ji8dqVh7yDfWzIVWr
zXrP/NCsWLDbtUtzoDUlQ5luJ0CJokB0IeanngwHlIh/StwumPJ5BThvDXf0RuSyr46iaDkVD3S0
iUr6qjYK8YbwdTOlCgpQtCAcidYabvBFpqGnGtsYuRQjSgseyBbFovJ5Zpf5PFDgk3VyybwZW/OF
vbBz8ALUEWi2EpkeWuXyCiNVzwnVwD6AihHJU1PRrpNXpI2gu8Qh15fbp2U8y+xSvLXmGm7BA1M1
eQwCcpwmI+qaJGxB3bKMM8QrhAHFAJLyrmr+EaOivRWK9PZAFylDtaV7KvNxezkc5VBZusWaeevt
DzEMci5mcWN95tmJcuskWq04b790FuVzhfI0b1AutYncPFU+lst67SqqOs94o4ph/M8oFhH7Ioyo
/CXJhhQL5CtJASn4pQYkHwEBIAWdOJ1WYU5h9gFfRE4Rs8/v+6xh4aX44KSIrFBmNE7yGu8Jphpw
lzu7sxJYkZsBub/La3baJquxOD8rQ0+QRl49o7THJ06/jgOlZGQTOrgPB37EDnsPHg3cdXJxtdXd
LSDcOAngCBFukaIWARiFgmmLJPQ2bJ2MRAipwYIgHjEMMMNQlt49rPUPPqldt3I1DrAeXEPPvu5J
Czeunaxizs7I4LidqUgqYFc6zUTL0IzvLbucRbhPWHknOtqLWQQWecXUtDlnOrmwsCKeyS8fPV5s
RjgQZtWvoZtVlTtd63HAR6iA7VFOY0awqVW5WNxPxagZtT3UMxJiPdipQdGvQNalwrvBffVtoYev
49fSN/bZH7K6oPcP8kAJyzAYMd9emavYjWLvsYEU/kNjyyNZu04hcjJ0KURXJFffAq+OwfMAtEr6
b74kaPbUtpXkpgK6eiBy6GWav8vD7ActBia7LQE+egJPkStILJzA5QLGykvHJrmJDXM3y/mUZiu7
ggjAcfYbaY+PoqI5Qq9fYHEWvj6axUhU5CvEjxzOcVVrv0gEpywGYeFH4DP+XfQ4R8OyJ0HBGdbe
8Wzg/NrJ2Lk4NedRxZNas3jUYx/hfZYJhzOaqQbUlVUE2cXclVmiJ5rVZp0suMd/PhEbOWg0UQgN
x+2GtOQeinXcT5G/4ankUu9rZJeUYt1zdkP7fY2weovgdRr3XZsu4u7fLhTcRpiuz5YJAZIkPAfx
oVaoGwqsAbehzhrRe5BAKVPpqk4lalShTJ8aN/e8TGK+NkJI4lzGX9qggrhXoDkKJO/v6O6llqSD
CO04xt7BVefIqzCQ1CLglP4HvgOui85wtNzz++4R1RvgNaX27SpYy2ba/W3TdiIRV4OwrULNc+Cn
7lypQaKy88h/VdB52DsxZ2Ul4RtPpPdL4wC3OXsA0IiGf9+e5aOInfsJEeoCLRfsmluF+f4k5oIp
oPVVo3vGA5uF7d+QiP3nsEFt7pbkpDUR3ZNZKeTloYEQQ3uU49jhnRW7zOQJd3zJkj4bC0CsWm0G
NGNlqVlHki0blMHEF5+53PNmf/iCKskXtYx3TiIw+J3pfj7XiKGEEHywG+xmNAc73JMP7ToJKC2W
tfoeoaPutcN+XfM/ffLEdIriAlnLcMq1+k5UHT6nrjd3tn9u46zRxCkw5TDUAXxJoruLbz4qhk5I
SEGuZygfGWPVJSTHPxEiSHi5gQhuFA7KuJRmRSEh9TuJ05zZyr+VxiPa+ownpwYK/p4mNBEfYUhW
wO/fw7PiE7+ffqlalVvLYuKnMEgOZFEqn++BqwFSV3tRuJtp3mo7ssb2LpGku3YArn8r+GvFGYJ6
CjPJqJNEvOqNeY0egoTx/8usFjKrFw3NLUMxi2NDQtNyZF3Mn1/sP69TZT3y/C89DsDQUJnuOZcQ
1IFDBI25zfTuRlZb/GOYxGSF1lmnu/kI6WLuFrqgKpiZ7be37QuAO7l4xRnh1g1OT8TupGGnNj0P
VNShGJv0ceRYxEKSm8yrE9h64An1So/auifjDEqvrsb919bOuMgg1M5q8E/KJhGqZZIRmasyqWe1
s91ilMWcP2ZewRYS8BzskHUn3SVmnYDIYNpViF7kk0+7uNByVgN4GOI22Zeve7kZyyxQecos29ej
QEn5xgc7GOyILl7oed5Nuay58ro9bx2UH5lbu8qZnJykcgryAAdA+YUi1DPyMZgPbRmsleWKnTPx
b5w3I/nzSEz83hhUGYp0xZN9KffxZBIhb74iUqXyzZXgfkPNhhBun5zic9fKJHP1EOuBYXEfb85F
bATkQPf4UVv2o3VszTvw0Y77Tub6odZXqtG9bm96wN95cNnru8PLwxplozUq7S3jGLcHcZwhSLnM
UOsRo6bP83vAKedIQ8vx9w9+xeNi3/NVEeoFyvv6LdpQ7DdhG3z1BdMHVutQHmw80S8uJ05LisZ6
qltg6X7JClgSD/9gIBROUprwjnZBjbIWl9qkcZ4tgQkLwoelFv1/R8FX4nRS3T2lWWKes08F3koN
JpgWL69CGvf4Jnide/Ro2mcMcliJS+EfVn5PFW0ckLYXWneEeHzkwjnV1lIjf7WleXMcuj4UEgCf
sUNbrszv539FdHnCCv1KnRZFVXj1mbPG9t0Sg0JEN2x1y2DM07H7xuIpmCkRU//E2fKvraFARIQC
zRSA2oIyFt6kKJKTL/skrHy1rhNBKss6ul8nPTxf3KhnhGDcoQSQtriCiMSqJ/y/yxlXIc+yRMpB
ze7qi5g78ZvBX6sNKtVScmwAtY0DfJ7GjzvKZ64kxoBMkEJb3i9T44XTctADzPJJz666Wrj/e6NU
IOTZOAXs0lMluB5+SydQ7FAuxcuhH3uQWYsn/tgRPT8cVZLukaeaTHCQCAo+1L5HQTJEfDTTc6Tr
vN2EkYI+0RNgJ/c1/PaWfxRpzcz7qlTxKhSmJQafSbIcRAerZweUhH2+UaTEqSslHXikmIcx0wOa
Irnc8aUUYiyYHg1M24uCtQKNb9aZ7h0UuzoHW5finSdGFoXqUYl2SSUR2HHGNMBzJln9sWlfE9LX
O1wXwWJwcUKqfJKzWTkYpY60EPuNJAsx/Lyg9k8sdeZ7T7BdiXyqaWWTxz04V76JzwhnjBCy2d/A
hx5Bb0o4l95tPD389wKscf15g4Njsuj99lJV5kBNp7J3LqTjkc2HOpPvbZFLovFMtsoaToeiwup7
PqNsCedwmm+3//Zn8QK/l9T17s4jKTzSj2/lRQXhAxasczDmLVwRjf8yDDWINitdnlV7HXN8GkXe
G/i0f9r7IivYt2r1waXPvUsMO2VNZe2PNmFw5o6tctSQlGY3AKgpq8jttQZJtaizeGiCtVqC+ImN
rdTvTf+DN72im2oJlD/s3dcj/8/DDmmiKu/0eK0DOBEFqGuCuyJNoVnztopjKwgYTgQdd9ZNViLN
izx+gx3PZIABzDUKxGe9KjWjKxKs/8S+9M0emh5V5DBpJ6lQO942GQjG/xuBAROw0Z+vP2DHHRjf
UzzRS+2vHsaL8PBeVuXY5J3bPgWLAoDNEPwLrjB3QSdozxQECX1RPJQ0ksd04+1T2WI3lFi17LX/
Fb2otPMt709QfiGSkLSc9bn8ReWHvPNnFs9rgv97ajBSBkKYOsQkokfsxEjMQLsavbcdRwxgu/R/
E0DV2yQtKa+JGvwE2ktW5FWYewXXx9AZuOMZdQ/HQyMrUNynHrJ+YaVGyteemI/5zk1Kr3+twH44
EiOxq45t/G889Vlg5Gl12zpJR6PkZortVGmsntLVKjTRENzkD4IvZS05KmsqoE7LBpD/qSLc9Lli
csT/UWXgL40aPYHgZlOrtawFQcbwr3d3hEL569wHhNB3+cFIll2KGhPqzZQhTIiHXjnkrfJpTffe
GhNuPiIXlh5SgLT3KIIWTNz70W98WOs15q3OSKQhsspsq6QcxHD9uOEv1JBEuPMrVRJUXrZYYMjf
RHXidQBeQArVz4ebmsTLGbiqjO+N+hmtb2VttzZmVSGruwgXzGOK+ssdiSlLtaxJVMbuaaL2QrKv
As3vxkHmB3n6nPL/tee5vnmCoz4ZUWqPHhuRl5X3G5v8dySjhNLJIFGaTRBR/vG8rPK4+xFUSF0p
yQbDmMrOPBVjmqOkPevmdrTKxkoYSuF/+ZSrpyLfZmJYjkDTJpkfCGU3BsoNuLpwqBUaMOOQkH6t
HQRqcwWfgRLGf1Ip0fsV+vEKDo86VRwG2HkkdwC5Er9K0FDdrReedTiOO49/0h4nddAcr1dZH04v
bGI6mO3sFHpDeZyQ5r53ciwR0i6Jbsxjd9F7x5XcNcWFFuIFJM13VZojIgTL+6dVbHsOct3gNu8I
qMyHx75FSYiEB1mPQheyS1cYlNscv4OShYW+EM9V4r/4km7M4Oay5glNlCJ1z3CEPbJF4vQxq4ip
SMHQrgSUHikyGhOHnvhaHf8CDNC3KfiM3Uu1n5mQkIbfW1jWZTTrqXBiYQow+AtWAKo7Fi45lgs4
PUWQwjJS7i5NHQ2tg/EljsgIQcnsNlsy2TOuX7Pdk7xZ4wuQKSmid6rqL1v+Wa0kgd2g/VewlckZ
WtaEYwQG97EAlG0ZovHSSe1NPKOSBqCamWvYlGATyJoysYBbvDFN7INylQ37MLKFPSHznv2Blf1w
DpM99XOliCA1e1Y0YcOAwiLhb7eS3PypbH/wHMzY9H5/TtzQ+iNmz2Z8xhQhZh8CjB9WarPjNe+K
1QQF/D+LiJDwZOnraD0dVtvUY8t+lOsSyIUCX4zBHz550oIrwr1TmnUwiTB8WsvYPNweEhaVUukN
OyTXWpEIT6mZjg5pKfLZt002GhRshytGmqf/7Ld6L87y4allb7FRDQ0164SZvuv36kyBwolYaa5v
7oJPdSSly1K9k3QLCyJzMaX7MpatlcaNiZFsUpIrzy2C6uAE3obP2tWzjNLBe6Az1G2xmb6AM6Y9
q8UbWl83o+rn9hpzKCYhYBIKQS9bO87XIt2bs6JRN3TdAahIA2HruCPCo1XeNcfr5qZlUs0kZ4jz
ojvFpKKASUf3MRTMnom8U57jlEzypuYVH31392ep8bmcbB+FmUZu7OrRqQyeH58CBv0J2JXWpLdy
3YvNJZU8ve5WgrG7uLxVJj3PgnWiRnF7Ye5Fr1tLV5SPJFR8rir4vrzvCnD8G0lfq8hkfEs4oVYo
UQ58Avmr7dkofO7T2bMBYSFdznV80fSTAesZ1PZG+vRHneSzFu5qVGhh9XD0Kn95rhQdswjX5NYg
dJevVkO8ZLkVQUmL8eKd6CeofDBiQngBNHvRCJ60u9USeraUeasYETqUuSv3mEklUsCYwhDNt/r+
Nzy28Gu8pp88r4WAh3HwRzcEoD4N2X5DSd5CMMUKD9xGi7da7WDaIt+QStRNR2wfCnWObjDcw41j
cJD2/BsZJw0SGHTcvtZCnfP2MYnnANIjxOS67Vnkf7raKwI0+x/SukG2s3beYKJL6MEVtDMNKcux
PUAmXv+qjIDh92y0oQZVMLY+D13AjPFr4rEWBSOI98fe8SjxoPJh0laWYxY4yLMcQ+Y4yOIZXybt
bnP6a0x+xMYny1vC2VBKCmRgTMHQEVkv0ANdv1GM4Qjc9EgCRnA8KHoFuctk4C+Vxk56wy3OVC5s
wzInk3m4A+s4JshgNpvIK+oHb07PN9NbVDaNFgAuAXvi9ODrFs8v/lPnInFyYGyPGLL6KvP0+kLR
9dzP1FQjOfGvbRT3uTkCOqMol19TWVnr0BlyPGFrw3ozlq6PcGSD7hMgGNTmLDoHkLG+dYzK0pvV
T1gxO72EmUJprAopHBmT2UcjUEUY9AGZ6KExvN0DJqmygshjPJrdEdFsJk6KrAE+hhvtg8Bfxr9f
/J3cK8Nd6yoarb4uMP27yNb9+U1x/+V24agOtWRZ/2Z9LFe/ZU3CsqHudJDI93PnPfr1RGVF8qOe
qAZn6D6hXnzmDdUHR4tDw+taxvKygWP44QJIRUlUwxbij1i4QTkh8MC1yuj3gNvjuiBWFtmkX+J4
0F8QzgHwawPvCMT1TyOu3c19qdd55r6N7lkxz1R+oBg/wveGqAy17LSkkGkCC7QxX5q0kp5Iejb6
FFpxGZorLBSe27TRbDZX69qP73dchSxE4nAK3mUwqkRqmRWJUueT3MF3RD3TFHSmtJmwPzh5BMFq
t6rzDDcq7eNyzqjs9fvtUPjTEEp0uoHeZJL2lTUvJF3zo9xl6Mhq8Tbeh3iqr+Q50HIUY+u6i6Gq
lDCnwk/CLOm/oJts6eJdWrmSOtRcqG5nu8hQJ/E1zQyhw+lHP5C+L2OE729SeiGjLuVGf2RBoKBq
fjK7dEkEO6TpCCulRjQSVkx5drXLAdRfGhWTIBoNTzJDzbLI71/Qoy9X69aoS/vZcwfAHbtNA+ea
pYGoPrCGx8vQZiQXEaHZNAPt8s1LsPyG4jB5nk8rRQuWbieQJ5hePDveMxDNzj105mqKrGkppyU2
cqoRHDZdfJyxpLAqVu062SlqoA0/WRZuAIhMn87igPSP4cEuErlQnNNU9jtGyqam0pgGsoDXGESU
5BUwppKLaMs3+lYIZ4kL3MYQ7YSWcx6LueRVxK3ip195OwGcSLrHcJHoUzV3lwvPM9jZzJoLkxtF
8ObVOqTWObosnbMTV2E3s/WmOSW7BqtYCSjbgBUCS2r2z9qpQC3Wao0Mdehh4Mk8SIwFn6415WVe
BeXcjfCxAOWg45e7BnhqyNtZKg5ZiLCRYtHXVvRjA60bMPMNDkmgPvbiXYINN8t0Emkw0L2WX0Ba
QM1J+PVqcS3HHJq/g0O8OxlvB8X3Eysrc3hgvXsxbUWpghnDG0q2RzEpGzmWPwf3qBUTcTZyRJqG
y0K8R/fz5wAVfQbv/c+AQjtzlj78zmEwg1tdkts1Qz53ciWNESr+aQh/zyCkYM3bSkq1MUZamTDx
qz4hlnznUSDePQ/+x9HCagHtEz9XE3tjqBpGqRog0+T+7UxJuOGQIJ0UOYmhzREO/BepN4T8gUbQ
56TJ9NdHFUVNeQ9FGlFmvsRnXKnsb8cYe0PMIEC8yH7nISTKhrt+uRhqvYk+N5IBGLEPXc56fUFF
uWo1PewkdWkP9SGimkQZOyHPVce01TPqPVsb1gW5PcuGeEue7SUiX4idPvvQHEwHDosq1qOQ7dcJ
N3sniRiqrJu8sSt+TdAAg53Ko9ly333sSZNuHNoGSxTix6XcLi5EXzXcURP4TIUQ+G8YVtrO3KVN
RTmKpAC8rNDujr3N3S2+6G14QJPCv33tY7zf9fOgEO8SB6F/2XrKlUIxDvmCcfX+lsmdgTSyBj1U
QVnGExkl9xS2xO4JJlRp+PPLlzD9TI52GY4av9wPnOCU4aYZQRAcaTpYn2IIvsKnWN59rvg7WG0B
hQ4kEj/wdDotq2XWz4w3/bJkebumOx+V/+K1OgGAna/e53qzXHQgvQwjfW8/GIsNJxSHcsj3uXkO
rCXKgT698I/RMhthIPXu2TBx8L1ISjNCV6urtOd0lkYIl1pTmF+b3pk96FdfkUCSB8tnxCV5K1yd
9DJw67FJjHqYRWtt+Tt/Om3ptTm8dCyrbOUgh8b4nIZ/zUnyCkmqOQWk149lySjhxQjS0v6yW5E1
OdAt4lIkyMwloZcfkwSWKjgX1OmQhEqKTYQAaXZi+OymxZU0YcD3nchSEdQiO5iUV22O8CNWvgEZ
SA95CZfDMpd+sDZjCVxYQoV4yZbZRfLu7jP33wnGpX+QU9EbYlqD+Zn1kTnplLywyjmUshQjATe0
70iQcEXRLDwJUrsl0VOiwZpQnTt7ZM18IiQXiXd1tsKs/yddM+9Bb4PydzC5CQ83rL3k/aBdL9Iw
UMScYRPdlUxHkOOJvkYIj4L40Tp0INRRuXj8DBnQZ6iTFRUGFUeV6u1R1VbSWhtqX/zIwMFQgoA2
Fm9SEDOgQInvuSmYHTscKlVWmthU9UXTa22VbD0jseJ1RKAjhD1KgJrDdmIsiTHcqDnMJqFud1n/
LDDK/Rfn9J9G7Pjj9S8OmgW0LoLqxQMRER/nyOcCy7NzkM40sshFnZg6G/aYz2hdhxjqrAMxMgNF
tPNLoaiLfvtDlIQXopyR9mOnMRUmxWV7t3hkhAcAhtKCgXp4L9N/GjLnPxPiHrE8J8rRQ/170NSi
aBRFVoOvwBIfUW4rdQ7z3geSp03HS2LNBhh8AT5CQgvzTdohkGJegGlnmWzF96SDI/1otJQAuy4l
yX7oDUU/3D+B/1nTBVdPc8uaJ8ZQ2x8KbVhjw0hp5Sbd2NC4RUF/pSnzH0II0IN0SE0b061xXe/1
87DGN2/sKYTnhscbtFlh0KZdD0q3jStQRz/zPm5J017ToAzHLSjSYNE9BCxyy4z8nJxU9ElgOIcL
1isDMwSgX4zYRTOZBwRHYuM+owwIQPr2vL0Ae/RuIhTC6rvLyyPeFpJLO1wikFvHBFcA2AgVxqb6
vT7Jt3cM9LMXJYd7z/9PAPGAs8Po3gqGcg+l8NSBshbuqmz9pcxTObkRNUW+fYml/sNB6s1C1x4n
akGCbEaVhJf1JkBG1MAUrPAp7nvtiqTaCNKeUzLN7NsWDHyG/s+yN2+EekLaeSCrh4ZxuYyDzbcW
LCCpbGEqZXitKLgALKOJUngHWu337Ql6FSGfQ3R4u068NFwvbxFQnqrws5s2kAMU24Q67HD60sMu
WqmPWHuUuwElLsAX+jGEW3/OCcDq9BWzXlUWtjKs47yPy10P2yG1vVs/C3psLcLsEwi3Wf3ZehAO
rN80CGxl8RQeHbM0xHmmOUUVdNxxBcXoS44+7V8gm3lhymYvT2mXvzERfMigcXvncnFRSyyOpCba
dfGQKCRoP3d7HmhM5m7kG1Tdlk/RGQPDYbKSC2SSn+2LE9yQi4HNLn5JMg9l3RHBzYyKIKbqBEok
XokRVwnwc2z74oEQE3GXs+2AGvfPFc1JggbiexkwxsKhcRVIGMLa+SNacwcPmjwocxReMPAY82KD
PqOXSNFzQgv6U490pucXxlBaHZlXkB+BzGfL9+1h6jQ10QWolQITCvUEWDKDv3127b76ktkoIGnX
q1mRepc27FB1Xca5I2Jdr/0JvjNDdMsYFSItqM1gRBMZnxBtrDZBwNOePcdlhIpGR66v076YT+V+
WAu1dQ5JwvNk1PkvLIMxxjqmCF+NkZYPmXX2JvGgKWlXDunwJ+pzNfG4+Rgabt9cegPfGf2KWDYn
k0gGBaIDgHhkVTIsbHoXmB1zIphNQ28Hsbs8qe1V4Q/zmB4hLyrBUqXOpaBTv0dDd2jjkydM4IFT
sKqWJYSU4nnEHZXfvm7CMZhDCUtS/VRJmv5anE+XsexooFHUlwFyMzbsOr2MZg3ew8zPdgt3Q2MS
fDeZRKGEXiw76um7sPXrfr6pcEKMmUmTYYn4R3S5R7qfmnQI3hynX2x6xU6pX/WouwxwcHxIH7PG
dKwjySCdQCgYJZUWL1dQ0wGpMWJBS80xS3oYsvaSaUpQiD/DZND2qaz8RuXRNAkKreEXZlUTrbp2
TXrO0GkRXjaD+su5rwWI4iCXi0NW+Tlhj69C4cCASe8AgNiIr+XNE5z+sJBFdgjRblCkoeLxgjrj
2lzQW74RXm+WzVYsaOL4a0GW28pyjnSdEJjijCCqRQHUxdCzZrA+Zm7Lr9H0OpjECGP5Ia4+FbDr
40f/f72hvT1f7Ut8repm2VjipPlCkOfsEh1LacWwq5e6Kmc9MxVvD7Ae3zMbOhFyF0nEvVys1UD9
kU/TuqVp6mBg8dhOBZt//q9D5h1sjKlG5+Mu0OP6uSBv6L66yzQbNmVIh8Q5sKnPvCxR/ToSUWnd
6vgwe3ZVeA8cAjHfNLsrYaln7TLhXrZEBSPV6BI6wgrFbndyEPt0bRHvxLPxysEuStH4nFmIQV43
SWES++Y6Dleuovk2pDJoKpxnuGK3yr7N2ZR3yY9zvc1z9hhOsHYnqNGm1L6Fdf9Z92QK0cDu/uhK
TASw7QqgPJyIp2zpSQSqgfE1XAaqkp3sppmDVtDuWbSFmHQOhMh8b8oGEKokq1t48LhvhUy0BdPW
L7laBiNKaZWNqVbgK/RXTbUGro/zTqMsz7tlpjrQcKgN9jWtpJc5QCVOfkbilTFjeY6P/PEhqjva
3mrOlx39VUwfsUi56Jk5py0Fbj+MRlmYqoc18ohUOxBJ0capkBYSsY4JkQ1eM0xotGxezs1bebTM
uOkOqo/wUSk16+fPnzVU0TObpZkV2zfTleF/sNMYz+IIVidlWtAYlbL4LaLhz6C3eStu1gyEs+WL
aLN2uilGSZPCggogkAXoz+mopOe0DQpRBXHDiRttyBxqAyHCeDdpcT+qS8//TrQh436JXZ9RSOKW
eLAmX61kgLOHiJ54GbQ1q+BE8FXRPRYHgeFLig38BK640/oDm5xpsbBbBokDYY/ai+il2KjltILO
QejsJ7zjw37aDJ/xH+BSoWx18hhuYBrb3uW3IN6QCM2e5DaqaHQB90sF2RaS2u1GdLq+epeZTPbm
4r6IBXvn17kD531k2uMrxCxwnGDaWNrPR4l0NvcexUdYZwjTqwHrzqNSfPfBgEqqOdO77WG21pMA
kccdA8EEegjQhS1uvvt+/pGtUKW7xtW09aN9h++AVHePWsIZd2SoscmHNEvLG3Cs1xhTDr9RCkWq
1FbLPlJIUfxCxaQKruhYl13dVv2zcB1Gjv1IjpMpWiilkTEFBrOdo1TE6gqZY8hhXsfhV1jrQqjU
zN4tmEQL9EuFClGgyWN47/NLKV5DQR1AAaBVGSxCXBFJjfYinnx8qn+vI6JaIIj6JZHdcqyROVHf
bfveNzLJ7fkh+5sNVYymUN//uj5z2YHXnF0VPjuiygeGx93UehFpKOfY7qoI5/O+EdufKXn3RaKy
axJ/LPdboUHgDnJsrKSYQzLl/u6xaKL9cX9HjN9Lv6kIq0CnsLsv7Kx4Lk3rfLfag3RKiEfD/CSS
AMLv2vkVFSgM1cfamAtOSYDlRmwjTr1+r9nIgHlvvwinbIAlU30H9eiDamx3azt2pesyTcA7ECBF
FyfMxzm5U96UhuN1aHmvuQOOCA8LhmiXB7lvfIAfdM1L+Qod2YvSkVLp3AyLwe3BYouK0WWKcKLm
n8pLIuJ+v9ewT4rb5W6s5CtxZ9v8n4bhOOTfxOOtB+FuU+LLeX/C12jt1RvICP0nLulNZGV0p6ah
UbRLK2vH6ZJG1oxHjNuMyrGysUX9MY7WOODeoPdBlN0NY9M38EXDcjXXjGHJDeA0GV53SNZdEGTD
CXm+FUA52n6IvZjSUCoc8UN8/tFeqATv3+QI4bzJQXMyhsCKKmXwIU92WULkYlR+Jx/f82ujsaDR
OxQpv0WSiB7A1VGJkCjtPCYt+eaOvTdJZc7/wDpmgleIEUCfSIIVrEkinGMA0z7jKYCdY2UiXf85
ALirwOCl2mLMkjSsk4WNx2rN/eJWt0pFcmX2iKuM7YhkGfeenX7xWph2vHI6T/Mh45DPcp5rdDcU
NzWnBVpo0PwmL/vtGWN1WWSxnGBYxIJ4D4DePIfmtmXTjAsTT66XvGazIC9dJq3Fdugpq8aT36zZ
BlY35wVaWn8rfEjMTKYe+8gXbphJzMH8TXHLA+J7emWN82NzwLJxmcxVPcJT/RybmjIXKHJtUOwI
vcI/NiTrVXLKkeeoQKBP7EcAH5pUQq+HbDBwRssqodyzHQXeZWmpcij1sh20BOoJ7cBrUDaH2aUX
WQo0Tg+9tNkPHqNU1htGt6Nx8Z6X9Ppy7MqCmRlmv2iNuO8IL3eBLgnw62Rg28jJ+FAPUy/LWGps
uBSA503NgSNny4+LA9NyeD8ekvvALP+ijysfiPpMi86SuMhbgNFtnaqg5AsecBv+irjQeB+VkunR
//vKSZpRA/rx1+iEDPg4dOtNpnZcPeiE1ilxRO5ApUdZ4qkZl1a/vX7VhjSiLL2ez5IfF/G2Hgs6
lDO+ro4hMyLBJcxruGR3Nq8szly0N0VExwhXU4fNnvzV1cYCDGdO2a6UbgCEijJhzCruYBdsibuo
sTxcfFCMiSfukiRAPKdJHUMwtn1zQT8NKLrB0Vfnx+4mzATfs9hVOk2t1J8URAGreB9sPv59dQoa
NOKM0bgOg9HuNMhA6jOdm1y8ArEs01jLsS7DrCATLZdWLQ4huXMdlQ3799oSdJs0+IoW08iEtocV
r706th/B4BvpA/ZQAaYDCi4d1mf9eO6Kxhie5kiO9E8UCpTCsIwTdpjNNp6Y7iktgQC1t7+dilqh
LPtjE77BZJgUDjHj61fmi77KhdyoDk7Dj7jpfPQOpLlaxGltjevubwhsgaurH6ZDlpu9KKLNKsGO
XJbsPcZQ1Dv3KzMn7fWBSEmXCzC+MKk6ufIbrsFbKs32ALt9fwBxgcOhEntsz9GVohKemqJFNXcq
JfPegsc+9VethdWbXdFCxlIjQ5cZu/aYVJ8au4LdkCZUbtBbRnAfE0IRA1IDp5SBpTKML6DEb8Ld
7u0MGOZo0lMA50/PXEWmarKhs75WSlI/OmaXj+oE848R+x5raJl2Z9yu9Q8qRjyyTv86PhwgU6sc
jNrBbJvh4Xsl9YRCkJBJAe6ucZZBXLh6tZWU5xOdV5hBJLdlzGVnK1rD0D8sMawRptlgbByF8I1l
VFm3TWSS69H2nBHX5U1R7dfDkpMK4oKLkUr8wXCmEh3JzbeutqWvHh3LQc3HJebrOu6ie2nz7OW3
kVJ5xlgmmylelRQRwvwRUGWEbuWzfTgEDeSRHSMb/v+P3hKfiDNAWTTl8R3a/8B8ML21mHCWOwh3
WO0zWpho/YIAZwe315VZiHK4ly4WLmf/VaTfh4R1nST/WUtGLYPuMqkNiItquw/TwAEpYzNvS+Mf
N3hBHCf6mPgWlw1MqlTE+yJ+Y0nblw5WokJu/+fwxiKMvprthy4Lak5brHkWsx6k9UcTlYcg7tyw
Ovt3Dcfl0Wu29jC781eQA0QK9X+1EUHUqyY5TDiZo9VQTIcYgHz79syt9Lbus3UXVFO11K4aUMfa
tJZ7+3/sEZGJsO4jxoAWFw6m5lEVbQvkxiwU/teCI1GkrQp4oqdG6shKNZcl+iwDZxAyrRyAutes
/DIGfABVTcQfnUkaUXpHJoBLvUcxTFiym06bUaRJ3JZi7eCZPsWw6zqdk044Z+q3cyD1TjHJfhMg
3/1ExTYdKq0oC5FXTmZ8zhQHBQsYnCxy588Ga0ZgAoT0gPheoZCetSLDU2TAP4KZbluS0Ou8Z3oi
Si6mEGD7vTcQ4HmbOUnvMs8IcP7/om6DWdr14vHINhT5tfgNxBQN32wTD94g3HieHK3LQ2Rky3LL
m/e37/bAOlzRdBxvWZpybJyUkW4ifaBD5Ao+6lM1Qz3lvrw4ZD/8oZQl0lMoy+jcFC7V3AT9j0Wx
JZ0H19xBRiZLSAIR+WQLNCLWc9fCnuwRnVH1747iAnKIzETvExwfmN92OzNbzKm10uUNsHijgfjH
3Hzk3R3Acvf42ZGOCOM+XC/KYgXrJVbV70HJ9qD+wn58OruJREKkLfHVb5rJyxu2ogc84+ggR7K4
ON3plNCBtLTiKZ0VDLiTTF6rIGDRiymySHnC/Hj0psYt2KiZQR0EyHbdCVKAW6/zwqCu4eio4LAu
MJ3IX2wjKQHKiOPdjNQr3IkAMbE/dOcMZNBXUISAJeApXUuVREWshB2VMgdUQ9hZgWhpHvlZ6OSZ
siZNOWTjTZ615V+7zqMZ+89gmD7QDGj5HAB9Fr9yXqyEhqmWiaLwqi/E2y7LfN99DMkZExg8bA28
SQiKcbsOqoeJMtUDuKcjF4nB7rh6ls6cNGw48av3sMaLoFc+ipIin+1FdWQYfEENyhEW7m7iV5Cp
1xbbQdAFr5YrIOKqNDgI33iH0ex3rbiP+i9zwjjJR1gbGahTaef4YPS0MNUxDGAeBylLeyRv0NVo
3L+MDqvu4NJaAYbBNFwEPiOBRTNWsy9MYCw6RfmZxz3/mUNWrUl1Fl1OnUXJdhZcTxQgvBKGxW+s
ojtig21dJZFVRVrLRBCwvfhIUUnf/LNCDHAnvvQYC1d3eu99vw0gjtMGWcWWCchVb9lL4NTcB0ft
SFc15QdlEJlvbwniZ2cEjcefldK3Rn60T9EHuZqrn50daa/cgiYxGrjmcfeCFpyREwy7DpNXSesk
V9Lyf5YpXuazWDAZeJ1DbJxH6jVzBUHkVDbJM+4qkW0GuLfQm8tlxD4AEZAC7yHifMxGu2wBThqJ
WEgS5wojzh9Aki4iErfc1hFkl9vSyCkZa3J9OVMZU8aNzho7sye20hwyt0Ywh3xcITZFk5Z7Xcn4
xBDx7GD8y50UvyIOm7gFfr/6+h3QDhDD/+aGwSIgMdejXOFVnpOs3uiSLF4SkjtxmqwtZJlef0zF
AmvWZIHuS1YiiZxLYvco11epM0jtpTH9H5Z9LvDy6M4aA12g5F1LfD2AR5wJ0dfQdz3ob6ny3Qwh
iY/M5zELR50/B8SyGW0Gxt0DbhfduBRNS7do5GsjBgPo8HV7jwsUKwrYv6EFpFb0Ld/Vj8Hl/ZNH
PExJm6o/TFSaQhuMUe4MqFTusFhxEI0uq2bfRfX/Ip471Ma1y9TMDBpsc91VbU3Hv26MFFncqw6F
lRCcUnVP6QsPuWgVRfMLwPAzA8U9pZ69U/kdLSOCE0e9hVf1D+1DAQT1rjALADWbNCp9rruAMtPB
Vtm+6RG0JNI8GYwZeR0TFB2XGgxbWATohlldNIgR26zdj/2A5+qhAbcQqJyjdR1NZsvwl2aVm8/T
uEnsXnvqX6T4c0aID8wyvNJ07d+I4JTzhgkWi2qOi576VYOgDKD3oE9xXwFiEBGnmuVD7bbBu3Ht
BkrZbwDak6veOlpIe02bo0BmJewD8Q65JVSQOWMRTyJ57XpSKksbMkGan2rGg5q+jU+sjsRFhy7t
HJ4uz3FBFQQltVA7z5QqtkL/PW1cHbgSMtlIAd+eHfC6kZF0aYs5MU/G++7Ul8A4lfuuBZ5K1IXv
JiMhInQVYm8TVtOVM6g4janGqLqvTfZDqgxZJrtikaF8eptD8P+wrpXCSCVtS4zIe5VpgHQYP85V
srFdNmgbXLPbnULAlAcZZ6PmbyWsTXoL3IE1plcbC29H2ULKAtgSiqYJMZ/nLAkO2ft6ceAQxjSk
rsta51EacI/UE2ctjwhLI76lzbs+mO3VOL7YD28Uhjf3mtPNaSk3YphtkQSImbOgqEyhVwLmENmA
dnmVFafUt5pOky2/kkTA9JJ7efjp+qqXI1oOGT0zVotOYmJYguh74kD5LJUW8YrzcEPr+R0b54ZY
CF4yvDcwW6k8B0LGy47jvMBjIwjDXpLzJ0rk+paHXN+CJaU9PBJaHqVLDLUJ1WAmRjyYr4cYMgVf
0JwTova0DH4oQNB3RZfaJXRfE68+gS48G/lJEGtSRuQhKZWiJK92HuNz9OMZREJL+Yw2VtkELObd
RZmpeN7csF9aPudQd81Z5JxuP4+41B63FG3LW75h9AJc3UF3Ctn9OG/QrqPCZDzAh4dogGpNpiww
as4/VOunMAs3yL2R08bD0PUhE8KRFQQo+WhpQV5AtUE2s2YfJ30FVqw7ii4TYh2TjXMumsjqmL2K
yFUUfLTiVzMcd90UnyNpSWyB5zr+aKAV5AQrqncr6Or7Oz6Afc//+VKuqADfxJafMnRbqeCg4dCb
C9OyLRaCFXht8JD5qeo2hbLSlMun9GCyiAhyW3aBhUH1RBNO6iCKCEtTRXsAy++46b59orkaJ8ux
UuP4heIG27SCMJu8AfolmgkXMqQDiODHPRHQFWd5r+u6pL2SU1CHK1D+XcfVLia5IgIDzwS/yva/
1Ua7PfLKcfQzy+BhQ8OOZarwY6/2DwMlKHNuim7H1o3By8Ni2oVVhD2pYs+OHHKE9Vi+i9Zpu1kQ
ZXzVH5T6Af+9WS3pNXVT22IWxnVPdkGcYCVgOUqxmfP9hOg6nmG+W4KKXE1WkjvLRRZhHLobdd9w
JBOkgiIsxveTLtEliEdlK7nqmAU1iJghNqr7F/qrWyVI0rG5d+pxAKKNrtPsQQRn8ASBvri5TDiU
kbpco3H/tisnLoMusM/nBkKOjholvU5CXH6dYTgQ6TQ3PSV1lMPNP6zNsWljjxgIew59ONe2G/1b
lWWgeeqPua0lqX6cnBRM6RCfbtEqA7OimXZcjSSXWWKiHoVGeFD3oDyCJISvVLcYiugRh1WtJQrd
mjLEiAkLtFxXunPm8MTSq4aQEExFJFBXhoMc99rFzrSOKjahtKoo6SMD28eABYHq3XZ23LSJ1BTB
kd5zaPPxnuBqBZJjPUMQd2ecNGQxPimRHcjrIjBuqvsA5ZeULFHI9dKUyLCvhPVcsILJNmC45dwR
GbsLaewP9dsUYibsMRkiT3iUH7V3cfW1U/a4xSe94NUQkoOgsyuZCpdyXhlGdBrZBaQHMS3uZRj/
Shs4WrLUaU+9FvMPlvg2A5B8qy3mUhmNGYCTSslpJt1IToS8L1MJ8GhygqWder0Vzi/Hm6FYQjZl
S7u0nJYsvo60na0s/soe/yGiRY6+71JOPFzB4FTOiKKCUYpd/6lRAqJzyLdvwrWKgeHWe/qaD3Er
mVITvSc6lDOx/1XUonq4PSewpE7aSD8RF8YcQF2sT80MIcas2R1CzXbeWXASEYO8vJUgYkwBKqFs
QRRPk43rMUQxFKzM4U7scFA4NzaJ9Y4FqfYZ/hXOaSbKjYGvqV6i2/NAeEE3YfcInIl1kVsFWHaJ
IT1QMCvIPiZw2wLDbn2g21WO5TQEz+Xi/ch/q5Sw129IXucigvDOFcLYSBO6glLDzvfa2Xv0B2Zo
4hpKCQr6VWq2HWdkDZrmEHwZGbuo5p/HGReL/KZDXkeFdxTqOQU4tbR1Ple6AK7IfaIeh+gN1dzV
9A345vbYQVYXMsbZgj1/xkQXq1aQaFUMMdvdN60nODQ9iSgKIEw18JImIqGJq1i1x3W6gX6MbQOr
2B/dNCIcMhbKFRY0mQ7N4U4lSz7xOEOhtWaFHplYMrNrbbJdAsjLil1ar1IXuPJXwDleyCOKr7Nh
ljmDq1XG1Ggpxe5YSHilYEdvenqSekcNSaHq9Rt5S+Mo50oed8z0xPr4kx1IChN47KtYf96Kf7y6
1RcDCTTWV+mQ1ywAHNWvTkvu1uj7wko4gQ/CLstS+rnq2VTopomWdQq8eT/AqUwbnLD7K2P+LZCL
CKbJA7H/6RheGmkT2R4ULHmzdFgpdWbFzVasvF+lXQDjsKxZtCJTSZM70WtACpUftfwJkpIXLhAF
uZM8zj1ICTcwZSpJTYOxGoTduNw89AXSyCmjS2kxZacPReJMBGhb8YTYJJB1VOoySkT5fDdSS6tZ
fABBs1yEqNwomi9N/hp3VPRw+OCaTdKTSQLS/G8twdL6G6+hZup6P3cdWqL2JngDZ0pVrUWrikvo
r5A3RcgNS/bXKLVImYJ55xBErZEzoDJ4uuiNVUf/ily/0k6ifsiFvtk1B/tMDtTuXc8YbqddjLvT
30HuTOYDO8aQkk9pWS6G8wCV6DVmSy+nZUMGGxBK89rYcccAmZYFjy/70ErFQEok5k/IdrlEuqfs
MDk8b8ZeFOIDRWQQmFxZ1LrDISMTbLeEfYIrbigQlv0OBsPBANvCSKNWNfG5oZUSDIGDRk5Da6fD
0LNLrfhojMUCnNtdAKaP+Wono8DO8XyjYHNJEn/GI4iFceNMV6DTyIltz96ZIYZL9dP2FLtweASu
RJkPC4Kq8CPy2+ChbpugExCsx+z+I4g9CcjXTPfydVzBmuv7BaCQKDqOF1yqE5Aifni80h/fwO7a
dN/XzsyIRvdBPQZKqeTkkH6ZzyDPva3f3Q==
`protect end_protected

