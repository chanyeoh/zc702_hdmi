

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
pDML3u9epGA/dqPpaSpuXK8NEksQzonUB7GrjhyBg4xmtx9rU8AqFgwUVIKfxFi1GDCYlQlR5hVx
tnCjksgEFQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
TrzIXaRW+CzIv5Z1S9GKmVl9JTQxA6Q1ZG4bsbXj/luKGQwm5qP8/reSml8WY2QMex3BfTPfrs3M
Lmtt5k61cKRFBNue5drCj5os207ZLmBV/emiQkmxyZL6dPfkfosBiZgwBhLbel7g85OqUIltLx7S
9g3E0W8CnkdPrjmn4hY=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
F1wAvGsi4SB4+Fu4huEGk3cttwWefJ5I7NrJ54VTmGzqUJmfer1+M1LiLhmG0YphHkOGfM4ufcKW
DsN4quSRsB9euev7k5+BGZACLIlh8442XFduQGzyYsOtkV5+PsWIC19Va1rY2sI1z6yTkXSlkyU8
XDSCK0zE4PiSbqcVrbsy1Y02vm7LhBYu0kUB41CxT+9dmDtJMWWjLFG1G+Tn2o3tMyM1/S6vlTUJ
jipPz3Do4SjEQI+de5vadpCtA1vjukX1BbOFO6aorysUKesb9dO/dqFRCSuHKi6jHz9uUVZrHGiD
dNfoWpKFNIJIO0HeilrkTfgq7AznL63NZr9E/w==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
MK5ljV3f6OvXg8e2VwSRDjtUNgYg1coasIiLehawmdBQmNdV9OfOGe3ZHpNEEzZlV4yvOHex2ViC
CdqxTYQD3vegXeKNlAFt8sgfCHvtkNmwDTC9/VY81eUqCchRWRXkvBlAn8dpjCKgoNU9bv9TTjot
9RdFQjsBlIEO7O6GLGc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cQY7BoloX/rHKxQVfKkwwmPMmtazTzye7h85GwheEj6g/0nYS7ReBC+s1tkNO9gKdW3T3DF132Tu
+fie+VgvD9hoEiDY7iJu6UsIEdjucxbtQHNtwjWGRf2MlixAm2l58TnamnQp43FmGpUcU7Kg2mNr
Oz0ErOtSs9nP/iz7o3fvm096Ly463VHd8WgMmqI01f0Z/pi4PoFQYqOVWGh1dgvNw2uw7hNLLr6U
vs2B3FhbArV1BNDX7PGWf4ywwvY14zMXayHOKDCpGKFlyzUVLhpSoUUwqBx0mTi3YgxoxPjGbjb8
HXenOSsnYGmPG6cOgLhySVTpI4k8UFFyKEMQNQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DeFo3CU0hqnJ1Y4qB5H4WHAMnGy8I2i8IymhSb8fUXDJaPv1UvY1JeTCN73rvfQiORkflu/wK2Zw
fLw/UT434z61pFwB6On5UYe91/6nPtZFYvmG1KRcn6rnUr73WPnEWi0OXGX8b49PAvZD0URcLTBZ
5yX3m3j5+zAmNP2DNaKE9Ayy81ZpCVUBqkKfTrsH7mQZzNaCbv5hwGpkwIQwwtUvskeAqY7oMXf8
ex5QARDpgkho59a4X1C6XMpliXk58TmAiTiWM4MMnODxz1++RNcstfGajn6bfFLC6FUhJjF3iYmt
5C0RkeIt+hQ14lGVEiPvgOLOf8YSLflx6LpoNg==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 833648)
`protect data_block
gGpefSk0xpZQ4oLZkpuJzlRR/WL94fOjD5FwkTNQsTNH+TBhJ+msdlX7SB/P5tMVY4SEe7+rihwN
JxYBR19L6x6ZaGoIUf0Z2I0cekuHsdgV8bg0JUfUqBnIedEKYFqSN19i5gAt3Zqb9Ta56XV48upR
cDvmDFY1HmgmdjsNUwptqJIrgvfO6GCK9bnJ9a9nPQfUdDNHhbzczAPc+VCG5redM8b6YGSmghwK
jmwdMTOUjBOyuxKR2ml0sRLnTa3/YqazC6tVQQCoOgnBKxe6u8Gq1ygozpnbVGra/6y+PYIwDv+f
sS23y6rl4SwpGZrozBWWe+YVbd3+4eJeaO65GnmOjqZqNEwZrcArINkCoQwOIGF0bZxfwvE+XbSL
dsd5NJQntWuB6V3B92I4UQ/0a15GT96bmXkrwy3qV8J7jiutnAkWh9bxt24EqYlZrMFD/YiewFKy
mgPwJhFvCbEvL9Rb6xXsl0Q/G8/s2Pj51aMCzN80ifi8Q4gewmxn/vX1ThiDj/PBP1XstspG5C6O
+V1D+zGzHUPHH0gXTHun7fpR6DETatw3EmB2jZJjFCTVvmfGnhJP6pcyj/piitro3W9syZeSmRBq
JkJgaoRpnqKBJJBXrfR8zAhO6emrYBkTz+oan/SOwEmkIslvpl+LaHRVFVtRekIseiwGCBR0Z8lD
IT7yd5Dl+bCp0w7Z47QxwYD6FY/Oc78cuNp4NoxOk/6l176+6339eJtwidNFuLatSaJE03Re6GO8
UNR/sxILsmM9OsWINuSRkABY05rDTmB1RijadEgzemnooecJkb7jP3O7uNiOVWfdHEqX4ipIQ17l
jcgIUaG8/OcyXc+4RqR1Rb5IbgWFBv9BbXvkLLJNCO4VDvxeaU9WjcOrJoH+4dL0b4n/UaXx+JFZ
6iZUFf8KJR43aIkWw7ar47ioEN1lZlOKkGKsv8NnmcV5URhmuYvlNHgyiNogwpNV1wr4gtv/YIG6
FdXXIHvqPXf+dZ5SFUjs2HwWDjvAS/de5hyWDVxPpDkwBHwGZPWN2e4irj0lU6Nuogp4hA6Gj4DH
F4SDeKphmUnTW/HqaizBJPizAwZyGymkKVWwQbwsfzOTv2Qdh+KJbhNZcM1SrxQxRf+UglmKBk5o
17Zn9JWZCT5KOJIfjQ9j7E9DFtOpseVwkYK2zH7jiyRyeD+O62X6Fv3/6AzEx2pzBIOGYUKa1DTE
0uPGaYofC7SwFZmcJNRT7o7z1nyrVvRgkCvIupuEkl8NyGniJArIurq/HCDsQyh3PH9UlNScbDaZ
sIUnsTSzGGU9NnmWtCqYfbW+1Auzgs62Xby/ukhVw6/iQptLxXRuqmkoN8XnIjZ4EZALhMCaat0j
aBst3D2O/piL4qS49w40IusgvQqrLRRcUI1Z/Fo3OvaEJxlziuhA8D1k9YWlzYzGC1CZAB73ZiWe
YlmWosozv36yP+UnhA/x3wHPu+Ne9111ZZW8EVO44DRdAyrSNr6VcGDg4iobpIsBqFzsPrsxIuxY
iNaAykFWfy8Tnls6xqjzxcXH9dLlTC0ZvnnS6OajE3MhiJAsEirypgwwp/WrviD/V6fDsVwAExBg
DpmLLou4PHeOHXxaCWvHiREgAj985HaOaN9lgFQRc42rP9V574P4UjHI8pnTPbt9vAO0D+ddg3tn
/DMKLU5DUFNwOnHMUM4UeJPQYQwe5Cz+t6AOVmH709x2Qv2bDuEbU5p2Ik4/JuKdCzVXXrxgVaye
yOUsEDrDaCWZDcQOATIBKI7jK7oHZimqw3P4ae9EQ6NiCvXtx28g0B611KGSVriLLNHpOc4pnxop
goKucbXIPYRRbOdzCtGAsTHS5kLLXELD6rCHNaiwwthRulQfH8yqBa2CN/++hPC4RJrpOVSJTMWG
7t0vNjPDfWojjWzlsUn/Dv1z1gKm48PDz86Wgr3cpNBJrCcNGFg/ugpCDWsPHiHdqXbMFtbUARNK
oFDgjKihT6yFpQx6CmaRpDKXNPuSzBuBXp3vUZR21v20qOwdS7yPR8DoYBGpgEQFsv9LS0/JuuW3
TtZiB+gPXv6LwqjS7ScmXXP859yiAOFCTYw20wgSuEmXVl0QfaeGCIzctLUaJSIEx7g0Dj4Fq+C4
iJAX9X++6D73F+BSyBWyhb5FtZ5JHLSGY+fmp0d3S+eOjfbKoi84pLhBT/iU60gI5N2B1iFdJUMc
VodSBZGclj/WWWrHLudd1TJeYSKhziu2PD0tP72vD70RmE3pfj0ejFumx8e+OxiAK7ZtRM0bTtaG
/wDyPdcVu+hS77nw9nLLkG1JsM/3wwQccP9PMExZkQ80h3rugZQ37snFvPrJveNyuKvPoe7cyJAh
SEEXRKjFFegekLjv/dILVwzzSt9C/b8nreOyjs1rX5yUVxH1wsH7siRLDUeuM5U8Fwe4ScOd2uwl
twCZd3u/QnDRC+8OAh+VYgCn+DuLeJhDYNvW3t5o6c6dcNBL4tkMVLtLoD3BJhecQkBgu4bAAbuK
vp++EZA0JvH1TEL88dj9XWxq/C3qhw+5idWCfsamRSlooAzE9XtsLJRIorUnmikFgHH6wKMI4sZi
Zwmf7u4F9u7gKd9cAJgIrs9mf5xXewUVD+D64CI6i9boFmqzfSwl8pCwrlkC4hcuBY/gg7JbfCwL
3NLqSX485IJXfbrTWb+xRh1E9i9tDBTHsuO1/nmIVzONz42vQ250QDz+fUUdXqavbcQjBfro0X0s
ai1BCgujVUInvnH5Qkl98qSz41YY27KbsNBv6tp0MJ5rGtRKubLn8vjiQL5rM3RC26WK6IgxD1uP
axr/WcXCoLNatf6ceP2oNe8DTz/pgp/THJqR3IWW2+HVLTR1o0U5twwpydMko8hpG9csMqa7dKc3
pagngFrSHXsx4UARkNL0w8FtaFMiHvPS/CVlmNfSVRARnCWptxSYw32MI3OQ3nt304LwwJjDP2Fz
fDJ/OfbMOhWAg+rXSkgqUqy+OFXVI2X/ikI3xK0D/XLmcEQ3w6l75xCWilkRm41mP8HY1zCmD2TS
xkvbPQ1x1xuQYleOZMOuXaqJUuV8F4EMWuqce6vrPQyO+o+QyoIc/JPRHWTmrLsia8iD4Vd2CyvZ
t8TjDsMx+1NB+dHoQfjLphkbUXm6/3yfrW6su6vpQEAjct/fFXui0FbSLSXIllfbRFr7jBvjAxA7
5fVxMavjZUB3UzOszhTYR5KwVEiO+suHecuOmlL/6CgwnoNKg696ohuVIqtzgtZNQ9yrBZhDTzXi
YlKBETBPHaoLBw3yWX8nBiT/ff/WK5HrDlQOpouh43mnJacdefxm2t6si6RbcxPFqGKww5O2bWQU
cedUVHYSh9ZAxhv43QwA/RwYgVVVXmerIyug527tlTLNTLAxeoQP4up0piFfOPReJkms1T563p6A
ZeEX6qsC4F/fhMss75jtxk6LF2LPT2Uejkh3qJaZ643HwuubDWCxDKyaLGGJJbvEZOtjVGD9Nln7
buztq4p1O4xgkkgSJnMVRLyh3vE9NmIHridEbfoezcCgfHP/+GstC/WnVm/Aldvsii+P+Qcz357l
7YUt4Pt5KWPmztuS9ei65HroIsspCZZNzb1gcPoOS1R75wclKQ0n+oPLg5XBfDfcg7HNWVtNHwwy
185Fr0iTjbsSTNbzY6LN7eLxbWBRtlsOe6Ou/+MG4DAxKFQFBVr9eYw2N2evCBihM4pCPrA0l/DZ
bEpOv3C7OxrNRGy7mU+/csC4X89eVG08wY7CInGuM4dGHkpFrDcKCU4y0Wi/VgTJxslbFpkAqMLe
5iqwGsYgfHPMN+sTy8gkg31zOLiTAMFWRceffyriWOXrZSQdyXDkYrW/XmIxJ+dmFQA3teIDByRk
XZasUkpLkXrabSQhwQs5rYUVndMw/K3Auc+pNCet4Ec8jmXLf1SQyT4njmvgFszf6e13FhDo77GM
AZnargn/dx7bxxmzrtVVPW8v5uzGRqUmIeA5PKaZjGYvS3eRpA1PbWO3Gkg4iY6Rs4W15eNQ04f/
gGu1pmiId6BYXC9cJ8HIREq+5qmJdngD4UWVFX4HApJ7D9BceipI+Cxv+GeLr1Hk+/9wjNKhG4NZ
BJeoL4Lwa7SCHqgwQtLKO0zHN1eAEqPNYy6EUuG+O50/oSDa9NK99E/pUXDquLuM/dXVUqzL4uDe
54OgapvyEBh5+K3D/cLM1tyOGZkhDXcrxnOJQYe9v4fpz/HdypMJqJMuhVQWsSv7lVmKJWpcJyLF
dB7UjpARKog0HchqdQWmh1ClL/dvWpL8+LGLacJnYJoNtu+LgsrUQn6sY0bf3NnFBqzXnqvn4od2
vEiRN2CDqGump7Rg7oxu7dt7MNmMVCUEC2GzVQeTTw5u5xF+B6IcWyd6Wkt95cGAXEov7Cg+3QH5
SyMBiiKe8wN5g7DuxvLPvYrGn/S8T9xfXVcT8WdElOPRDL5sHZy+v7R8wF7H9a95wfI2BTLMF9dz
aGrvwJdUGXYcUFZN/+4S25xdoNsL89OeRbONSdfD/55SKDngptBxOktbaUQaL5iTffjGaDZ83oVO
fDcXQ7roVbc4Pw2OwJsEmWLsxbj6c3WZ5v9l7n7E3yH8LsS4tVjKmqKPWu2mJLgsT3Cqvho2foEh
D47tKu2sx46G/e/ApCN0mkV9BHe4IgjKTm/zzGcYRvTqcHihfCw/dKEqnQbe+096uLRr8aq3dw6v
+9b4mrq2oZdDQBvAyNlQNX32yqvyhjeghyLGOMK8Q+MH/iRaLyU3/qrqFUmv52XaWCDmuuLr/r2i
vbc4cF+BWmpLjco1/58UsXu2g9Pc+XI4vILO3HNUYf75MDqxiGLsdrNcdMOvpQpcW5C+BxzTh/tZ
BNzL7TbrS1B6Kac6+G0HWYUdID19+OpHpIILo/4TEmMtIUO18x7q8KikHw5cy71Z1N792s6/wP5H
dZOB+6d8le5LEisMC2D3PlEv/mPko/y4tegkGZ7U3XI1mQ5ndAKptL3+WE2bLKd72PoBTefaGZj0
l6VlKgSDz2GLb8k6Idjzzt3dR8CO3eVObcE6mIEtG0JOtabhc6vNUgVmAG+qqX5oX56Mptew01k1
O64Ajr4upi3EJ9xc96nrKo1gzVKtGr3LXJab8sSq0c+zD2WaxZSF9Ib1FWpknCu8gYL5JoOfwKs5
e43LXv1gVdRwLOqsEpi4/3SO5D4msxoUpWdy2dXQKNaVV3LerG0pJ3lgpmNuDVi/ME8StvQbTgQd
0RRO/HH9ElbH+5VA8w3jX2DAXcx6gB90Cv3Afz0V1EcyHmLlI6WtGI36hDPuYX4/cX8f6ou1PSt5
pKKnVam+9zjEdrDjLCWRLOK0V6wLwES1fFatxlTEmz3YO0oSJJMfhsXAIV30ZPPlM9bZUkzcuHVR
FfWhH+iMaLXWXLPi1pUXdvHBTlUVn7VES9xyvkw8iQzjZgGYQp2rCOGJigiNm0gmoOwcbqNg1f1e
oQrCVryE1UICwpiZomQuF0zXOL2Y/pUZ+zP1GZ7AI6vssZn3aCtITOpvB1WFRStWTfKfMY8tJa/g
uTanHRK4mTnxx5avGMQnw8ZC20iLV1bwE8/r3V2hGgpSgoicX4t3H9j+AGsE9ngaNmMyTZMMNOli
nqJkE09u83sWr0dAAtcXmJ5RWt1CkbHoccnrPTk9Xh4sTDGlxxPf0j10rpZrChIXSaHwgI2ZBiuh
cpN9vbboJ/eXRcTbwtxCRGnmMoS6lktwQLPDnKN9tF1q/CBwGDARbcHMyJzAXUjOxUlYjBSGw83x
Qx4CT5UTziJOXt7t2htD3RKrWUYrMB9gdmtFPnIqLvGc1XvHzzd5lI+WQ/ExX6LtdqLdRvVvCi51
SrxNdG1jW3yC9Pr9HeqDrMOaS28knBcy1VvLozfGbWwE4M5992V5d7tVB3BHPaHaqrxjfLSO64Tc
wNnw0SS3qxcBZUcZ77w1ExBi+GFvkkrcVdlsbg2zOpkbc+5Cs3FwmHY12lx0Jio6KhTax4ZZM2hc
HCmcosK3AiJZTRlnoIAl+zB6dZeGW30igT4+v9njEDkB3xTfDMJLC3tL8r1qxVxBgrkReQPcp0T9
l2yPcGmtRf7J3xlcy483tipKhHq7jPaa0tNemtRfouNTSOUBCWv5Autoicdhuv3lT+Pd7YR1ga+l
a82NLDZ9aOWOvqAU0Qy9fFPM9JK2FWSIzPqpYfoNa/jbE5vE5Hc2Y5iY3qNG7QcdTPL0zIOK8x7A
6c0i8zVDnegZIpAZ2Ah/UtxJkTPFUsMsQ/RvABlKdrUMBieq88iV8BSHUXpNfMRqEfUVu53TARPa
rOhxtJbOkfSkpY2a9W5F0CkQLEnMVsmkXsn+5+Zfk1W4qd3ACD4+4VF2bY+PywoNqCfRkiMu4Gr7
XF/Xjpr5u0QTARAqrXoSHTyN03oDGZtuzOsfkhRT+M3ZW7yzSuSYxaNkTI+8AtmQprSSOD/Q1K6a
p/LDp//Bk1Ub6iWiC57Pyzf1nnflfMA6y15qvzClZMWm15jVesw4DK5/pkX5ubWQo325NA+RhwnB
QLoyuzHT98nfrxPjyYxjeGKpFggzcaA+cgrjxvTpuIrbRoBVQPE+CGiDLR/FA3yGA9UdZ1LoM7ca
5gnKTnJQIZJxzH+Ho7cwmUx/Jd5SzVWMyLMstvTRMWfQ6wJ9M0CsvO6SDwtupnjJVfHXy+tf6cxa
uie0V2jWE6mJn43Ln4bHWEcBb57NwsfIUfM+IlM0RVTjnL6VgIDJMmNm3CHQO3chFjGxLGuXLSKx
+lwoXDowenvBao1fUdbEoitsghsTVedMGhiR9VxP0RelnlU6P6SrNXfXR1UITihpyPaqjYBXodnp
pLGSBQrKI/sL4GQdw2OAUmwbgyueUuCm6HrozshjjWLJ7pWdh0FXdgcEY44hAdUJZlNw/M41d0gi
1lhDmFSR8+1e594nskRpLAAXakEeusx/GC3pu8J/tANTHVyTiyVV6t2/Oy7uL8IHNQGaJKpZ0okx
y+nAptaFAjgJjeMAijYtUW7G4qjgkczH9+YFv7HvLWTuW31ilYlIpHscMMfSezV5Lo0UfZb+eIRD
ley3oc0GJNp08PKMrrefTl4wc01MESlloWFTgIqiT94J83QWWT/ATtdWMUo7TX9ntA1GBy+bPgtq
Kq75+Cug+wuXzr3pB/IZEWz7z06g6Hv41xDXNbXiv+IhyEEOH33acYuQIV7LKUpHgMcOK4LPGSrr
8yF/Dyp6o6yIQ2nljbl16UGubVSdG/tokMfNIyaPXneYD4/bZpYMa/spYcDq7jk7tIEJe0TzFeHw
gOeSVWn5qZCUpIGIc2FeWhXv4RYMpPDPsBMSw5vMb8IhJXiYB3hkuW40q1Df33oVYiIx8sHzFIx6
8QI26ZIUNzfG67oi5cnnynejs/HxcjOO3S4XTmZqe31E6mlbAy+mnmYGPCvyGgzRQUMeJk0Qvt9Y
0jWhNydyzlDBMW11bxDKFVMKk3VpsK8l8qER1yhYD45ujUFOuFiN/3PTB6DpxkANfizxfZZrbAmZ
ik5MnCQB7f6b1j15UNOFWXoAhPZ455CwfN/eoiq5e1r4cupzHBkJiSAC1HJFdJDxql5gKICHxhGy
ATSiWdjMsthURAKojrRubBhMh3hz5MoTftayMNlot0EHPnMHxNLerq76rlYGXgkd9Upez7YUkk+H
fFjP7pcIrs9Yt+JpPU9JaNucp3YPsvDrbfUUrKF/9+ax8frhG+WH76SMJ7MFc68Dro0Ej2BrX3a/
cxhp+L7BTNv7QgMMPS3BvK/fVl1WmipEEgSN/sNCQfMcrZ6pr5IPB2VDDcsmQBg7PrTQ9TesuURn
4bG8hDAjPEbQdmELlINBa/hbLTWxr+AMcTqSkCm6i/MIHZhg1ob//EFQ1djHnvUhXE06UKO//r5B
MCnt7yKL+OaB3pHj6q5WrP/8+y/8msYNUrvxbBNek+OHMFlpbPImwCsQIJpiAtXOvo+GKIzSvj+5
MOyhZjQ2COL5bV4TNqzRFsGhoTFt04dPgYqsDYHYHGLd81+78FgToYSY+kwHLYD0nPXp70GrVWPg
SL6ZCjHzfpwWJ/efTXofzxyRBNEZxZw7eDC0nYr6bvD2V6gq8i0dVhZmrbBFq9pX7AoMOeR48UvG
FJns2lpWfvrHaZCaQ+dnqumOJB04UYtWydGpC7v4Qa25YylgVHKUvyi/9f1oXH//729PsII+4rKg
jcISqJ5Y9Xdo1bq2jxW+fxa7mTABRg02nzBD+xOi3gZ1eHdge5pM1sZ5nRNYSQ45+kxmb0IzBpNT
V3bpjNmxiqXZG5HY83G5dz8x6qwiaf+gUjAy4undpuTYha/YWrvwxg0yvjpm2ls3Iy6qxk0FpE54
mfcxqnUTekb2OfRBaun8hFZVV9twpsDPxiqVrGv5PuE9GzRhiA7eaAHQbJjcsEd4l2yWCw9wyyml
FhnWp98BuSx4v+mAifCFNpn4aQtThZPF21VUORZsR51Hn0746k9oldzg1p5HrOs957P0a+E/yoyG
sBKUtgTox4POA0u0rGJAsIL2YPDYrCJb4jJs/UTRCi2aQFNlzavXtCz6r/tRo5RMbR9vgjVPxyKO
ZyjDJkbeAP9xledLLuN7pMN+kAA2nqTlqBR3QHQZlxtw88MFPTfXp2MeDxnSwaW4ciRz+Mq8bDJ9
XN66VXkZrdhD9tYSb9wKFKl5gu9joKvDHj1dBsmwkMMS2336JacbUy7XZTj7XN4ORTLAzt4zrSDO
BHBHHPblviheoAx1xqxw73BVs3sT/hTFxzTIs0cYEz2Eh0ftxB6yXas8qd3Xk/p5hl4LWzg1djT3
DUcCwR116PCkqQaryzTvKabhkHSm/nN0JYKOesKjB8EfQmLro5FdMf7szSAiCECIGok+vPWe6esO
+3SQE5VVqdGc5jsUgnfJaxdDJFnImzOEPzhL3NhBACiRsOgg2L/A5/XmlFh3HTEeGjL/CjXaGfP3
jXQUDx2uHV1z6UcIDEqXDD2dOrxeQy2kw69rHLszH1+mPoy0PwZZd3xK2V/m//kZRRY6m2UPDvk+
+RnQrUff6Pgj7zxcx2BMH4WFUdevo82q8TQlLpO1DzTnRwWKC5+eaNMiKGZVQ5AwJZ5S9+hgZcAG
Q1thsvZa4UvK8pDGgYgRaz9RDIc+5kEA99YvbWx0u5O9bymMnLjMiEO2IEtxf7/ORnDtgLTxedzD
tnKMsRy/Z/wzMyUIlAl3TD5KeyHDWJx5gMNUyw/Fm0uldMUZvopwg0mVhrpspwDZwnvS9u+a/Eyw
e1HavnoHzsmeupR2kXDEDHfRl6Atspxp/3sa6uRZvngIYENnJCkxaQ5OsNWAfsBnTFbYcefdcVw+
MzvgQxuNhURAElPoLOwIEfwWoiivEeLsVO02/JN/+NufI+rFI+w1PZXlAzsYLSx9pStQJv3evX0q
kg9RlN9AOb1oWnhHc8Dk9PEhkObYaGObIEuHGo5BzUTurPJfA81bwNofhmtaqiTy2vhl2tmx0lXb
5lMyJa7LOuQTyUwQlTlU1F/vZUOAjjl+t4JdT1vECvdIZynMtxFhZulngneWW6C7TzPSaTWGlB5w
nISq0VaCDlSc2L1zAYMjUeW0zltVG5JwUOY6TDIiTHiwefMiaGUi6s0L89LBI8rdu2PIe89BWEl+
TTMCmyMVPYmhfWuNLq/zrFSmWvVZBr9HzyQ2THUgamcX18k/jqz+pghfQBsY02Locp3awB69I1Et
sTuWrA8ME+kwvSPlNrV6L4/hFwLPeQ9X3osUvl2GhSphAj0ZjRcwps2RMF/pGYZ0dUYjrls+W/px
G4l/azvAvAZ62RSvnbDs8pazSHh3EF4dNQbgLELqm3P/YY3RgnUpO2EWuZ38w2ZsMeYotNGh5Mk/
jJR1W8q7N1+WkG32evypcCR83LPSrDHkna7nWpTiHesNYHMrMOTwsKINljjb+sBRu9tncUZ37NsI
IW9hXg4mK+FD1LmD2WGQoz1ragFR3M5f23+p4+A6uWpgfuZjctrJsxw99vCRNFr6yirWW7X8AOL5
rctrUFYtulSF43Q+nqFSvctwW/rRNWiQcVxFkYYhZQ3pdQftQsM5wCFK1ObOlQHaXpdj5JfFHz9Q
ExmxSj+EdlgJSIe6MVXIqEU4CQvwr5U0ti9Z/XeoYjUkUotzTPRR2XPZB6zKZhUIigGyfXNBsBcJ
+ecpaWuBTlm58+e8nHYHGnhSBIkyiPlXc8yYEo2hQSzeTog5q87WGk2lnwGai79jL8ccs6619E3r
G9r14JE/WPCXYRb2s7bgBmAvop6iyFSWlK15dZFxh3dk2/N93vAzq90yNI45Tngm5FPTOPlASG/L
LnKn3E09OwKWa1bS2OoJP6Jn4sd2ocQhzdv+qJxeWcxDcw1Awct5RRrs/6Ylzxq8veY5QW/7lrr2
+xCzGLqkd1tRRhdsQAVHvU3Le6MDINEEMeIlNGS5oDDe6WW9VgOSg8CcvN74sFWDSmefmXJHQOFr
AU9WGEzs4BtyMeCE0HEtgmIRl4qdk7SOrSl4ETMIxEr1GjYeSMr95waz3N0o1nTb/1Ok7w/GHIYy
khb7ZVDQkxne2lXHK4tt3lEei4VpTkjcadNQKKcxOjsRW9KXpO2gp6fpcMpIUAkcmIZMC/82vFXy
BUJ9p+FR8j6CQUpWwXMhbsHNO5bMMHjai698PijONzizYGYLvJNhh5fRgRyiVpVxVGDifInbKKoa
WwaSfnY/OayopmaE5qeafWuFhsReMCZ2DPCJq/oK9idIYH3dacLkRiB8M+uwn8vP4rwrLTpGiKbj
h3S3tNrmrknsy/ungbG6OwtLGWR1rxLEJhaxV0S0u1kdR91whQOcEGXrjP7AA86h2Ei8KNXMtIAq
f9OW6aGsyECtv1WV1E9laV8QiLwqpW6pYvxAAiDijOevVdYTIsRhgzBUm0g3FX06INo65OUmzV2X
dnBfwl+vG91wYa94BIG9deQvwZhKvGlxyliiG/HNWm6HkqNRjQN5vyLndE+AxRtX+wZ2l6PzMsv+
r6Q0jbcZw84VnzVERxi0Pv7byS0wPsN5nlC6jeyEvTR6RrYjKsk7qAuTv6Lcq/2KmNR5n4GpLtjj
x1geGWVKJpjSP9z12V4iI4fL8XpSiQkhIWbDR85a1XDnw4brbaPd6QXbl5JFZaMdn6y2NAWoCWZd
6rL8n8O7WDuE8Zn5cvg1HwljAV/vqljpY4JG1w1PnR9/r5NpepT/0KO7lwW07M9uRhyVCeAG59ZS
7O5pUNOba3tKOmEWQzIeQl0vU3pFCJmPk1rQp42yeFh4V7wzGF5NgTT/74Po2AhUqFZTq0c3m4Jz
WEAF0VBlZUOnVlwOjFWWgMiDZ63OGlQmEhlB1bPEkDuqTyTbSngrgmm3AUYJhreyAQMP+ms/S1uR
6WmEVNljlA32nIVhMIvgqhXopc1LZzbc0UaDeCrJ/lmuzg2xE7rdaO2OHguC4NOw1ovtKIAUXM37
ZJ+thLuGI3Pb5cSXoHm6vTMKvsL4VJGOqewFhXaAsdpqeYnOCvl085Ivzc8Aoc43Ql0XpfIZy5ng
K1b5fRkegFFsljhoTsnEt3f9+o3KLWE2IEm6lij9wqBhKPs2dUnH5/h66edRlX1XT4RETaNYo26V
nn6lw5E4YoNKhoUe9FqMBI1DA9awPV0+SKMBmSGFUF9OaOky2sYTRhY13nYoaEEbA6L/I14uCqNy
3TZaIgqmNHOqGs9/ZxlqPK3cNFmVQ8cy0H2699R/5yyVraE8LB0tlhoKvhHKMkDRdFApfWXJNU0N
IfXCtdf/6FApvyY+7Fjp8FQCNarH0K38gjoZR41itabw7C7r6Z8fqh2uS/CoT+oL6ooqTBsaUVyk
xRAKzMZt6mlgLu9gxLAyDtstqm7162QH9npoktXORXQyBf7ZoBXaUYKFqvBgr1S+aq+O5YWAmJ+y
GI7mpk1X3ITiZmWcF5VCi0hJOOdGkaAs9KOZT4EE5OGe5azX68DqTYNLNfS77TorruHqMy6Y2g6Y
gx3zQbXDQT1ccSgGbkwF48B17J0zL0qKcxOP/QgXR6HAd4CniaP+ibaVxOYyKIs1+xpy1M7IGmvq
iM2rZQ4jmLAoEIfSse1fX415sZswntlC56F4tzQDLcpd13XvBFTSV+qdPMShkG93qi3ekIe+jjjM
oWFfvEdBI36dtgelyGrLPd5lZr9TEIRtJSeCj1Y3n6OjklM8MOze2jMw15rx4OWdJBz7UwwrB230
hLsHq1YeA8U9S42xbaAtu6StIGy2ejdKtUb/GgV0jQuhfz8UsjT3ipo4UTOPoVPGBZKjra9fL20f
j633NMn2mIaFt073cgQjEBTHM/frBZibCOl3VuZhpPOqpLTxNHDZJA3E/mUjCdfcATWaDwJOCmzO
5IRpRC8UwEz6QGmZ+blO2eAYHBBMLIZT1BFrELr5G0Xl2b0ARWP7eUZ2rQ7mepwE4esPhc3vJw1H
jRpIrjdrqNUzQNNJqqfUOPclNopjUplMDWQAmg/5YKxRkuECLOFTe+RiuE8PeNTfeiAQYgREJcLi
FNYuM19J6FmKbFfUzaOMGjF2qGp92IAPZJHSbKmiAdqW/Z29F1/9rN3rclHT1GaI2KxUKAJ7Duvy
0dKVU+TdqmZR3c5WdjJRaemBHSKjgnH3fHGOsUBzQ+MoUEkpCpVTWCRHehXqS45J9uPDddwyNC4X
BJeEdoWi62dR2MlNLrt4PsKt+4m5DiOZrTDUOXkTY78HtQVgPXvUbeUSlTIBNs0BUoiV7DiMXqDy
31Oas2lSx7jpfBDvEeYTfH+PGBw3+JE6Ad0zQp/yCMpiaPXADe61rcGphjrQITv9WKi24RoeMPlI
HL476Tup1z59lB3kY2TTZGP0QLXRp+rurntxyRZx7TJ/cvYsx+D/pJzqvfed4udDaRmY97Jk6WNR
zxekI8wpY8S2aprJ8iDmEPk+B3PtKFygTyhISCd8EY+fzaBYB0InBhg9WjuwXQRG0a9JBl+8o/KO
QdPG6G4b1njNwMDVHx7PvQ2F6TSMZ3jIpsbYFTeetp4ftgxniFRKf+UQJJtkamybvPdfEnxns3lS
/YNdc6Fsy/rpOHPz6Ib/SEthuSe+50qK9sS+9w3aVJCmhRWQHcF1hw29YBXQ5mRHwgHWSrP4Xask
T3NoZiY9pPuky4NwZW+AZsfhsUZDMkbafdaCwpNOinD6x3GKjtItzGVZY8dE/b1nnLj3dMMcIQi6
PqGAHdjvAodHSIJNFmmEHSPGInJhjHssx/BnyPupEHPpZZuYuziQDOvZtnagA4a5Sq9iTx/rs2kW
cgeM944qJP7q7rXyc4cr02uzaka+n1W1Xcsi7rPrPKQ332EU6I5CQIYVebQF0Sm/pyqoban7cWhd
VUkYeT+Vrj3DHjHrz2nVBQZddZNOFncgrqdz/uH6atg36QtiY0bEYyNRju4tmioTAEYeu9c9UNE9
nH0JFqZVJK4HLuhKcC2EUjPSOwoTB47NDQw50Cd4FIX4yo8iZMpfqq0LDf7rWWw64OOMPpn39itP
M4PACAbSM7cyP1QvbVHYXP82+cUcNjGCiu5inCwJgO5gr3fov/KYWzwRhpivQfB/ErkJp9MvkWvb
H/+bls4YNIgI4EowWNhRrLlurK7xSLGf1IfLcfcUj6cEx11lCqvxAYnyhTsglwk66BDFg/HInhQt
/arKE5oLcvVfyNib6lM7Ec8/Sjd7yCyH07a1jmEi+P1GARhnlRyrlHMWn85ugslK5YOyasUNNad/
Ehv35nO6NUXWbQwjYDJytHrZJ6me6c2GdM0/dBwKx2Pq+pUb+RP/9PyB662zQwujxtgTDd4YvABq
FabuDgEvQwpw8vA4IwDsCAeMGqXHsnxVW17nbocwBukU3lNB+7DZ29dTJ3QkgtC2ycy41y0jTJbD
L4iviRosNJOtEEyxYWSG0kLXf/jYNF6xMKL36iY5eJvkxPGLg0zWpWGdMChJ52zJU0tUcolJJjlK
2Tt4KWEm6Z8poAWyoSkFuo3A7RRkIJEKRCifTmnhB4egaZL8mffXoM1K5wgfGcnJ1I9Lqloa71Ma
m4XekXG8IvF7b0OxPr3lOCM6KQmyZdPP6TSne1jexoS1NNZy3NJztsw8x/K4LKev0w2mDWN5obCC
iFq9uUD2/SLN4rptNe4OOulXnAGHWZHmDQjWvoMyzkXxBSgqfnzxAO4G/YOJH+o4Ge2jGV1j9yIF
vVEME4thCgCtGMOfgmztbwq6XOk7AHnbB8NIFFKKDnynwtJhw5VETczFaipUwEfW6ZVwVKJzs5re
aiWetFNffA+4fXayLulJsartop8XVh2+X8H3HIws4WbRDgg3Iu9eqgvTKII9f8djttHhgb7EmyKi
GqP7RWk4LmtAYFT6aWeQAiDh2Bga9QGgnw8zrIxWahakOpGnQEIctWqqC3IywUrV/nX4/vKdfQ18
XjyS023D04/cpRu3urRSS2z+0TbMwmAJQzYOsKACk2TlSqONFYlKljbX0joYuX0JNkhgC0J8JfQD
DUnYOKe6NA7ypJ8/QPi8WvH0vCcyd5Nu2p+MZDrLU9WmheIwReYWrO4piLJnWe5KWl4FziYKEOjC
g5Brzsn5XAUnVrrFHyTJwQe4eE9zralbGa2x/BjmH3bZC+jCXlSMzrH2kBaew/5L1kHmndoA8P6l
Zkv2hDV7tuus19sQIHFnhJaAh43KTVdquz1NNUhPNCGNCnEgoYtt6CuPkYo/zRDYsBxsr40oG7ch
VF5/06mzFOyRKQNQ5xQAHxcJWbozp9uMv24SshG1N3ixRhrXY0BkCn3pRKH13evfImSelWTjOR4q
D0XtkLHpRYae7O5ENRznZYL7xy6TDffyHMS0PrJ4oyp6k9dclbL/8iccjZdDuy7VSo0aG3LUKx95
0d2HtSQx0YEIpUhNlH80KzuqZmgbGX7f2z2ZTbn03cKb/aFrcPvcL5GUDox6VCu9qFQpV1QwM0ET
pF+pQCRPfaWl3WpGqLVYnXuhQav3yE7lSXwHrL9+Ty52TlPVz79yvhGXzsFFMBeRlOX4h1WJCJ8x
PD6LrWfWslwjwwvXUxK18wRNZ0PMaHApcF+bHK4Lis60zfbR3YsBKtiOds9KUKOx7h0LF3oaKCBc
VCljila5yAYdD2TX0JiaHP36VOETWUGJcg7DP2Xx8A4TlTndFsx6srq15lLmoYFu3zIWL+jtSU+p
BRPMfXRaWEzTlYkMmC+mPPTJO57jfWDxBb7nAEDvDJocOw9VRGRQ/Y41S8HrPHYv+L4UrLrjQ/4q
tfVv+z3raY5Aj98UWXmg4fqH7e4Kzg9IQH8B4nm4QWFpKYgiPBoIlnDJl5qeplKWv7Wf2Kwy5+al
Cd6JlFxkyvGJlwVyumAKbLUdci0eF42+2nn9y8FuqxQOd8nKGS7d0w8ypL/oQS6J4wqWI6rgceIF
7SVRfhlObo6794I5OEgbncdKTEsplzBvLCzKdno8UPNFFKJ0SBZIZbdBmLNrZoIJ33xvsByEUIGD
NfIf2vkxj7Mh2PdxUJwrHz/5EItIzbXd4W6gH9GfaAnXIpnXFSX9UbKw2EG00EjJLTNiiISiU1tH
amkf14Preg0qKw7SDy0jIQEyxho7pbQLB17bDu0imL98EsFFxS6zvgyYs3qrsCmc7cqRGkhGAWEa
VjeUHpMCyqw3RCiBDoxCdn1VQiqzbCsLuovZlN/t4L3H5QmevJUsXMwFGz4NcoS9c2eW6kYIyRt5
vbyPFxxiV4PayKjAfH9VEa+o2BWxxgHHqLex+wRZZk/d4i7wcL4oORlyGItBhgm5mJDm1kRYlaAh
DzdM4wQB4ACJ/ZPOF+UWgrzQuqIj+PTGuVEpEbe8KC79zRINg0SrHq4IvW6GD0hHKBG3mFza39HJ
JDPeu89N4cd3nQ/M3pf/sOohL4jIO+dLFbnbKdKeeK0DSwbT0E0NHlat/1tWftp5R1HASmQXA0FN
DmY590aMx8SB1ZngpCnclmC8FV9mKsquLzT7bA0gvE9DgkrMlWc5jrcLq3z7tBY9wlll7634IHiU
6VM01huw/fDIp24+BrhMD94tAxyOKQbsi6mVlFDxNMlxArCyCVpyLHZEG2aeKqZvsIDpUrg/yGml
qE/7C+JY2Txa/BwLER7DqDQohZzHchSpixlJO4/bBlhdGMDtk00zmoi1+hj4EmtOQ/OvTJseFFji
2lVx5MfcFY5w2ufh/Xb7epP9OBzOTdqWqktq9guvREDrlaOeXj5gJXQDPBsLRK0+WD65QadpPKX9
dei931jrEiDZBD/EoFmNuh9f94tC4J7evRPcKvvtPc3ggCrqSbF90IPlyltGYEucnEcL1fO5QzGB
/6n+COJn1kjGZePXYLo8wWZpKUlvd9yqcJCusfpAZfsNpxq/HcnVS/JYXqjvWoAgO3rwkcgLRivv
Nfscmnl4VSx489kirKQxp3BF/fiSHHC538m5zm0fJ+YWJTuzTdDmX3ZzbyFGCR5eLG4EM0xXFKc7
J7n+SEOgniAS9wFbEDAW9kMVSBu50d3nwDqVCuqI5OLhZBW/kWb6lh45GpTzfkFmo6gkwBuc0NtW
ui3ajR+/uOrgsZ50xzuIaVCXJkXRhVORibI6Q5e+DNIBPHj8Q1iHACWzLar0tp7B0xKW8BOhnDsK
AmXGg1sqWghR/XjhIl1+sxIbwPtz6NM62Pzup3ujh6h8HxmHcXV2dIMBiPvpCnvBYw1EEuODB61s
OxJTxtAWhEP7HAZ76xY7XQwvpvDe5ksfDUHNtV82WyU2YP0Hxd1wm6B2D0yAQCyNcpmeLZrI5Iwj
reHH+BwADuyzjnZHgmNiN83sXL681qgtHt2moGvWALJIQ5X2GvNAyjF1y/dWBn5qdLStDOGaWs6x
UoiWbaD1U/ApdhQ3PjhMxI8aoZjFlotmHn7sDBbvGQkVjO73TZ8BxmW6ylwKw+sCKNPnaWVlcfql
BdyZFjfCHHERuQc93J4kWqFhaAWbOXuS0YabvrHTYDxkEQ8lF4CTVt7pTdhseCvl0A/Exx26uzVc
racUBqKa14sid0nufy7amieJLkU3FUou2X0R3J+HVOxW687McTgOZKwY0dVhE2k90SmdB0ddkTfw
v51u9wg/YqlyqN+Vi19JiLJ5fiOLIgezqpk0eze0DYXxDLCp6dwvoucmO+cT9yBhC5IEfWBTrKAb
9uaGIvNXxB7M0zXJGU8sRFni9iP9BfXwuWstaUBz+/lKMJY4zFU+dz7SEX1/htFYE//QTkDS3vI9
wZBSO1na2pHeopljZyGJxeASFiJIj85kukyO0W8uYqrUVUzN4j9JHXiQ5yV82c0Mz2tyH3XJvKcn
DbPGkLz4gQIJq0wWRDzaXpuNs4AjzXiJ124zz1VWy/C5Q6Q6h2mM05Dp9xlBbIv/nrfvu4Ja1C3C
St0mJ13W/0a+Z4px8/UpXyx2StOr8pLubEP5fvT0ZQuL5sQ48DudpZWUybUEBhD4LjJpSNDqfEzQ
4vAlquC/oYWszgJd+PgHYUeLYalPbtDCVWwyxQKQI15WLjrFQE4kfdS4SgURekhtzw0jV2LTPamJ
Ogbfyx6GAaw/RA4JiG8hrS9z9Z1efreZpGcGdtqgW9y5gzOW37TH43WVHMzZJfJnttNoHXmHqYu0
VazP4gCSf+OlOzb5JTrNvWvacixChLHIJQgJezMJVGhabmYbnI7hUD4lbReCOIUp4il8ByGoSWTl
WegeD7DQMXFGIE9WM8dbRaexCRv0KppnR+0l3xp373RAAF/cfqWuVVTvnGVWI139ctbh4/2ciLsK
S6ozLW6EgGCr/Gk8ck4CM9PlQI1YPdJEVEIT14DHRTMhIuOwuQau3+T42bMsAkRey7NIpjesmcDa
MY7dmvvNFTAI7zD2+hZaMOZv9B7z3riaUVlQxD2hHoBtddB+3N02QSLOcrCQo5dSAwzmg7XOj67p
1xdyR57rCL66Xz7UBJh+zIoIAIjlDjEZfh1/VbaoGMtMbB5llQFH7q8MBxnTaGKRnowa4TPAvWJS
9AGSw1IGFpZXK17usGm1IsMjqNM9y9ocYwT72AJqtdb3UFHmqbUGlDF9DFvJtsKAVH12mZ1QFfs1
VKSkhPxFn2PU9tUNtQ200HCTAsohY2KIk7oXF1gxXKauuFsEOfFUCcZsU4DZ06Nnp13G6AomgCph
su8jUzvBKEpnQFudbd4IM/eIU0memTVCzqXVlgNQxRQjdRtPASC/NAlA9JzmV9vIBneXYTTTpkEJ
+GZ6cpG+W5e63CkVFOQj8XNQfT2DmgT8KbWj/jOTUQm9C4Hr3mWjQx4kJBj0NXjaVG/jNV2Ubq9d
ldiINxL7SO7fHe0G3/EqfAiVX+T1s+L1vJ3wO0U+dnRwAl3lv8pveAhyovPo9CtGVGZkXtp5J48v
64y5R+438OsNzNVHotGp05wnZtUdRvnyxR1I5GcyVcTOiEwzpeavUyNc+XKSy5jGwnZUENv2xL52
3+aH4ecoWcO13J0Y1bjgkjPtcRPJ5xQqtwoRm7dYeZojkfBgI/qHrJvnPZLIjUvJfa1BtPodrBL3
jnvKNtFYlbsT6cKWn44NrTzmmE9D+mYDQCDgX+p0gNePWCN+F3cRLAqA930ovhCC2v25m7n/JMjp
uFzkNdCagVZiymLOcH7QsZulyT1verVQwXkHGQpyR4gm+F40TD1ef8NccSKnkF74BNmrqVUqsQiL
rMF0zJAvbsLR7Rm9gjzOagG8OT2/UEPYo7xScN0svqlnmWSh0u2QCt30yA1qJlw0cXDoAvIKid4D
eQiRjBW0/f46WGaz23MwbgPFI9FOU/jIgGjMtD/BQnl5sAOo9MaiNa0PZOWFfzGueyhhDqrUh16/
V5L6llFwoOH60Y8F6X3iF4b+6Bo1UscI1Rm6DGfuzOB9dhqiodZPi/VvaBYY5zL/Pj90aOXeFF7t
XEMAPjlBdcwHYU1D9yh1gpH7Kq1tc6Wl0oyjqJSEf+xNQtB0265Aa/9E2jN3B4lrmHuPher2q0Xx
N+Ncd+fPeruEByjQ+Dq38L0JEu+rKDtRFEz93zVQ+3+MmE2ZfXBSCST/V5Ot2nefPbhjIXCEklfx
196RmgvUgfE+BcGbBEV/mdqt/GkjNIw/HMz58B2Q4cR0w2XWHSfXmCL+9V6jVYixKCxlOf4164C9
d6hnsIEyZiyVgsG54pnaavUIa/E/nCo9Uru+KB20onSMTKnCBJpuuYQQ8S53zEYjcrmjQW03vn/O
xmg3VepVa7rnjBHRg5IZPKkFDfP+jnoLZgE5UoAJfLFkcIPgZ72kbolV+oilSmqCOcg0R0QzPNRz
j20FjChOcTXCYeMUyzHXnll8vrTKjkblKLXa+u7lXe2G2rHg9rrZRMwJmvvAxxpKF0fts3P9YnVn
OHX1PBbRfnbbxjnEAb8GCWz43bnt59rRlojcqOVqQRlVDH8RRyzDfHSQknHj6wHPLbSYIbYbxAOw
5xeefe3mkaw3RB9nkm3w1abnvRW2eiYx2xA15/+6wNeCswQbI8HtyRcXUr2GIW3Zs1vy5vpMSSDn
VE97hJ0WY2p+BoNe6qF/cLcLzkwJlzNqHId2kZ6728I3tSBTV+jf7XwhbyZYzPUk8BTkNcVxn6WH
zNg6ILtM1G0TL/W3dD4LPkMKP/d+F1lP07+BdL+mrm9cMTkcmHP12zIsY1HkcAqPUhv6xsmtvhcW
7ek/OIU1X5Lb3ZDpXSpTtZMNkAObitpg5vpvyCn3MyK5ew9XUMK6fwFcMUm9/h6HK/mx4hhg9vdY
8YvZ8OTwstYymDeZJWx0cnW5Jy5lGh49Ar2JI3su5UZNP0HcWwqt9uUWkAgJtnKarbbEVUpug523
iUdPkGQk5g7QpE3YdCWaigLKk3DlYaDIjneowdaiRn3kaDLFFZtydg165tqNnKzG4bab26qFAoJk
2n4KZ42+4BO78ofZegoZLQkfGSMvrSJR5KzXSScbmZeusCf8p75U0UQiTlAyDJB0ajfIbGfvNKdw
Xy47ChMNP3D0gEP90wDiAaSlSo1yJfAFIgTxQqGbJlv8Td17d7Ntfj6voMIfm5wddf8dCBUrt8Kx
b4iNth/k8IAgE/TmfE/J85eMPx8LFTDMZ9/gTGd3oxC6QsK3zpgYFJDrMs6fb4S/vSkBjOqYW2ir
7DeS8Wg6Acs4BJYrYPgLFGTskiT1H0oLkSOr2HPqqaZddgHSBDXLQjZXQpe2N9lPmJ1TMGqaGIQ4
29n0VqTrToGSzk2iojrs+0os1/TyaXcy7OQYBw75r4LirnSAYXBLS2dkmI8N6BGm3f+KZIFpCYXb
ufSIHj5euBENd7LuciawpWLU7IePdSFisxdIFjzjzAwYtVUCrJEmfkxMfnjEjEe9vgIonJOU9aNj
IeJZ9ne8x0zM470iCexBq75BRYF1uSmS9gMvnuG9oSlldfFa8B1BWvCrflz5YCUiAtz9TXNIL7hv
fsftwW/5R66JA0IJxgpUzs912hSXK+ZggKEX32EABRavMoqvj1z4YpFN9y/InhZzpSrLeD5nDNLT
bRFPFvZ8QCR6MpuelbJ7DqVQpX9/1guWooCLj/spxHESVgXMglhGjebsoPDzjCcSaYsORTpX/qU8
1gg6WEenUUk1MiYgpWt+HDWAsH6D/BWI9w2C71ski6ETpU/a8PpyKz2lCJ/9ImIQOf6WBiQOSOGu
olaKBe9hKpHPcUVANQcPvWAOiph2o2YIVhUGJdmOOHI4t3kf7rLt/BYsoBHmxIeEusnWEMgGdHzo
mqbFl8rD0ZyB7mAJYZMTZoVkeSZPdlmghWtXkRMc90Q9SyJcFIccHvZwL1mOrDTvnpp1KMGav5hL
NHiO5dG0DV096dJHAjr3NO4eLJoANFkUcmNEVzCyBY1QRCJwd67Ehpcx9oLh9IkrH6NzYPMrIyjd
s4VC3+zv9FQy7htk1gRt8/TMdy+SMJ5ubWAlrYOYwJh4Rg370ZLY0zJb06bSVMipwc5ekdtMafKY
ndPU6f9VJAMcgWk8lOcW82uW9/ERvbeollb7X/PR4jyMOlNhCreY/KBp/7hN73A/h7yFH2YweurK
6Al2iTbFJiQR4cZSPkrh7diqIAk52kPcNpEfuPx+YZ4GUk5ifTgXKSNWNRq42tf/9UKuJrvQ8iKf
tOqf6ADeAOwbB2EvEh3sD8GqneBvR/0x4KFy96NbeluRxCH7cWLTp6fP55/DMbbH8Bx1IDMGWwMC
8qhpnQQlz9FbOMQS2xz/ptdDwBsXm05vm0FD+3W3vjGF8hF7zVzGWZaYpA3mLT8UC3xOoUr6ipfu
n59N9a52VO8n1z3SQXx6LCUvWmCG0T0r8dPV7meaxdb5aOfw+LVY3uLQZDWvC1fXBhTpr2LfHlxq
M6w9w1QDezykj4B4tiwXQ6Ngek/bRPkDKiGCjo9+HamvXyCoD+6eEIGKZgxapMWOSQqu+4kA1uZE
2D5n7CZ/rj4wdCtUT/bD3/kLaW7hsGJlHcC8BptxyunHBZKzIgrc7An/Yi07Bc7jLIwqNvxvOpLD
NaNpehuKWeot5xEHtsjjR8uygch1sPXEXCAvasamNYlWJ9WafPzoKpEVIFev0jafv/643N/xYVZM
emd+zcV63iL8nrtkdLRyAXaFdnAItm3a+QJiOXf71KztnVJJbqSDD9KaUTDLCmTZKDNSjz1+i2ef
DQvhDtv9/OzJnr7dJmxpbEl+c8QNC3+SpV3hRRd/IInqwbTF/ZR+x2zcFEnV+/7MlGk1JQwlxi90
5K9ymkMtGlbbAzmZ9WLPOqgC+fmhhA8u4KHtQmgmk/fwo4R3MV9J9HG9iJjohdG/Y35pLN0tkKUM
hZhGqVA6qqQZxi2dao/q8Mv4/mxjT1ACu4mNFs9gOY4Ohn45p9PolpeOl5Awcfb0Ar9ufzy97N0A
Y8RHGRHyfXbdjhkXsQmoi1ee93db5zUD0yPG89NqfdwnCrX2VUafVjXUrc5qlNePxLYZV9GsB2QB
8w8KijpkquRKW+u/7exiMMxWECQMe2lkFFDrA0Um1/n/6XbM2sHApCUWlv/NrGiaA/P58c/Xp9Zb
JClOfuwEgXsTh64OPObaCwcXrv8jxCAMG9Nh8FRVvLUaRyqGF++mveIBVIiU0umYm/Y8uImjWA/5
5k0dZwus+jUiNMPeP8swUbwGz4JgfIq0B4J7WtjnBnPl/BPyeN0Pe8kmZ+r80vQaMKiotxNzgqef
LOmP8B3PkDgfhbLGZBp/WI35hJbjFjZAVwc51HSwQQhN8Rav32sRXwgiMN4CGM6D3FJgcWQWOARs
z2CKQdy6q9mKmGxHlB0D3gCxoklOjzHU7D/Bj5/rzTzW3TB8b+r44XG+pC8sjQF9BOjpvQpdXBXp
eDqZv3NdAhsXLznwPhH/NNlhNRVBOw2e1OpHHE5UfqeP1I104nOKTnnusehis1wnqMO8COJSn+oM
dIF7gB7vztOYOpGOUCDDNQvf9QDKNEuyfatjZTFAODd2SyOLRWByuZcAMMy/0jX/HXavCWLMZYD6
4kZ6p+dVB+aNptIlWKC5eSObfN+fPkNpIsL92R+CeAvdboCplu2ISy2FfxG4m4VKD861mVutmSl7
ixbCeqYc3i5sNfoQ1hwsecATMEHMzSyNZE3ZSfa4qf6vMAUiMOdLuDpP7e6O+cj0lF+oDkht4KlK
PFnxlRUp3mJjJJG53KkrAiaQHQ4CIAY60ndbrZcqYDQvW6t28jSM5XNMSmZOa6/BCXazqAgQXMLy
vS4rWFFbCgm39wSo46yY88uaM7l82IfPL6LFMptdw8ipQ6EJU+NYbpLpK9ggIea/aDBAI9e2frC0
Mb5SsNKa5rakeNDyXxKT1BAscCBKJVU4d/CrTFruT5Bm/zfs9OefBtokSJz06b4HuBA4tGQv2jbj
7thuRl5IYTMJFfVhFSdFR3NnP6Ja+EsI5oEZH/TGKfhMV3WppDVSSjWFwv0NCWSF+KE/XiUm6Ctb
tFjdlAQ19ZiGTQb8/7mBaez5Wkaq2HwEHa9UTbMrINfUIlKAOLhz+5qF3DsVbgn76Z0TNrXPXHiQ
ArDe5e/qfeXPP24UrXBrDYYdABqtsVUBpYK0Lu/uiFCBZ5K1LcLAnfz8Ok1r8vMGhIaRBm8DJ+bM
5E2BqHG4agsIEiwlhBF8tR+0hqygrP4IhPaQOpvHOLXrjfa1RNB30K6vTC6rDkKVxguCvOyDn7GY
wALwnrUjTTRHxUJCHiLupn8/8zuWWZG0YWeD6i9nHPnejkaBxi8N4TiqfKRUX6fYfItVKU6uR0Fp
DSQovRMTwXv0tp/F1QfWq5ZGUXx1V0YN8KLHwVb7biClJfltPlQZZZmnjaHwiPcGzvG99Q9OMTrw
PX1xfVwvbeIB19PRdjnjTRpep4G0Gp/gKFvKf+qiA92w4/Qeo2FWomxkzmddWZigrOofMX+OL8JS
CTnZVv1ypJJaXWxBHTpsyVqYzv1BsFX78oH5jcGbIvzSBEup7hert6AFRwmBccgY42fbLFyBbFAl
vWhT5Jnnq5sSi81jsrjHa7xgIaJfHARYdZ6AAq4BX8JKphbua8GXWh/Y37KTE8XsRsId+Hyi/Yol
6Q7TvSQwFlTFcXYoDLtV2HEtRVPvcfmO3q7In7u1BfUFaGE0YxqzDtWOzxJhkj0euMV8YBUuhD1C
ZcT+E3MSdqcDe415+y6ZXQswIpv3JhLnFPeOLT0NfsKIW2ELKTKp4mF97WagMzrNSxyGc97tUjpG
EYLrUABvjyat7GcdxZzdld88NZrOudg3yYth9bz/6YuZWQe9+GLwZFZFJqgYquuyDFgqRhEfJT4E
z4u/EalASeRLTPNaMFAwPtRmwhPzB6L7wtotiK5wsMaD6ifADbnIKzOnoyucXuT3mGC+yf8FrJxR
dbRNS5wZR3h54Ge6/VxpCQJqtkaF7AueIcMSGDrkb1PP4Xu+izHsBkro7RRvqMuZpgMrD6hRidMq
sM7LFQQy/HxK8gxwvb9j6KNnTarYevzWOxMS/5fYI/kxSit53MM0cBUFmGKGkMakpTfbOfhks2gs
Yf72e/J0stXWyWRCGjcQtIvSDPqB/Fs11vMKuGmBvWXCnEtGXLbHnE3qbyhIlnyORljHpISkzTLG
pGY1s/4cyHJqzC4Fd1RF8tOa1f6HOQbVv2mz55Br55sex1c0O6nd/vuiiUkYAFhI+VScNYhYbYiG
oKtv8iICU8VfbTuNzDo3E9ckop8Rms2jJ02KTdpvqAbc1holulkvn9kwKA/jjaxlvnqHT/mWRKBX
Ro00fvKuat3bb+p50Y+/RAfHVLRQjGxZOEJNTO6CGc5Bi9QtjAba0jcTEIwhISXnK8L6JgwfHBxU
BK3lg07NnlWonDRUdHr9iaX1Snd0brCBml/Nk+gQCxdjgdT8bHCXJniek502GZBerFd2xWqQJ+vh
t2jhydsXc/32LHKsz75aVgA9258iRvIQB4wuQIj2viD7A0mq1Re8b1KFf/3Qcbbn+j4Tcsdkq6xs
ZrFPH/dWSnrCnVTmMjMz75nvSOhQjMO4DQSu5c6hlez2Uum3Pmg2pKKikb/X0nmuYUYCykDwuIck
aHygD3N5UVxI7WkIA6N2/+xG3gZ96rFO7FxPNFXRtSymqBPI1LOx+/gSvSZ2tnK1k3mcMtcraPg4
O8ROAQioowRIgYE8xMRKwLY5fOOXgCsT8wqPthIsqRbobpWm5O+UrvWdoz6o4Mc9kjLnyjWQkBA7
RZffaThuK1w92KCq073nglth8F0r+Y8pitBvdsbctqXqMqqtw4GjbuaYYwjvAQ6vL7TUAaEn7Mjr
gncAcIcakMi2AUBAT23q6B6PPEGq4XZ6KkKuavNT3Nz1XSdQEArGQCptxrxyWIJCZ5RGGfpnsa4h
DpQxWVhjGE0wKM/J01zZ5x6HRIl8kDxsLbah4wF+g6PXQFP4uKOOj1zyeLX1uDayS2WIAyzSbaa3
LEgNAh4GAinTifSbT5TFLukoS61oFHjiOcIuhckaskPljeSpGhqzy8LwZEL2X7A+tNwd4gWjzZAH
bClM/w3B0ChCRQotNVxWkUEeXgzh6ZY7/7vmgf8ggA5m2ZUZfAXRzDMOICQeNTxUXHuEjrRIkjnj
GO7CyOBcdRS12p1lJWfHbzMWxbGGjpXyfF72KzyV2FjKtaXGMLAQbp/2z8+E+6RyaYQ2pPT02Ssn
pYijlGq4oM3XSSbPmEsEp80TOI5EGyy4DF28UtnE68OkKePl6rlEJs3mj3QgcReMS0//NKRHhGc3
Fru0t1uNCtDOU4/YtmBBq30FveCBiRAD5nRjpe5thJGZnDzRkZuuxMFDXEKpqIjN8JbC1Hnwtq/n
MjuXqYU8JrP3xaevgmYJ33gYwmBF/NtozMM5WqXIHi7rOKB2AL824Nn9OcjUCEbrLiRv2E3NW/2K
5tQGK6FeVEW6hF65/vgz763WUwptqhEoVtGD5upbRTeZ/QcANevnBdiiwUukdfFG7OYVdA6+VQaL
ahuyGxOqniN3FS2AChxlQWzwNUyX6QXNIzUZyCXX1mYBZioEXW8RQgCKhj9kSi4O3Gctxmln2B+w
kACMnNGjuQ/XNEORZ9ZwWINYCOAQGtPSVaaVrfYRmkLQ0TyNE7UucFouEEYNXbXYKtv0V0ceiWjH
HtzDCKOwnHKIXS5u67eporDcM4Gj26wnTNhGaPdQ1/ea02x95ZhYxlHZ4jxq4bqVQWEqxUHMS0lU
QdiBnUwN4HzHJDd7mf2H3M/BfJvrz4cYvKE8zmAoXQmC+xf3M6WI4fyisV8S2BOvl7szJeMvQs50
Ad7hDukO+T9k49maE+3EOxUNp3j4eWa7GgKspRg67pgWaGkNsQ6yzh3jJtsC7ld3N3qlzgDIhC/g
yZ7yu28MXOzN3gCvfx10acfZHYAL2GT99/uPTW5nf2BygJyyYNHw64ygO2r7ndghabU+yQ4RDoGA
sDe5GERf9efEniUjTSeEkd9eEX3fg8FfjqRcKqIa4ASETj7d/dKGCqeZDaePyKL7gRB6YPgIGJ6l
dqkici/S0k55FhebjoNO70ld4NP0DT1NPluxPvyeN8+/8/qSOePEQlSalt4wT2xJ7IUSG/40v3hu
FVhQdhk8x18RIyjUtVl2UlgQGWMQJGk+RixDjulwJJ8QhDxPV/r1YEEovHpMIbOK4wZcGSW6RMow
bTkx5n4yvNX0BRGK8IWvc4IomfEHqZSp0jSpwy+vDpPbU5hF3WwoIDRvaTWridhYzmEzfHRff0ss
Q9eIH7GnAFixALtvmimpEH1GJ1KdAKGBZTpC6dBikteRXreefJaCuugtDSmPz6DeQMFIJd1hf2ur
FLWKTsP3PWm1PmPXnVCSAZgw+m/dr22XwFJAGquFoID+vAxRg1HKBmyqmtUZRv2sBGCb2PVwQHdd
lWE1Lu78B6EncoFMXYhiwAbAGkFsXpYB7jTHKO1i6irAA2fwrh4Ir5thRprSYgm3MO6toB69dsQc
GRw4FyStPz4f9U0dGTOD7ksdlBX6JPjRei8FjygB6UcCTMhw/iR67wd8Nn6dBm2XsfHpwaG7nBDB
a72ryAG0SDIuRAUGsF0wRMevEEzGenwvT8TBZe+w8/EfEQy9/y5Igy3C93P+ZCYKMKCV/D1XzWbv
uqSslgEimddGRL1rd4DTH4iLxn3JvQ7X1WnmJlkBfJtNbRSxRgNbuIWL3YgVslBPGtDpW/T/Rp2m
CChBaKP9x/Kr3qPMrtnkXIRw1mKd8Kkgi74pp0S1wAFc3Zih/ZWVpYGev24j65MCXCYr0QsknNBQ
M+55/qqfkqAGF1FMcDdRGfZh0RaqHcTNt/j2PDbqpUgNYVVIoaWUrjR/ui//0OZULc9HeCpDnMEY
woTy82PGdbpitI5IAfNAWzm4+MyfOLSB8nPwZp7qReevhLF2w/mniFQiRmF+QG2F7y7KMF07+/L7
P8QEQ+HT7f3y1WtTvVSVxfByM4R1HHC4x+96T8bJLe0WOMzyXSp4yDI/GPEJH6osn6tM0BwWM0Mk
W/+s0Oriag/9fNQEet4oyekpeOeeo2qTq9D34fRB7SAktxXs0buf9qZ2BPvUkZJaCrj3PcVGy4yO
oXaVRQSt764WWXTJR7K8nqYLN1Yxb9rrIGf0b6Og7F5aVHNB0T8iH0ZgHXdjIJ+jPbY0bu/0+t0S
yaCwma7vp8mSGMDqyXBJMcQ5ufaxTnDu/fPmuR/3MI6RkksJKxK1j9G67SrkZLGCJ2H8qSj0OwkQ
yyUOiNnjAP93K0RadaOOSYuCmjrZKfT9TGG4c6V/dXs0JY/7TaVG0R0sGC88I85xOqSsU7XI1R+r
f6ij0d/CWuZKFMy5sZHL6zN169KPr7UJOtLuixsKOB+vIEhYu/d+C27GDhiKdk72qEooLvXGcyMi
H5n2Wl/4LUMOp4GKmSk5Rl+IB/Ljer315cm/lFffJ1EIj+b//tX7xSjEl/DKHHz+HSPHP+lBMBx7
W59DZLNmIAu+R1BxybAwRyyxj0CnTvkxzNb7gLCU5S7wga23YIqv5i7llkkK4vg/CDrBLAZVtsOv
0A2mIt8mXqs/dOLiinOFG+DRLTIltQ/hbi/gwcswVoenvqll5dAwvt9tYBGBiS1XuumG4B9Cwy9b
YwrK3hyzKUBjaxgyNZDa7FP5xsG+2lknRl1b57KwPnO4niLh23866C/KfHLbZnerZD731M3Ot0mK
2XtzGrnlQmLdeiabY5+4jR1OJSu7hcNu7YBjjNMRLW1DPaAFN/FiVu7XOwuWJgsC7NCqMF+/1+ea
dKab6JFBfHPuvlcim913OD5V3Zn1zBlEysc1kngOUSNoKhcdm06ZnWDSbpHqPtIkqMPoMNTXYKPw
6m6YCnCpADxEkKXJLDaoW/p7bOsQ1oZRGGA6Ylm2sJtkzJLKkAOIP2gII131NZG4K0fGu/A8w5tc
2rZVY7JA47vx+mWDyrv3yZ8I4PhJQicayyD7GkdpEocrCscZRydnoCh2QSek1llOruQFhN4hm1Ti
cs2bTmWgmj27tpcwLZ31HD0JDJHxHBMiceaBMPM0Fma02USltyWtKlHYDwoo8NKX/8aqTeJxLI0Y
pBMjTscRWcvVCLkSPg1CPVy33kiT8MzoH4yOmvmsYD6WenZ27eV8Y+CjcR1AeJ9pPxBcDFpPtBed
aMaKmU3VN5zSq+An55b70VQxYXd8FYcCYlWfNpL/X1Ok3rdsJdBtuAzrRxqCFwSQEpTk9UD85oEo
E9DHiCXh8Y5qP8KAi2mVM4rvr/T9ix0+t4fTrM+EiSo+uZu9n2fdJeneZoBxFV9C2yph5vpVctpA
Oa3XCe4ptL2FKOriK0g6ahtGpwBXliBDOQyxlj2NnWRZ8FIvayebkoaYE5LX8hWzyemtv/G/6wR2
0cxvYk3Dr1SAZp8xKMkOhqS87pB9Dx7UVoRLMVHafXDu/jJnCspfJMVzCZcF1OqzIpx96qhPaDRc
xDCQdDG4LSEspv7h0MeKWOHBuj75+U8mbuisZ9eD0t/H8CKuadFI0taywfkokW2Qefs1odFHs9Sb
th3G82Znj71bwP6qqNcVnRkNKPGkEpr4TY5xr4OpjwGzKu2mCd7A4iBkucQChFsFn5kCB8hbsSDS
FvT0wQ0s0apVCIOarmEufI5lr8MWV60hj3y4nnlGTx82w23/knyyk5kWqdTwizH6UIQ7Ed3K48/m
uzO+ORryegfaTYqPJSXWZiHSFo9chrvaLknP21bJRX1dahkQmm2TApBmWQxSbfF7fMTGgDaqt2mr
U4U6bj0eMoVsnVKrGKlBD1H45lS+tiZBhk5R+AkrXHYfL5S5iVcvkbsW7zJKu/n0LP6jG/n1gfTB
TuiAgNe7/OGnmPhGqt/AF7JLuhfKTyG+N0a0uRNDXQdjbqJCN1DQ/YaiUoowLR6dIjEQ9g5/LdCC
7xw8+BfMAbSzs5flL9FubdBv2Uz9FY91uJmI0Yzr8OS3PJFs4v9h84GtIWZ5HtlHmO8P2S3WQcz1
RIECBMfVb0fnoZIxGyY42ubw+mC1rsAP8IDhYcKJYCeXqtk17+r5jx8zjqywikYm4WgW7KD+VbKQ
rKy2OpH/vca8YluXaTa8/8ZQ1FBxjI2V/4aEHbyvM5XRWZer85hVhmcVKP6i/vmvyr7SP6SJlhCS
a9xl8ux4PJBMKWeZkFV5zcbesfyh4YHgfQ7bBLRyaWa/rdNgOt54gtEsXTw4Ol40h4pljJpfI8Rg
Tlav7krLpzhqlqL9Iv4pGBfi95sledfBdaChmgVh3L7Uk91iKXB0yQjFs/6sGqs9dIFmGbn6dRzt
EoPiNplKZPWCTQcKZ5/GnIOmfSyguQiUh++Dx/TmfQaRAIHuX60kVWNFAhp0KTCxKwdydAPQH4gK
b2gs9cwVcZdbDe2539Yzke/ARbQH1fvAYX1hIrI2Hf/jbv/NbDG+mG/i9YF67AwZsFv03v0CwMcH
yJcZ5G6kC7vNZOaiIizEj3b3AkNv2CeJ1mo4ff6d7qP+EAvnr0+t0v2qmARQoKBsMci7KUw9zbav
oo/nTJh03f7+e1V6mA5mWG8I898xU1ukkO+wWvC9Dp+jKidXCXsYnMo1r1YXIGaJMRB3Qgc4f5Gt
XmeevOOLPZ630SQRIqvTKpW0sUBBISszIIEVLj24P2rh9umLa7kEEGVdpMIsm9dd/GXLT2MUOZNk
nEt5BBSRtaCqgsJCg140nC14uz3oXVE3STQmAqAWdaIK2APHgo7WCoM1E3kT9zk+fApXbS1o3t6D
Z6bXJOG+SDxcErfFAMJSbK1niAzni1+ngLU3sgjI0GSrg2D1kmwaVEFcYyF3Y8QwaoqkxIG4+MRU
ZdLervqAtXsltb5kLBOLG14hWMCoKNpWfn8nzk43G0dCLz4/0EI/dhM7M658YMHI6NJ/7U0+KCyR
oq6opIrSKHR3J3a/sDJXm6tTkiKVBT3S2K+jjg9SgeAuQdwd/RO1BPnEAIFPBWjjby+ULWUg9qXO
1dM3624AOTFavrMmi6keau79NlMvzimMrRt/siS+x8yDPkeu1m5V5bGmVnjpe9oLozdTQhaxiJoI
KvUvS99q38DvKVp0c5QNiwUTEw9i02pJbGK5DdCJPRscXnK+2T7CulJ3yjj7z3mxBUiBjvIGUOFD
Z46vOqEB4mKZt3GlHN44C+TZj4rD4MeCUASogFhlOV+fo0g+olUCvgFDlc3fFFi+ScMGpfkyhYZv
GxV3HhC+m1NKahs4DC1+aXpU3/fckpAYDCpoxZK4KjWiLjxHDqg+VeTj60xY9DNBtxCV/qMVBzfm
m0tYt+plTWIjeIDJwEhidbB43GM3uUPczKU9RBVOjDKXDprQikIYUPaG+SFOsQw7/NIFjPguSGZI
Sp8CVARM3a+vdF62p5/SS2e/PXC9gAZcEnT4tbcebxzC4P86+GE8rMFfAuzp39xkksGEDO/msdeF
wSNYSqdhxIs/VEZYeSDlWL/PmMzl1tyToQnGH0w0nq/TK0ZrCQF2v96M64d6LVYVcqr5YH/cOLS8
jjQmWFSoRiJiIpgEohxGhEKCOM6NNCBg7tzOY9/Iibl0gafMimlFit1sp3C1Ufi0y6K0P2CS6PEr
koJJHTvNRuVG4iRfpFsRd/muqIrCkZdZqQizYE7KZ5Eeyrg5yoxB3yvaN3QA+qhzCXlyYEftTzw5
IcAdWDyNzJnaCZ77z/mDsmehzvEu110S2xrqcUcQNGwkHbeIKMT5V7XlTJk1akibIlRLCUC+jl0a
raeog+X8ST4Yf3yfs8irGEO6V9gbJkGQDpOnT7xgjDzES7JvYV8FfGePc5sHt+MwZBH55TyHTB7E
jVvNABowlzkhc9onqDTNi1WvVVxstehV66iMTU0BP9ShsfMZzorTv9sXVQUn6TLiIVc7oqfiG98+
S7SKnV9140/OUOflEkPTfOOsRAQkjlmDpIJJasPbLW5ftNc9lRhWX0/CvaXfdTKrXHHOOE4lIoIZ
bb+pcBe0IPWF19L0cK1hLR67HGVUs6vXyrHgGwIyBFMxTnFwQzd0Bjtg9o9AC6Xc4uluf2lTQy0B
+nllTuTxeWd3bVpO9aBPk4Tu6JfjnjFcf3KAjwFPUBkrzc7BueQoTqBbedDsOcRt/ChF/nC345Mp
w3vGzdYCcJpM3U6pIZ2HlLCP1rnew1AXS8kypsqISKCi8CsQ0kBYqB8QntwGn/c3U5FKYUKOvmt3
4ujlRAettjBHmBCTWaU6Is5lbg5MHZt3AM6fx2vPMB2UjpRX/hXfP+yT+Ufp4fLtKSGCSeWtCZPO
7q5BMW2UElEfn1fnxt0myBgqw/+J1pHZu9TTuQPd3Ac7+t5XdzgQjU/PHKGeqKNXOLVJRMjTlhJU
FGRDwiF+2M7mLgqywTsAHtRba/P934aKLH62/2ZdD69yZsha79r9MKV/sZO/gc5DlnS3IoJbYQM3
zWTy9j1kjMPo2yha2ALl8xJG9E2NmaQOOXUmvIBmPGdlJHpkSX/c5LbNNzuCMH9seju+KhBTqsRU
f4Y77/F6/yBMtrMhQNAWUd/sap56iZVjt/jFcwqDsqT/cUbaZY0K6rJoznTtYi/wLj2zaKK8aGD9
NxnOc6Lr2yTemj7mIyHiXDXoZL0ECJs3mM9RozkuKBQM3crYyGRV8+5A+jsdrBGF2Q6e6oOWGbQF
kHHlgRqRw+Jmkz2vZqLMkkidnlsgAdLKD/0GqQuVrj/6kcHyjvgiEqtR/VKV10WKIqmRPpdZP03c
T7WNl6dmi/aZgo0rVjYwKaumF/7L5YJYZebSQJKXuAzdlldh1uacwUZIkSL6EvHPJh95/S121zoL
n5OdSa8NkBny9+OL3ZcQwz5sBySDqrkfLsnwz5IQnr9AFU/KD3kKlyqS3P1HnEceDN8WmX85/fA/
BjavcdjOVtHj1y7TsHYgo1e1QQ6HMZvLKzx/AIPTmslKUV9mE2O2EDADn2ibFJOeDZ+RYY6IAn+G
z0eMl1yGe/jNXVEDN8cT3Atz43MJPwpP7/dCB9kSfmdsaZkdqyeTBnonTdhFGG6PlzOcxIX9BqdA
d9i0z+fZ+55WmKIZL0aXKgh8d/lBjtAB+97hOzMa/MGEL20BMgxu/mQUV3pSu4tA7VaHY96VExvD
fv3aY09RnCE8M72aeTC3/N1MmdEzT0MEKEXjxlKVjn9+WZDBx8SHzbvRvOKf3gio76TfEVSUKe1P
haNZWbTePIADW+Yfunq9BY342E2Mq1P1V4ZGEA1noeMdvTl0rh6OyfHPZ+NFMQVTEbXzp8M73/mt
FpSrN4yMcqe53spjqIHmy2cn2bbd61aCRzcGoghXPNPeZyxe8g1xlOWHyDccjIgr233GAsDAHAy2
w54VN7MIxSq4dBWqTZ+F7ga2/L3+9aHb9zPbSC8RIqRa7EESVU0tC/FiAFAsJIYtWo7g2YbJdhb8
Zu5ZUruTTruAP548eMcQBq4kXgEI3QeANUh59TPjHsp7F70Bl2LTqOxCAae12Vn1RejkCsRow3o8
+8oQtKH8ysLH0r0FOCZ0GvPOdT1r3ANmEitPGbr4kD+b3PPJPf/au57cE6gdF8jYi8SaUd7pTfng
f2/auoI97gFRuLPlKrUAbN9g4nmrro3FzBJ8/4Dg9AGqfDcXxUu983nWNOhXczZClGukb7mkk6kj
qOwCrNjmGCt17WHgQHTFW55bBo2uwPerh1KdRvKFO6ohVg4ClT5dCgVWvLrGLNzLU2D5jA1OHyyo
FcMTrCY/4HPgzbWJSy6q4f3p+4JnaYEtH7jxRfZMF3Em3ZL1mwRH/YaC0ofKflzbWxB7UCicoAti
A9ZetQoEHfHzONmiMJSK0DnfScbz51DMjZnJ39VvEfCGaTHUcyBoGE4wHdnkgSfXbDh4hgEUjbEQ
MmwDe7sdDJMOJJyu3X7pTUxC3Qr16ziGJMohsib5Ckiqpq5KMwMNv84hL80y6ckRYBkJL8uBIem0
l8Q0Nv+kprZcn6jyOx0xnruLVB6tRlwnUltrvwXyhlltoV3VOGE2AligLvlt73WNbglVjpymrVsQ
xn8S5MRYZwXVo9HuigFFADENKZgA6DeqJvV4SgrR9PZGQOGSPKK3TKSp4j8A856VrZnaiRyxsO44
t6ZpSPkkme+RWE8Y3cVX3paCsdU7aGDW17JXhW9e9I/jXi+kIj8ABYAmYN6QSItVCtyDmtezxlCm
vHlrQaXS02JJ7YA8pWGapDvGYkZScesCMUOaueeyGjpFlum3aIdEvszO/ZiFgO74duY2vSPbBHnH
0c/WHQJPEh9aWLeYh+5QZfB62Lkw+sdqjSnuYMNs8l43/EG3+dAQ0nDnQdttx+HbRx78nuOMNiBz
JnA6l/KYF1F0NCoeDz0EEpK6dA+d4QWK74LQkESMSzz3HPHvndwXFWzygvkIDEgoCNvkPdqscSAS
va4NmfgfCw2IKpoyw7YGZDlLUKgZS1gIP5Ia80e0vwzFt2URwxaxWPX/USS3yaiv1lX1n45VDXMW
uOjhgPWHzh0C/M1Jmnhkqm4/OxXr/YnAV5Hoaa7BuCPkimQvvPN5GvgGNvmKliTpf/8nlNfIoWzv
fFiPNe6WRINQi72zknUCDzWRZVh3EwoTwnvjvdkORTE5mvITu8iy/T5nf78jo19gXM2+mB/mAG7/
O4E7I/thq9YQT1I2btjfSVsHxAtICSk2yErBJxTrT+Eh1wRFeVar4ZnBFHK+4CsrDigxqYIVl4yx
Wo1V1iGoV8eif8rvN2k0AItjTsWi4clAUThDsKmJSfsvm429i4PF8fNTv2db9MrLdOSSijMiV3F6
DWgpnN5+GDx5CfzTQjsSa14ljXtr26QUp8Tziz/MSQNbewEkouVFQ/82tWCBIGdtE3lJbmJ1/g1J
KJ5LWHujH0B86j1X25C/Yqh1Vif34kzcrEe25m2lO/rHawF7RPvk9nOgCb7A9FqvA8yR3dzuKKXy
hvK3319U46C+jhSHaw4hkQOKo0SDKfLIM7lYW9qvW3htpLk+STXYTNBPnBj+AZ0RpzYPsmx19Nda
CR1B2bUfKBFtvdsWO493xIMhF8dJhmgkOvVEcId9QJFeRmhQGfdQhfoFlss7kidu8syBewGKfMMY
GLIAF+SlCb6o2xbUhqVTzih9NlmqSJAgmQlUxj/m9RhF0sbJbwM0laMZaK02DkgLjQ2Gg9qh3IN3
ZJ6+/QhUrj+gNxeT3V+6c0BePBejI0urEL3uvrJZ+LfbYlqAeFhwd/Zqt5zGOaGQsgvjQH5+JBQz
KQFiyjV6sA8g1EblxgD/loZvRmRUXmU3mkxuWlifQHaTnEEdlPhmqz5Pyb0Gp8X67CWQ1KHJdW28
mKZpmuB3O4sgkur2Cet8yog9wJ83KfOW2APNAAbnkdIeHXROX5YuphqFtCU7WJWwv1+1sXiHPhtV
TgRmd/ASrj0VEjGXGapaJ1BVPi3h1gEq4av4oD6LU/USlSREPuluwhqohABagdiOw/vQwS8ir1iD
AH1kSkY4XBARIBKFk8buTCYICtBzO2rFrAZaLSqlLtgS/dnEbiMpH7E+PKXcO67HFIAihOzRlyov
HuQcIdO+FrHoacfrZw7HFVNLIa5gKwowXWfJ7qR4pS8TbtXuavixThd2zISf0JEkQ+PHDtjlGZHw
4e4f5uASc/JHWP7leLku1rWu4ZaXGqUUqUh0PCC9UPASDnoszc3Rxf7qGF0o4G+dMlqZSavbqlfE
utlr3HZ4WYa1ePWIyFzAWoksGpdVq9E9oAns/bvqIlKuN7+qsmyF6Te+FLHkex/3wSCdxm2krrtY
VoKwx5+deD+ZCNFDALi37TZTwjqFiQi3Eqha5g7xfNa7jd3jA/y34Wko7XJsKgt5E1N9l21V8Xbl
RtbbTV2+8XrNZeMkI1/pCnB8b4Kv1BcGme5kTQUk0BFBMBdSsh/xtcJZy9tmGLuUdHLVAAAhJ+3r
2WAbXOZnofK85m4z90+LWdxGS5CgKaKLryajn2vMp+TwjZUFI4vLcCFPjDvMEjiKNYx6dBROBGi3
CkwGIk1I+yYSdKaMLtq5DabIqiyWDrM6D5v6TRZtKd1cdhPBlcRlf6inmDG+wK7HlKdq5+S1+wm9
FJJMkdAd9z1Rn+P2FYufqCBWZPvC/NpYD4Gk2UghP9LJN0rKBLdQW8lanTNBAoHtt6pkwpUsoK4t
hpZ0m8ib6WQ78Cion24eGCBd5TqjIjx5WmFa21LfKYFsKf4cj0nhyhk5GfP6Y0D/nPdBkUgpuBHE
BJTSmnoYzUWvLw5Zl8m5rMKJes2tX8vFF+OfFu6uBfl6nn7aQ5jHy6He59H1TXpnT/DBuzBZcKA+
Zjoba/ifXe16ZKPe8i7rXITkqJLgee6jqf1eok6y9V4sdOWIKPGwgoOkXfhkdCYJ6IEHsCUp5L4x
Ub4F3CNhynE9K1WAZo05NTJ0TrM3PQqKjLU66hxqJZ7YsB9gw4aIQA3OlNX9v6S7AqmmfqpWIwZa
o/RqbGOApaqL7PYvuGYyusvuJ9yhr+JoGT8rX3VevcOLvY0b1Qf5XpxWzi2qadg2vL5h7QPZLd5E
XhJV+LTWJN212LJIuBky8pWD4dT4IUdOrasRw8bcy4eYeY+cVIc/+Bf0El+FsTPKagQjLPH+QG/v
9uiuf+MEGZlrB/cdi6Yi8WKKnRXH8R3meo2TjMMtUdHr1b5XMPgI4FdFpr+yGH1Fn96u1HtvMTDB
5nh6cQtjGWIfvhXMeWPjQHOZbFqZ7fqqv+Q+JGc73J4VPbPtJ3J86a6+8LOoC3sCBI+FPewSnqsB
ouzgVpomhUUY4CfNRokTgqIj9euHkcQzqw6KQ9MwZhetdlnkkrTQVkHJMcB0KRQPE3V1/VzxVvSB
X5Rag1wmsbu+hTGsMfET+Y97J8cmfmeOWcL+TnHipn/ffsxXvaNVWXbtZrwEeeGOPEJncPq7MYOJ
6UKsC0hGfcwGI4uoDXl/PQkxJn70ObOZXrDz7wuzTGhlfhlNa7bV3Jywt7HBbaquEtcsYZQ7Qc34
tbuhVc5MFKk9C/1tojfDlqYiImrazm+y0DtjvaRrxIZ1LIbvoUzUehEvdUY/5vyisQ7BwBlWa0PV
KeWxhgH77t3YzqHIhqoIlXOasR21FUd/kiVD1ua4pP67kWjpenGGfbq1+R6AQR3geywYkWt5mlQg
dDLx7/4lxePQEzq2XkVYd3BLK3wdhj/+zbIwtAQPhDtjYFeqXwF+sOP+t1hCZmKvrUV1tg42F7h9
rhlRspyOCZQWkAGb7o5eEOCplyhfqlcn3BzAfdYMKwSt9tYX47rCPeE3n+SYR7bboCkwset39IMv
Gd37DegaPFVTFXsmqoCr9cDXBa76EYTL0ohisC6nN3ehoavlSeED2OR7GkBX/Ugd2U1IY4c5UcmP
wYi8F7eWbxu4TkynLK9DtjiX/MlJs/CHY2SL8V9pTpbgVAZy/4cqunQBq5HQJPby+sdfjqlPDopi
UI99pLp9+FCGE8JPsrG65Qe+3AlV7RfEVTPtw9MDPO25BGun8foVzStiw+AFsZLbSjsg7dnw8E0a
SuxxDmgJ/HWcuU2s1uN0pl9sQ6x40nYAozuYKS0K903JUAqyhoywlgL8Ui3vrpK5r/XQXobAKIXs
wHfkygyrJhnMWmcByVGpIa3djBrqYn740ZuzXnwWdCTb19iIUIAzQ6ijHP4lTw4mX0u4ihDIHYD8
WVeFWdZyTy/cBnukDSOv+e6ubvivmDZ9VY9OZoDZJS0B0KDACVx4Kqe6q2NIyeLs7/36/1y5Agdc
Au/o/sFnMw3v+2YpGLRifECpFZYbY5Hbvau9yuLbSN1ohXSHfViTkLcyEFtOGtyjzCjR9b/vxizc
uHGeKvH3R4192YYM0fo0Nru24TcUjDR3oPj3f2FZogxsEAxxwRkYhHgANCtB/AdDNaoZuIBXDeXi
0Q64f8LjmYSQkm+pQKnbbp3Rx1VpD3Yd/8Y9xZKYuTMVNqX77pMHyGeNQTtIEc6z0zc/5qdGSrjU
NK6/54njJgkwba/lJOQOtuULulpiQLZYVBn11W9O8FDVrhEAVjf1vcm43IRecrm5He6hTbP5TVa9
NZyayvN5ilioSavLmG5XdtzdKBWhfhXDj+WHdtAkTIN7j8vCaDUFp4nMudVI8v3sTP3XkesoMfoY
rwpdSZC1/uje4IfPUqDEE0ovsshrt27eX/VODxaeVbiMdPviNOdYdEAm+/ZYARSUmERWxCwQnUuP
Q0ygBR2rZbDCiHZImXgIEuRSYHh8KRVKupQYWatFLSsH+REgxWuDaMDUKBhNw0tiltgiDTCppxfb
+Zw1OauqmK528KM1LmZfPxP1OR76pkkcj2V1H/Vp9/pxG7WHnTIKRgnH5ksoNyZBNAaXWg7OKmLs
B66xiRnS4uf7jJ/bqgqLgz6MLkxBK4e0WLC1h/XWSCbXxIE0Utj35AKtZPo/XjU2u0E3Dv1wf0gy
Jddpsug/nX7edbtx0rpzt2Piz+9AMFOK+QSaCYUEQZEUYqCO+d2LgjE27ChfRqn+yTzVmEELl4Fw
9Q/qGKIGxl3N4fy6Z2wLL1WBNR6ODpODNmKv0/ytNCpm8DvM+DrdraE+MIu4PE1AQjsX1yYQTBTB
U41Kik5ocdnO4lUwSv5wH4/r+8iICYS41dH2horgMM3gkX+8JjIJCT5owg1QdemcDg99eMQnBfh+
25YL98OWJnW7WHCB/u55vG6wbWRuKJ208WCB/NgDZbfyfPef9g4C7wELTN7WpwjIl0Ln0/h+s829
CkEZ1AFdLjFQH7ZFXPgw9uEoE/QcDHI/ztoJbGH9O3vj8eVHUIcP+mxnEf71NyD0m7XRMgJgLRR4
zWvxxsC+ogjxoYCXszqcZqXjbqwpbbJD25gW0smT481E+RZfuC6omkjfu528qlmBbmdFXINX6DNr
0WfY16nRpQ0v9TP4kBTGTg7td+rNd7X1h/Q7kzx1DeUlgn+m6+q2N6ky1PEdHK5c126ZMHB5o7iu
jWkYurmyKRs1Bj6XPpvkgFPOR4MDYHcSckA5vSvNqBTfDOIpmS5HdlRUA4HVvn2qQReQCKHURrct
4+R1HyGntCfgerQshAwQ9rkucpsXwU7SkC9yCYumNbzEdqNE6Oj20c7m4fVUGwf4AGiWsM35dfgt
a2+yWHkjKL7qdRP8GORFD6Dl+jXZMCZcVXQ+Xjn4YUO3zoEwqnehhm0b/a1WaDH3svETS98xPjJC
WrwT2TSNTvCw739bV+ShBTs04QCHMYQPzAgFvV3JouqcPGHwin4ZsfQIXvqRK7mdoZADvLNwzf9t
eRwXRkf31l0cAIibSTm/DuLdQgzx/edKVjcTyB+LomoHFyd8U+vyEGkDhMPJENgbDMbrhxsKeI15
FWzv9154ipXde+8IpYJkV8cglyGZWDTtlHaYRF7TLIzkRK1SEUX0sAMX8HA85NZo9yEKIy7Zk+9Y
/VdAtnP6YmxGaqq/bJe5/HbSUrVZKu+hccs5gUhom4WixuYZdoat44pwb9K6mPT7aJH8M3KlgdLN
5N3dGq+Y2QhHdcoVUF2T96r3uM3RypQfmmNZS9N321c6bz3jJzm3FGv4gCNpyVCx5fyWMULcp2nn
uEwxfaJHdjYkFJjt2ndOA1ah2ueq/HdFrpy4oiSgQv/3LI7XCx/HjDRx3+jG3nHw1cehO7lBTYUI
0TwQStPt8KIm7b42TKylEVsR0OW+34e+oDfaxiP6R2MQL+f1drms0gbMGQXu0QCXqPWiMBugKmxH
DUajwCDXuc/FSeXeg9ubJQwZ/twtoH2Q7mMfblFfKEpRgA8F8AGzTX64ahTiy5uRQxzlCJLu7KPl
WQAoQxkQOkOvgTg7GN4+kH6RmC4kqrC3BxZULUfPm92cbZpC3drYoQkG0vEPeUWBrMtvAHGU/Lu3
dN51zujUmgR0IBN06k97v2ye6JCl5FkO6pmuVRF+FMtVPwiOYdLSLxCN+Sm5+nagKW+AarUKQLSC
0f8uck57QHZhRFt84j7D5VG0XxgQ4QcqHdAi1ZaUjc/QGMw4y+P2MzQuyMBpTbgqlG7RBim8fPJU
LMVFwdjahyGA8JZsCxNY7azEfmEo9AJ7UsU+b9sVOlGtyQpMXUgPuUJ85r4kBrS9ZYw1YrDmAxXy
ucPSCKlGrAXXxfPEcSvifApxIEBxJbonQWs2S9nyLR+UZ2qUHHdI3yzZlXwWxN25ChidaQtzCrJc
0K1syyWIfGPvjC5dRkSALrKBPslWhd02WqvYQBBALP2AoIVcHlnhQKiFIw3/dHJgn7a5XntuxQWh
tz+IFi9hEIZL9d2XI1qb8lTvW3cSwxro8GN1iUeqqxskmaMI/QfLTvoRgUw1E2MIY3OX8jlS4OVD
v8UMNduFgrdRMUqCt1rOYJOJ08xnK09ZOpCMmjmrGiiLTxo+gO6nSjHfp3SV4Qtm9PAjc8lV5Sx6
pYRub4YQkA56wNJkQjfLh14rxAhkAJhKO9VR+/RVg0G1q1Q/rs9Kcia+Vt9w25BSzMYcN6S64FId
X/zWlV61vrQj68+1rlmvgouLgXK1QwWTUYNGByzxwbbT/KKtMiSHb9plFOeQKfKPA6Du/HkMTX3r
4Gp2iuuUO6Ti0XP5ldzXmx4T5zJn12tuevNZDavVvIUo0zV/+V6nHeKsbzPHC2pktsXfr7irKsjZ
ZWHXhvz74gyQtdETAa7LYr7YGgtVsh7xLLKEmUi99jeuPA7xC3dXPcTxxmLQG+IvMFYtzVvuOrig
D+Ui1620MIJgZOlHGQ4XYU2OpJqnIdQ1UdkoX89KHxBoZ3tX6T4dDYoAKMfl3dh3JAhRusik5+n+
qEq9KePB83CbWmnYRsyzOl/wXsgySEyuFK6pviJCgLKYd1dw6toSCg2HdAaNjEMQAbszezbLbE+1
Hf5CefVAkWhO8T7um49NeKetdDKPxhA76Ef315faY6wnISEU+ertvJ2uUzB4B+2FZxIEDalK3D6z
lQZHgb3fqjbT5XVXeweGZLltYQ/Jp+jQHnVO3grmA/cnKal9lG9eyJNUSnVvn5sH76daa15mSvUV
bH549PULlhSj2+0OdCRZrPDJqjkxRBoURY5N5UPnWRtlBY0Eg3wzLC1H/12RVQFcDeiFVJmFu8eX
aXmkeeH3CDZhk1eOgLtLA/Uo3QOrcWXh8jFBJKloGQw64Z8q14FPmS4jFAQ8YGCRU5977xSlafOm
yAU6oaImjOUO4ooYyyKgOH0ETf3QMtAXX7zVsXahStEjMPzACLWTqcAltf0vcjUiTKDw0mBC9xey
Vo0l2N5M2G17MAeKSir/B+cgPuiZh4G9cxbiVSA40UcyHNZ2Mn5rdb8y3KTZzduBY6Wc60lppJf4
HwVffp4y9n/Eh25ummh+Da85aKX4apvWOOTeLNGbAvi+Cn2oNJ4av8f04pgOkbOmXrMKhvJyMzNS
NBxhghHvSOoS3HZouVaLft36rNe/cUZftscsw5eI4k3ZYUDSWFwtk3PAiSy/rd4hJihJxXXR7yud
9mUyBAtHwKbUfxrE5Me99tX4nME0PZ1gIWrEt05PX/ng0rM7fjYiEk3JOE2YuhJBJTlYxDFhqG/O
n8qxhUwbw+zdQxAw7qgfhrKrnbY/A6MtXPraxoLI5ecJ/dTLCOsnH1+W3Z/IDnlrEPkvDcDtodGw
5sXpd+turL5aWDqpQRb6Gcp+5imc95LoX3Mu3Sn01GiZlO8+4faBe+1Z7TL1q8A3UKSt/dMPIR+E
mtxJl9PhLZqpjIjd6E95jsAIy/l0kbSQnXNB4Jfak+GUeV1Reb3bze+zEHZevqbi1i5S+EAE6Ixe
+m9qoVo7VYoNn3MqS7luajp/8guxoQuCkRuhpLvSpwz7Oh2rqgEZ35wdQgxwvdcmfxjIpVJsY5L5
kC7eMPHGDsckZLK8WsjEHiGiAwRhVSlhomJQR+7ED/I8Wu8/WlOkdK4eX4wWxL22maBDTuYq4lR2
kr2aX+X2+dcBmUqq9prI3hvsIDReDUOY+ZEc5Jc8bh9p/gqyZX6SW5tWFU/1mKTfo0uYAQ3AlPvl
hfjb0tLRLhXcBCoji6nz9o5agRgRrA8HXiiHA8+9G+PJHiQVMqgzD6XxjczEtwQO7qCvTg4KCUU0
VNitVxZYSa6xRSBLI89blC47Wm4Ox1F+l35FAlT5kH4KEXkv1aKOvVcZyqG2bbwBnatsE2yH+Lq5
IHHUQswbfyZb9NgiK3wBx0AFc1TrivLTjUV7J5mxcKnnQbHLUkU9e8MbkhKX1kvMGQnDQpiwn/2Y
UP9Ek9sEND3CMlvGOaYNaxmpNAvir2yzS8yIrSz/Wp5T++YtyxMmEpmRsiAfsvRcjvxgvvSgbfh9
MZ4hPOtsqyiTRqNiHN3B/YvuDJFP3RQao0S6XBvz+i2B428MV094JebnkQt7TxRY2g33c3fooiCg
nshqZkTh68Whe/WL5CTHd3Kcuy8JDFwH4+OQkQnipz15Xz99j6b9fYcIgS99CMp9Hk5f5QkmbRY3
HB8dSUCw4cQIQB514I/s88wnvvBB4QSjlJf9JkRMSdGGXyKb4uaUUQkGDctCplj/O3KSyw3D5hb8
mWpah8MfnyjspezL5uxzjnN+IQvaApesDFzLtf76Cmg/gxxMu0SJ2eOIjCYa0R/Kpg7XJh8VhWQ3
Fs4sJugn7E7FABnQqKJbph2R+SKbQ7ZwR9L40MvQ2jtFzC4X2FAG8x94ICwge30P8Kj6AIuAhsz9
X2iYyJufHfbhEzK5Z8nLt4bLIioT6TpR4LzHkHR7xfmY+pWAMmN5fWfGSt2pT24XHr9S/kcgyH6M
mo12QGtAMRhnc7sapzMrg7lVIqtwh2R3Zc/CpOJq7tT7CczN4xp1jmeu4JxD4zOwCiOY8epMBaga
iW2kSmi+5t1IdjpZ9SA6g5JQ6dnnBN4u+32FXttEe4fO2+5k7K+wVBNHC1dm35qo8dl4tsiQjAET
A4mJKjJyrwEhMEl4STqi3ttYU4HtaYPo7HO79BhJWhMyDku8sevM6/hzrWUcDxDRc9OgpWlCN/M2
3T23CUDEOlYKtWYM2dJFJiL7/K3lzyuz+RoYXGDheJvGcE4/I7ni3rWCyKvXHKg2UAVwcDeHE0aF
W+2GBOimE0HmJ4PA5Hg9r8Sc28ssXLhw+Qve9BK2IIFwAoOcNZP3CpjoaQj2p7BMaJYoBX6xg0Vn
bBV8AHMwshS1AqzZEIF5PrL4v/oov6b+2vytRMlB6WJVSSJPvwUvFLT/M1bTuRi7aHEsdXVG3SSp
SIC1g7NOEO9WPS8TmAHaH/rxVrrFLt79mznuCCqURuTXM+mk2ITHkKXLw1g5Ui1fy17h9y5Fbh61
zkvgT2P1xfpYhQlGIQyC1jCGojPouIl5Fsr4tm1YC3haesPO5eD2TNn7hRprTv1gSuPXQXm6hvzH
RTWXlkIaATYIqS0JlR0T0hQhJC1JfFDwegC7RBizgLTEYy4wod/izrcyK8n1bdEvT3qwOenr7uU2
2DLep0sOGUsDG2kyMqrBZ4Jjkyd2p/0U4XRApXUWCDzI747vC9zFRR5FkIUCJcRqGeBCWtKArCqG
9+OvIDhAIXu97kXy7sC3RKMpBTcuLRXn/SNpJIKbDkBJNx8nQtQMXsDInWGsQuX1ZtbNU8BREtqu
YS/sfOGN6nd/xCQU5A/uyy+tuukGbCvCQx4v8DIw17gqusrbRSPey10rgY/HCnSwAK7s4oHzSfbW
0K/UNePcpYf7SS+vcxlQPyf1+8s5KLJVtazlNMji4MWEiwAT73hU4H/I1lS1WjBECTExIWmyUKW6
5AMiwFOfVdywsizltZawDq7C2Mu1oeouKPVdycAjeend0ko1dTHA3S65eALFDNzljA7aTrpTdJx/
V2BubEiqPlDQ3qhdM9L5MALNb/Gqvq7Jr3Y1A7bg5Sq3AXPhh11iidrCullYj/3sxTjPptDc9+FU
aLkQhj359E1IO05tdqOuTo4zc336BTKDht08vkUGdnfL3MkWVZcRE1s+BtuPoj1/QXEUaNjAyiuC
qYW++U/ut/IgKEXSy7aXLjs0PQvNEGRXPg2WuEldLJMge2fJT4l1l0LGRWAY3SuooMivU801g+uS
+t1qwj0+sN2y3wQ55VX5YlhLlz37A1g1eDIctner+PknLIHtAaBM4Zc/TAInkfU5GMfDH9vg1F5a
n59Z4Y3SdrTN192MWWT8Tg3J0uV8IXGIdmX+XvA5IvBBiatcDqpb6CbhhogFcJB8hUGitKvrSwYk
3EwtT3IfKIjYuVYw0sPG7OHuEDVa+q5EdBsMo6Ou39+T4oRLeq4sL8pHx/8Ks5ARAXH2b+qi0RCF
zhDsEk3x2o4NCjuSL76HKb7yMM1vUoEGaTj6akZf8pWrDm2ApLY3jfgY0wkSK6+jyJvkFh71EmM8
5jFH2PCe116RJLvzZEu6kCm4mXfVZZJWdd5h8WWAYwHkG/7XOZfwHj9fB+C3BveC+qUQau43VxUW
XVgPi+3XxB7Q2NM9z+a2dKaFnxewlxI4JUFl8kQN6HOranIPsv2m/Qb4ogGgeFntTvwJi2uBbOcT
+CM9ZQcsBm/PFNhmY1HItw2LS4vzgKdkETBPmKkTZ2kSvnERJuKGcZ3F6F72YTv3OIU0YfVnekLF
OsbgwkQiwHCENcrji5FzPs/Zst5KnDNMPMUfupSky/hhUR02iagrH40lS9gyRD2jAac0sEW7s0k6
L2lVByMDWyIMH3+tVB17W1hps7mRaLR3ZHBmlkTSI+JiVExFFEC/CTeoC0hoM26f9IiCW4XuVrLK
1zQGMKF/w0k/AB1r5U3Kb7Dk5dZaf4LDD0GgUgXcXr2AMrUx8o+OrVlwSqcn+rkmR+oVeVbRGLcr
HfryYC7JtHI4bSFlMqIju5jcGap7Pozkl/rTWBrNO1a+K8xCoWXJn200VhHKwI17cGUla9kiliAK
t3z43Z8Ds9N6APpHk1s0TRfNJd248VPF1Hc/6hYBFjwFbSOuFuhlOWaZz2qhxADgAY3Kg6j471px
e28iomeQX8teuacOO3GzTiii5vvP4CgvEFLO/+vU8ph7igGgSP6catuado+iE40g1RUN2OyK3dlz
IJtp/tN349LfMeqdWDOB4UFVlLGVE9FvwxQD6/AArvCFIhkc4dgFpfa7BGZmOFeQcGxrpc8NK2qC
31dP9eze1PAoo10uhZ+rqDv8KwnYgKn/m8poWxSbwxoiFYYkRJ5FZ+7m+jW2KG6pAco8iLy6R3BE
T0K6z069yXJ1E/Mql6JnFsrPhVKpKsRe9g7jc8DNj9p3PyO1oHFSVH41U8KbI3Sb8TlzX/GtaMx+
BE77SpKkh8fc2K/74qBevq/Mt5ye29r9dAPb9m0OpzTSDTXcVsyeHOblK9ueatA1w45bFTgXRRLu
rDFafSNCRbA1ajgjwatyaGi2UfPn6EDxipFNZkJy1TkvUDZMs16r/UVWTcY++KL6a1P/ctrGKYD/
s9kYypGGMq+S8xEKvS8CVk32ZE4bQwstVewGRxZaTqnyTC4BqV7V1TWjebLkdTAiwzKx7ql4xl6J
/ldf4Qj8Yaj2vP046xjWstgrVyQap3tWTxyk+qjLG9dlTCSEjqUV6EMbZ2bm+NuioSLvc2OGG6N7
PXK/3/iLClAYMksctL0lSmS5cbXhE/rWvF+jN1a52MOT/qTvobob0WDA6cI12Nlzmm0Z9h/b3G2z
bUucUPlGtDGwYuaNZUoZKaFypTto64yF4Eeu7STSuy2mZVxZvXr7WZ8bEzmculr4oA/FFvZaWIWF
l3LsJZH9OAQn2ftzaoB9LBO8teuwRqHJew1LWrzgKLYkq1Spwb831sLW2yhGEXFU8mP5sCuEZDaS
5A5Q2mrSV6uXbH9fPU/WgkbxWXy4HSK2361eIsKoDUMhijAmsQsydsfJemioj0HRnrsRxWHyItIv
XqSC5GIhJVTyl2Tre3+TJP1zslnr550hue66p74u9tYTE0M/XahWx/4VbPBD8F2PbNc8CdIDuQ+6
tYhdZHOdSRIZ099V/i7tSUCFPtTywvTw6/GyBNc0Avly8P1+skM7lQ1UAimyG3Xhq/8St4orJkq/
vR5u35D/A4t8jyeCRUOHHwCEeZNvyUVT1jSjpMoCKKH7yfbrVw0FRqpBFyt/oadL21UkDloYGC7D
OFDyWZf7PjG1L+MBwbWWkxMF/ocys9jza7T9j1j53ZhmAvYZWWE52bxoGb1LbyNf2g9+4To9zPEi
lm5vihWRIrPlvEVN7X37saN9FIds4UYxpaekV9rMbYBIcU17tAr1AwFyMn+IgZRu7TqGg+0JYbc6
fldh+gy4epLhzEyBTNJgg3SJGcNa/VGb2hNIxFacYCrmAN7TaGymYwZsahcxgZo/6ODjRqJCp9bL
4wR4APLJjx/PImZvpvad2o4LeXu94LHiGfKRtobOqXJ63B08bRY5yVSTiMnCXUUQoFdXrrtn5Z54
MCSIjjdmr6jfF2R/HBlF9MU3lFvYNKjKursjTqPYyV/M+l/YB4tAWXA+P653s0p7gigzpFUiROxj
BsPJeTHh0kF3vZH4RL8owqqKQIoPuiHno5oL0tdUVNUovlKMEVNTDnpy3Ep4N4evA9/Xx7Ch+peu
cSVBYGhKIjg25ULIEhv2ou5/R4+gl9UaAe/1/dr/TnUbo485Dlepr0ofxAf98ZRROBK4vDVQJBB5
RXV+/LwvBJiHgNWxBtvcO2OHMW0Ypgyqgcvo+Nfx6PSiaAVtnjkhAVZP5bJ4sAu4Ha4B/5cIZZTP
sWz/Q2aCYIoeeX39/ZRrpXTsWN5OnPZqWQuS8RmaTlxXDAkSVxdCv9T1VM0wHPafCRlbrU81uft/
E3IDcit8n/6Kkl35GUfufJFaSOVPahKBvAvVVeAuJVo7Kbf4jpy6/wRVpCKt3o7HYS/LztgNtInJ
Pdr356yCMhOUVd8XJpwLgMuCkVdslQenXcZxAeDFHOVMxGzhJQrKLTG6XyPXZyS9fR2ugZXMwr9M
AzwDahzj1VehyqiSvuf+lEgm7bdF6/9YonFZ6gxTtZXIwNKOdl/LctPcZbnHlkMP0mAuoxrLQyzG
DILhlVICI52sMH+r5S4lsTqhalva7rrZXE+PVFkM6mTAEETGHnGQl5xBWMTMJlRd7dzIfvHLINB/
pMgNmn6YKpoNb5QSG8HOjvkDTgfVap0JH+KexxLwjZstGv5JNTpQg44qKakMXbF1yrN9xsI5Q9fz
Y7aD4nNCNfnG903PpnFeMh5QP33anaX9/ME/jhG5rDsm3mNB6UbNOQ6dh4JFlkFwtU2cExE3AAe0
9AV5Vanw9ah5V6Fu6R/4ZHo4YVzWgMOeGTWfamhOAvXin1bW4+auSPxvVg2vF2f+iUTR0wt821/M
MX92mRbn9dqAzWyQVzZGjvf4ppAJV8zMwYYBrM4lHZsNVuN1bDgExs5QpqhBPM8QktpDh0/FifjO
0h2rzVk64cnbFarZMS31FY1ZHG0WeMeudyabAeSkcqRl3xy9MjT4gEU5MIuKWJjCNeZq7KyshcA6
s6xvPDRUdSDCfMKDfdzlfNi5UUHd25J7hXyLQ2faMPT8rXLzDsWwUpQauWEkQV1xr9b+c2Qutwpu
fC3Kh11o7Q2LhQRqrIzONRIRBbY7qCUq9LasQ/ycjBFgTKQL3v7a+6PhkSgrY6zl+ErD3+V+OMAv
uY/DbsvE+tPgNSlUwlIzvNi9eqpxuJ1Cawu1nF/cvU6Or+wAbjOjqUdOltzLM5J/izY9e9xIK3wD
6QbwhqtUyEN6q0ZYjE11f/3JCX1X4ov7AKlSNeQq1t/urgKdwRX+0ssHu5WSWKkZloQuwXPkpLv1
JmhxCPmTWpRkA6/YLGiESoAuXys5Z1u/CRTv/qazswDH09bOYUuk8h0CRaEbAg+nkTr8Oyb+5UA9
rbstX3JIEnnYNhACqyUN0ZfeHfCLe2+s9r9F0RvJonJdFyKEceZwlrK2WloBevoSBg5XUnW3/mgU
DxFGVUSl09/CAd4vxy5Xpq22ukaoKI3vt5JXzntoRCbTjKlETBBeqKHsXzV/Zzf7x0tVVqD6Q6nT
bx2YpWcLCJV6mkQVS9YKx9Lmr48wrICNmEiEPCOMDTFYto0jy0sEeVvKMecLWlzvlNX2IDpH9l++
ge5GaRHJcv4AR7+f/S7LzOwaOkQBndmbQrHTZ/LCAjqXlFFUtjuYt0yt1SfuBgaReJk8I+8iFjP+
HdTKAtrmsXrssN/zh599uBAIm5F/xzCO4l4WyHm5BZ9cRKqUmClM4Mn2HVu63QxK9TNIaKSIhOuv
zHo6l1lKBe1WhFKKfKNezkIXQAuCCz9hN/LwOesgGaVULJVszZm8k3BEeL/lYCG3+uD57YtR02XO
aaitgFj7oqefIqq0FR0wWKe8pOJXMYZXbqKjQ16idhnmCYiHnFnhqrrp0jDZB5hzYXg+gYLDIlXn
Cd2qkkAujDmHWOtLUJhI4g1sirbnkn/AoMurzcm2fCCr0tyMoJW9WeTFF2Q5lc7jU6tL2T+zU+DA
YGwtidly68ZHSEhiePM5ohv4DZfkmuiEtW4H8sSswHRvnC9+krRnMjvtBFTwPuidEL4gu5VIX8IB
Mb/TlWLaY/eIShgnLQQi1LoLLqUAzxitz1j4lur4mGOe3IkDVSz5+0yAm/M3wDTPf544Y22uqsev
3dAdzE5xGjrN1NDNOYLODqSR7eYPS4Zh9aDF2/EcyOFXd02XfSZE1N6dNm5ce/aZ3Wu+aVAtwSGT
qLRRpO4ItilLo6cB5N7vtjhgGQqPnWFhVjkUALIfssxmCK/B605+93lxwXNwGyZJZwpkSEdCtrYr
g9LMMh6p9QaIH0vaxCQbwj1NTMOBPmKHndejEyc+dmTNJVLg6zBKhbzJ+1EKCczPF0IN59CrVck3
Frxp1hkhTMTi9mMoxRhGku1o2vWuO+AjpLFVArJc1DigKqOwvA+DON6iNIhex+zG5DYVxW4GXzHV
LJbR/gy2aMZHzumhAoYtFkDOP/0QzSHJ6M4mZfZ3DkgJZEC5cvvVRRVvgIvOtqaCZlmuKJmwsGGc
AakMr0FiiyXlU5JcFFtDM0EllQ+YSvF7FHpt/isp6RKmeuyjCUMABvLNVlBl8MN7vAbcCul7Tmy8
6vAmllleAsEI6gbRaINrMdxdrTagXkbPCnhS8dyUaTpJ4x07k/7IooGQ1jnj/Nxhg9ei1kDbDeCr
SRUDPTNePdWXVs+zOZ3HTQuaGPrTGc3yBFodvs3cxAwolVrU/YdzZB3L5I7b9cWNMeUpfqkWzXqm
/l7G0/Ezf+icsfzsFEAqvxcXvIZsJMnDirLWdQJDYIzDR1kLOEoRGy7lRX/xPW6nxkNGJoRBJ7Id
C0BUA8TDg++UhdQ1p7bNM0JBgHUmH1Oe6Q+r7piWG6DJZm4Dhj6Vi8dZ7vpkXbin0tkhafawNBQT
wBCsRcOJAT/HCBOJUICEcag0UcrnH68lR/rwUlPdAqb781f5fHTbsq/uWslI27N9Y/ArHl63vvaE
6OGqnMH++oyMMOFLc3BAJB+gxJD6tYsROMPiFi3016a4Z3eIKgf8B4w0zrZ1Uaizd7MBFf/HMZ0D
vL4a6wmss0xkqYtMZHerviEUw9jPjSm2LR8Rgum/hV9yCsXFBaiSqnV47gzFv1GfGcRPu355Uoff
8x4jVhxENsVN4Rk/iRx5Xt+dLPD7m2SiKcfqSr/39XUktKeU2lBw8FEpcAOVbAZEgbL71okTNo4o
eTBujfR77FjmsVR8dLiGMkq3hfaWQ9znT/aPruEsQoh5EyZoIVq4LMY2tUFlk0VC+rGE9rlE8HLp
f1wNWPn0jfzSsjHNzb6qqBpA/svroEHzJcaZAXdfIzztoMj8j+wkkFweL4AVy0mihaVlJve+gvwm
7JvnTEsvpLEmAljuFWS31sQpFnnAkHkH8xkJM+6YBZNDldW1qP8WwdD5ihYqyApbTRG6i2zRwtRX
PBiD6mMUOlLcTtGGPVCRcXUtKWXJnawlmtRCTfNJq8DAOuET8LYxLhcRNkjwR19cRmYF+xSU9JLP
6R7m1KvhY1xawUgzfHXNa+w+Gc/a/m8+f5xZqJJkkX2wQMHovFhUHZvcbOMOVJQyRaUpa0O7r7Gh
eVunrVCdMlrzz3q23/oKC9L2rW9jH8xIvByvIbDGpeXuxVy5DDDhDDNaf7VR9Ihq709HwuLzj9uW
gn3oqvwIZyCsldoafsv5g0y6dZM6//+X/Fu84GhKixftkRYZXwFeSmAfmFxIIJtcbhyS6O4cnHLD
n0hHtFPLErIkmNGpZ+Q2A7TAeKjZ5HEir8wANkyIbha6KbgiiB2odNV9VPwAkmckeCMa3ctappuc
/jt3Vzs2Imp3lxZ+ZWezy1sM9/M2hzDOg4gzxiKY501wAYu+VkMb2fAADjZ24+MsBut5hHrhFRZV
ruQiEshYuGekLEDlh0wlJs5gB3V/w6qS80nrDUgGSCfHEr4oG518IxbZAu5kPhuemnjn+mFg7ZvI
rD5/EbCRi9ci4nUvDm1nKNKsrODXnA52CKMkyvzPK5jGm4LfM2YVebcM4M5lkqMzV5gWri4VTM4k
/HAbZO9jmBqvc4QN6R7yKY3zhUROpVb18t8iVSEiKBeKX+j7Xx2FH3jz1F5fTVYQCbd0PehBK+V0
5iacGiOCUlBvdPrTEgIED9bMwDmtOfKplZpjAsVSZTaCbueNH89XmDaUex0x6id5hRcr7T0Ioy3e
U99QDihDWpnKlIsVvV9u0VEIS2ibK6TPvBncAvLIk4T9vPow63ak9fhkz60ULbh8dfVOPUdyRmF9
jqP9JUmvAz7elSuwRY2MR/GhJ4XqIrRiC2Q7ej8+lPzClM5zAr7x07r1u3yQDfmAJi7K7kvgiwOS
mJzAHFeMrYPh9VEn6Y2uHtyPSE/WwwoLh2PY+yAuQOM3+RXaLgXLK3kY+CvA8KX4FdYeYJ/j3qv9
Q81JTDvE8xQuz/wWbQE6u5JHeO4ABIM4nLeDq2LiwMb/KB4+oZAYZ29jyyTZkbJSAMtqqXt81Rqi
igwkKdRnOSzuDaYrf8zwvKz1+knkA4y9LH2tjlhDTB5K+kpjyeVEtB6+hfw3WUU27+Eq6eZbnTa1
qcr6Tq5T4Y+TPKY+0J0cv6NWUV9E5gC2ujMinEWmkt0HX5Qxsp7+igH864Gasx5np7O9RWgfv/fJ
/3q6T4oMsUmusjZ6O68afPr/Cax13UJAjKC7XBUyG7K8kzu53GeE9HH/CD5rRHMumuxE0nnbuwF1
Bmu85eWmJ3eQOfSCXA6N1ahgENrvJilqGD7u0tJScUdy8K6VGdswam4AnR3ugWeBlpmLHWnU+dhF
HI4IUVdWBXZaQ2sg6i7Ho/P+VMIYeND743hYrHc12UkL+/s+B93fB/FZRJNlqp7lyF7O/zHeqrRq
R1P9KUSU2JQGNRbZUAxmpxE2gPrrbOwKQEQKXyocD4JqcVVPvPItsqQjJtU0IkoOJZIZtZkT6BR8
g2r523YBQ9dVfXJxc4RBE2RmhXOqc+tETYccA+8GWQQXEl/6eyA1XXLWSKa6NrsCu1rmh3nTcZiR
UeKaNu5TOvpUvGirZzSHkB0gNxVHav4PjddvA5/TQH8096Kuljr3/eZvqnlfqc3aey78krNhINU/
x06VkA5CLIcl+Iu1sMaIh8/lmwjzmkeUoX09RfLERz0zPADkUPAFieKFnfFM3p0RnF6EnfJ4Mdo5
SodLHaMHU6uWdgyv0OEo4CyU3lWN6Aav799DHdeVPIOXbm/UJ0608pgCl8HLHLTUMRLX1ArR6Jq9
rQKjK1K5GwtE+xMT1ZABqNa8EKvgEFaVfnOKvV8BoJ5mhbSGZDi9wcwvvxx+xwXvQqQgnEgzZYfS
3xkTNQcXAzZsnY8KyvIlbH0fqZdTEreYmZto+IqSJM5gCfhfI+xEKehWAGjK+UckMMIG8lp5es5H
jQQf3CitnRLXuDRtl0PmmOXvqOcPh7nv5jZasJnFkJrgtfKHtgpA8W4XmTNckKF9JhzdlaV2TUgo
rOr5zMEE3fcb8ZTJOTdKG5tBd6IvrBbzHkvWXuZO8HLfUwzwCQe2bmWOapnkSq4HF8ieIWfr+uk2
LGLbxbu1PCawPytSjvT5wt5kskCHrowyfPOQ3m3SDtv5euYGraiOE9OXfgWlLXNJb5FqBOxogvaS
Y0hbBlsVBR4BZ+SyxkbMC5OREZSZ9izfuHXp98TWduqXCYSPCiVMg959wJYTdf6VnW9A2fqPIeSi
tKV3akoMwQfHAePg2fdEvoaNfycsiQin0LLG4wZHlkpBl3nhmTLQcD92DIFIOggQdrT6HYD05l4+
x9JlrRb1+W/+tXgz8rSrj+xXGGkAorYsdg6SmeR3oEzJlCJT2yJXh0VGzn1++t2jna5cdluN+nBO
MQ7VwcmGHGOUzAdjS8tLPVi6DID4I9BnKcCxjqQn1g5aOOWr246ijjlgoIL52DmkMP2t0vi4906Y
YrhxN1H5vuL/ADNiHTIG3HPniLUO6CLD0UVaJFhdxet4EyIhatVX6uP63rqrVYwwTvKJY9KCOj9y
gW2c8Sq2I0AQzpc1coIRMM5LHhuMn4fAOxssQBuheAx3CLGKkMXRIUYDpxr65u/TN9DhuPWdieKp
bkH9z6lnFDLkpVf5+jepEEvyi6Ih/aYC/AcRGDocAs8uJRzgbKvPN6SNAZG5O7pOr1ioJAl/aS8W
TY0TSW5DXeULjPM3KHVsYR9X44Y6xpOU9/vw9NTbc+ZKbLQvdwGEJ7Xf4GN0hrDNuz4TC5JsGfhQ
GX6DLWKC8TYPrqgMajeFKcjkawL2gjPTeUZWo9Me+hQKtohmCV7NaBMcgBcwT2xDKeAmzc0jsjsU
50k0pAoJjd/jCQoBpvapRsU9wQm2yHxof7jTiNf3usiJzfXHrDPtxF40uvsMWyqrz4nFm+jjPcBe
uus4IOdjWeOow3hx0WK0ZhBCqahrWNRnbvVWTUI9+VMhtJvpEk3F29AF9gUCLAQZMm30tgvClI5Z
u3ddMRApQmNgqUJZlzIQh6m1wKuYUfbQ+OYYEUgC6T3a++nwTvl6vvGnZ/VaXo2Pq4Fe8sQc8cVe
uuLEJLVXzZkMaKKyNP3KJze0B7PigAHExXW4FILQtCrF9wa32M50HvSMbTo4xzt5Wx6TC4ItWGWC
k0vrVPBkqu2AHCQF4Z6AWi6Y2ZKGvUMNZIVHDaRA/EkM+FUKWhV1hO1S81wGhurVUOKDF+RtMpU4
E182+hNUDCwady11ugW6JGmi3rbuBylCokFolqNvz+Fi+BLSBbn99GKn74bT6zklyTVNHpHwoJH3
vY4nG8aN1y64mwoDu3uoozk6cJ6fytEGYiBkdU9upSOiupr1pONciqoww43sFWFAYfnci8NUx0Z0
jVd33pkS5uMk2zMTvpAhN1klWfdc0ypu2WGP/ae4DRYca0nhhjgWRhZTcUD1tkKvo3EgOgeEO+vU
XaXEnb/CluUY9DmUN+6YMONl7p38HWRbBcMyJY8hLVTtBIV0RHnGXah6d2ls9ABtT6P3t4pInczA
2mL4sgMWmkPTBLEZhrv1YUt1SJDsOk8beOB4jtMY2Sk6uXKq+smeNhpeKXuaK0ZHtN8l5ZBugU5i
kiVKLSUR/iYAVyZoryEvk/PFiSwa1iZundTFPfuJtXO2nDKnOH/Swg+a40aARQMVQkpcpheBE1V4
+cN6W42iyOsCegRJ4AN2gwdu1ksKV9AU8kWYfA7i/JEDH4ZCn4O/qyi5sisQ15XOOsFRsiS8gCsS
8PR4ZngdoBmHg0wy0Y4jsFYYmNTsMJhxGLljiVcKOmYLXYs4BbIGvo2M1Py98FrarkAThlZAbJ3X
fCdB4e8Y6YTILdYljOdS+12zNWCsU8It/i2WN4/8r3/05GjEgUvsjySPauNsZzzIAbdpVUQ2aecL
z88eVcWMrrKKPoTJfFRmxa3bYzfffAZQNfRCVoP/RLN5vu3HNhjz1Tct27uoB3Fk27of0/AAHfeA
WRvG6lqVhihp44ajXwhI/XS/XfOam24+XtdyE21GwEITJG9rlMFl/z3SUib+hcWAiBGYyDr1tQdG
wGPjC/K6coXg3/cYl5IO0l1HVB/XMvM51tEyf9uCoRMEAAY9NWQdccAeGqzNr2AN4H7N1He0k3K8
VamSoY6gmHDkjWVE/9BK3lvxEjtEFwnTqADs0fndBJnJesIeT9WRzK19MQQT6qvkTSLhck7tZ2sL
U9NqNKenyVTLc+Gtc4fzPo1TVyz8W4WygdlaPTvpeFAZ3pSDS88N+9IoRKabOqPIy73au2dOk4gn
2l48l79fyOcRyY0Rt2BEWha4ansZxO7UE69GJVXcQQ2AREkZB7ObivSZBQ7FiYFr6tuzl6uH5uJa
X3HXucajBsUUw2gm1nqkJxxm/Yetq699Ab7D28qXNGk3FPSusbUvJASS1UrvXULfk/2+di9jWcfh
ftDXD1CCnXaq/pPvKRZXy+6pEE3RusACL6RNDsmWPIztYTap7qA3ITVjxutXlnQtgf54Odd5tk5z
6iW2PuzJL5qBKGokUkNwD9I3y2Bju/YV7EQGFg5pYl7ewunuVhmxFRW4YId1aMFaL54+i03yw+VX
XxsDe2DztPu6GSsnarw6aNNoYvgUhSxdVsAnvEhd4JoiGXnfbC0g38aB8lXJ8YPWsSUxjrTlOOdE
2qStjJGk2phYoF5xuzZooz42yBemk+Sg853oxErWwgy3OK+75lEaM6g+iocCsvpitBHYDGv1rEqC
OZjYuYxOfWMdAl0LM3PquATeCP4PbJdPgHusiplLHQE+XxtMCOjJS7pD+LumRM4XSzmqg+YDlR5x
jCDMu7jIHVME++iRV4cMlFwtJwZMLq6HILKGgF544xZdaNlqVm9Wrn7Vy9LQNOKY4hI8P8N7WkQG
DCcnZylLM8Fy9RP0/AJD/DxV+EO4k0+IpYBQuWyzuB2Uckmpw8AsSIoRXGcGlUbHQMx0pRnpDr90
3byEI4SDy7kSCD6f+py98oq+TweDLJmKXMxGdivykkFrAVuRVWj0u5ja5ATqvKvaZJc/p/KRK3Kr
j+NrFD+MOokVOPP+bGbJV7CvN+UzHQF09FSWENXtnJvEDmoCPeUQrGl9y7Kvdmf3agrLyWR9d0qF
7ZT4jVBH4JrNF7TGjIKJpQiEdggBa0mQTQMKMICBpynIrxtHILJHxegcgy3vZF23uIoTM/3WpRsu
bC+6B9qFtpbh6NYErsaz9l2GmsL9+pphErzrHcgee6X4PBcpxQAleWWc2civLcZ0jC333zn/J/dJ
B6GSJk068/TW/0HnBKsxDTYvJaWHbQ8jrASRfTKuUDlvnEcNZMIxmqqud2AR60U4cUXerjaNv55c
XK3oYUZNr2BPHeZcE9Dp64mtEeCHfX7Qm0Yj37hi9eZRrOq7UcQuvB5l2A36VKNhG7pSRdxuQrj8
0tpyfhvWtQ//Rge0op600rq0Ky29XCVjpXF2Ad6BL57MeoOg9r0mqFqzxEsMtWslZlnAwQ3xOXn1
q1fjwipbo+TPDiR0u7lPjfY47LMCjzngbTy4OCO/rlHhzzhasKr24H6VSdRfDkPumIojf/QlUhiC
hRXXLIAWUi7Mxuyom7djXv2mnDqJqmh4wujX5iLKUsNbsKxqFPH11xijQJ23jUF/6nRUJ1hfkwUr
LR9H3WDzWbPitgljZEKhYqMJ5pK/eGIjEEPeZtwfnsPaQwuIWU3sdV5HXM8ot/wY4Sla2UP2Al04
U23K0G0/C6DTJsZqYIgpKqZF3Kf0JMsXxJQ05hUOzGzlWtdqRETyGBPbXagEUk9RfC5NwQKusyIQ
/k3WXya5LDu9Y8u3DTMRG+nBO/Lfk2kJPGj6zP72367MZ0l3ys/hT9KohMg9XkDLe73oimhqFeSy
tkTy7fU/3a1NKelJzjb6QwPBe3aaptCGPq+Kprmhlm0Zznk/m39Lnxc6JPKW8LUK6CiCK7waK71D
z6dOx73hiBIR0ERcJj7/zsUnbvJJggqD1idzJUpTqcASMMqcpPvGAvxKdA5w9Bim2ZkIBw0aWtpo
iBGHm6nzmCBNfHH/PxjbAvdKvZGbsE4VCUvC860NT0OmPdoiebFSwRrmo6yzAuDRMVqnLfAvTID6
Hxm1Zoa8jMSe0eXWOlTgYk12EYgE1m95MR9KjDoyplKnF9CqFeapOmL7hOmSiUbzLPV7ygzeGWtn
HMos71aHOk9y8ER7EETnU45QFy6SgBQOIVuFT/pyZxU90pNuQdh40v22DewOVgrePI65Y0w2wVox
95et5Bf9y5/D8apPXrmXKKmyfVsotBUa/KBW1wpUw1/cHy5gdV+xIlmO5ww1J/NgaQUKfM5GjaVL
aWsCgyMHyfp6uK9NwFb9omsPDz8u0hzFYfSYVID0ocpu14kVcy6TCmN13ZaJIkuTjynn0Fr3cul8
WrxJeFBM0VJSwQ9Uf7gjbHIuhvcKAHCyK6E0iRUgLJyBgtldnCRqO3o7/lLAhw2n1wYyjfiKYroE
RKpv7R3d/vWC/OP0yF7L+9lnma/ACrXTviCAdf1kXN1cR9Y2tw6zvs/lrUsXWrPqTC6QWd/Bmo0b
0G9KCW1PWKRLEMvyc0mWqoHBpuhtkYP74VqmaBUUAwmL+UhGCp7aGfEv7XTp5/tP9HmmPZIxqhHB
akkCGczX/fgDLBptn0x6R110cTq4AXxLqjdkYG8QT3HtDJCrm2LMxZsOv3uMhpxfkjctkIYzaLM6
dRdlAlDoyk5DXs94NkqvENONLr/DkMxTwcvGEZahyrvgfZrsors29+kUPfjHU6SHGDjJ/oTZdhoy
f/yGhLlfIQLhyIR6PHLvw8i4A6TfBKLnWs/FsFflOp9m4rXtBYirxB3IUtgcTmjquuNeysdv7/ih
cQoYHrSCSufFGtDdc78jNYYJj21SqSzHylv6X5FqsVZ5LDbt8wdPpD1ehl2NvB50oX7qSdF0/nyo
cgkDuJu73VOTEFz1M+cEss+nvd0nV/+jkQTkK3ROf7QYNNb/Smgoo5DIsU1OCdkRMIM7dQ+7Fhxc
AM2arHke7R82Ok4phk8ghmd7Sn9gKVr0BGW82SJtbs0jiAPJPb+tHfVasM1HjtN8C8CAqYT8ZmjQ
DXcdvjlXMnqqKCqqo8+4230gjMx9iHnk/P9gW5aKFBTeGvZQZJ3r5I55bZn+JTbk3bXbaYmCdIJE
Sz0UkwNJGF/fiTYJkwT7G2Qk09CSPYTBw/lYMHOGch52txCimxwmN3zyVzWNt3cxYzl6jWHwH+kg
nmLJISkKqOmuHAcOI84S2rRW6lA9rWwhiYLVNImzuNfvbJ3PVeZCxxE4DhV26Uhk+Uzk1Ynikfbd
c8TKHfQuFoZMFnZ3Obq64evZKHlBs57dPvBKUMlL0eP/zUQFwOgyjqnMvC92braXHf7q5xAj7W6h
SUvu14Oj4hf1znAy57H54plvZmzd4IpHxDGhEDFEX9BL24kvbcqj7wE9TOXJcMVzs4hiCRKtM70z
g1tNyLMzb9J4T/QbsuVk4ZNj1v6HWUccAozKRvVwUGtFNgI/YP84TMk/55kZDkij67piuaiRoh9f
dfIAWZGf2F6SODl925xjPrWrLInFUqg75O7sOywbQg2dolB52tUGHVkzVxHIEfmwGr5z4etbMse9
7H+7+0zBLwR5ymopdMCMl+tKFRRs9UCoNRpaI2HGfyTyoPC44qW5GljunD/t8IGcnqlUs2JSdNIZ
8RwLEC8HGb24OzKDkIVtg2r4DBnLgOCBbvAsqLwskNlDRHz/J+pSNRqGgcPrUs6JUn8pJUNxRKgv
bPJVJnQMGxpb0gRdDCIJIagoXWldCyoU5Dvagq53NQTNdqsYPQQ2ewHVHD8kG5yK1Uy60X7JASbq
5Zm6scCnWf8y9138l8LyvDTZGHezrZlX0lFv7lewjG6CGJznau/Av/Fc/crF+qc5dnjZvVJnxYd1
e8AQ6ZKGJNzo7X+XEBeJR09qK4Qz9FoB7aOXT4JVzW49hktHc6L11nMZkn9o8bpmiM1Zkj/CuxoN
qYkC6Gq7OZVJuFNmvxjR1xb6hElLz8KzYQ1U6MnQhkqvyNKF00Z/lBr4qRT8WHSGStS0R21MvGJD
S6f2pLTqlS7DPY9YfHMLAHwwYiYfM7PvQlsmZFJojUMhNYBxbNQolCp9kyrOU9TpL1dUmvq/ZTPM
dZUZ5aGNLD9oGwzHteTjhbKVBpvE2LtnwvFuqQ9/sTmBUlBAWLJtNZioAGyUx6jNYTY2UQPXK7zd
EuYcwRvNMoF4c+w815kGRLEFquefBmB6kb3BpT7wqAdZPQ10jS/NUbAdxuNSRW9V/7me3x+72Ixk
jm7Qhc5A5puNt61trccQ1pFsLwzs5PA2c94GvlKmi9RCMUDaMoNcMg0pv7SK6LM0Ieghmr+Y5t9R
uQmJ12AUOBUM6mMWEqOzH4dICAIowwd02IHQV3oWkwcIh7GXV5fh7kxXFOYSxDTsIv+eTAzbMSg+
iRecQeybhYfJMbUbsckxj/wlil7dv18mzSlLReMoG8ST4pJc78eDGYTiUhY7LkyUX5xgwcSmxxqg
vnaGIMbLCGuaImseu8P95z3Ak/K0Mi3zl2BMlqiCG5fFkfO9GHhnmIUmHy6nw89+xOg1x7MHQrI9
CmRN0pY4UYEv7RJCX7wxkCODK7WRMBLxsI/zeqUCZ4XpzbZMz1Q/tJNX2MWOYEjT2/Mq5BUxLb3b
4NRhpKfmmMGiPgnblUioL8ubIwWz7ma1zCHOvSTceBHn1cV2Bu8rntIjwJAC5ub0iUX/U6XkNBWZ
nurBD5pGjise97fmTA6fr2+T0s5qj8P+jsdupXs0VZ5mb0+k1B9MmMqxmuEasJ/7KWYG7Wu/DsbX
D8cc9jFNZ0b7Azl7UFHA0oNc+PDkEQ4AHrU7dgxmfw43STRYXC3DUGljRmP8jmBBrq7XKB20P4kf
X94EXfzqIQ/ArLE0fQhbvJNwbqCk2HgRUHCnFl0Zt2Q4GMg9kpBi79MJYrGSMbkDLdkKUDEQbsLS
UbdNZc6/WqHvrMzEZPugaAc1Z1Rq2tAYUIXqIlV9cfjXx2rgOBRfzaGbo5CiuoZHK/pkGp1WJYXy
JC75eGJNnh1D/Mls+DzxQT8eeH48Oqn7D6Q3+mwNGMgemVQdvmwjOQb7n79cS6UNqtT7F1rgtZuH
WN4MpdylMv0YRbRQzRTVf3MyVqurqm2+qHhTbRyMXJbh6bHJlis5QqwP9WMpUo8lXLSuaZ9kuhMv
i5l6px0/2OSdDAz3pgZ9EU2jiGZFh/LsYFMAtsKmXk7v4paXzmx1QtlMp43tp6XNood+6nPdyl6M
Nq7iGpoU9ZPB8LMlDnnll9t51eP41Hr/EyVwm24kclJyKCGOdbWGCR4n+yH2aI9hx7Mfsa5mJaAE
gc0NTE+d9gJpdCOMeGiY+gd3tImo6atuQYAK7HO5xIuAY5XW1hX/a/MGeMsdEgoNZkYU9JOIAe4h
QUt0OAA9Wgqt9BkB8OUNgqHDZZAe+c9J6tkXx2Bgz57flJOm/SIib79qYYy9anfkhzxXASXdG8sZ
RSX+MJQe1jjiRQ7mC7j9TI73EpaIxxRS76gzahXDyV64VgRIuckiMLe3tY8cCRHYZzJOuly3k6We
cD4GFIMTiDER+qKTLoHiEWt0tizUYC0wfiN24V8Q2zOG7H5XHCxtmS2ofrSvdu0s5IwoKRNOsPgL
+otq9B/j04CTSrmRIXkeJ5Gf1E0rQaaFEPyWLG6EUqc7rcNG0wNZVe87/wVxei+z6ZlDscJB+Jmw
rwXOseyCfzgArLq9PjPfM5rz7FvT7+h1AmpuQlmei9UK668saa7JYSxvevJoSRzZKjYZlk7vbkfy
l16pEMNJxNGWbWrPVPZjhEUG8IyM7DKa53h1XGF8flHFfGTurMpVKaq1UcGOHH02dwVzK8q5SkxO
VlyG9IELezouLAkn62h9pP3N8JrZYRTNokubG57qBLEq32ATkJ+NuOZQkaCx6yu2jAQ2EgR8xSTB
otQURt2qsnfnJJj9spxHVnDy7NJUX4hQJCtwoyE+u2zlNeY81Juno+/FZMu2qxjBmUSVzDt/QxLi
651xupHOqJhZQtApFnbdPY6gYPZ/lOFROQfeCFaDZp5DcIcoL4CJRoYI0YVga0eUDkaItlDRuSFd
OfHzhyEvdjcAivKSu4w+RO4dkBVXmpbIY8GgE3t3NsbuYbK2s6mDMtLWn+FzRKTzBjoE5XqUJkNX
KmJeFp3/dD+wGIaLSj6t737dd+2lFlkQUILKKNKRnn6YhswnN6sB40dz1XByVrtY0wwyc1yMhjm1
N6horAJus33HXoDfhaembc1c0w1r1SrVlMUhFW8MYV50jsYBBg6CeHZy6wae9VcoCT2yaWydZUsA
93Djju2eSBK72QV4V8ooAk/ZMozhYiSAHzUStboPg9XQxDVpODiFqz0J2IwFVQmr5+h0gzmpPBHf
lN11aSRr3aUJ6R74OuD2WVWa2asb3ieHeFQCi95NGfxGA53ofUgQHJPRvm7alYeR7c4klwkTXVP6
vUSm/SlCwpncGKL+lo3unSS6SMA18xfRygmXiu4hNZ+I4vcAq0ucUz1qMueAatKT9M8SSydxRPIO
VEsWwv6lTM1mOxx2l6kMnIDgLtCuzF59qWNOmZYTFcgW7eJblfK7e1cbAKsmB/mz1fWVg5pVpW54
iCTlIllRr1UdVKP0GX582odZikqrJlPrknIkJHQK0Toljv/CG6RbbLwzoiuU7khJPKSkVvhjwd4P
ue2KwcAfSrgVbRWoVGi1g4kLOqSOv/lOV6CO/O1DO+t05S5D6Mm+AB+5itxzFSSZIdI31FHj7B0l
/VVzxoB08xnWxrxpJHYbDh9S2gu/b3fX8y+22orQDzKm1cF5uEbls8PseXCG5vcFaQwco8a9n4j/
2L20aXbdkdbVYMOrj1mrvj7PoNG+85LgOGRdywczk9s/7WI+evTMqLpA6YijbeqFhMoDeY76H4O4
TDQeVe5V8BlulHdpJPgqB0RpVsLGWMlTSDD+6rOhZdqYeEuPnAmI4Eu7osgwMjbALI5h66EJtkiV
LXvugJRMCz4DQ/FyFHq38TTCwfKaLXp6L8tWPZxIxHYZB2fgm19CxIZv9ZiRNfBi2NL3YPRp9apx
FkSB3B8wtCr51pZc6AFgeVwxtIVYQJiMFpeYabJVrfaB9KGnW7QACXEI3Y1NPm7m3jHt+2ABhAFX
eQZf5M15lKiMLnDas9cQobsKspttjo9J4DiimfT0kl4EnOnEulFyK3OKY+mUA8cgvURF5waaptj6
mSGELEUy0blwWX4/HD7DHGctAkgPh4OwEKrQTRtqXBLIyKgOTN3F1gMwjnYX93616HYEya0oN2KS
hAM0nXMf3pmZLng/dzv9uWT7YW993+EDIzPE36h/zoVlbQmS15bmdgQGYd3hes17mAa3eF4BurB2
XK++x9Tdf/K8W2z9io0f8Y+T5rQtH5/C15ltaVZOxB8i13CYCXB9u8eyYFu4kobMgUmCWcvmCWVT
2smP3+y4Cd2BvKYvl9vFSF9JQ7hD3z/GHPHnq02UTgYNyChdBLO7MOA3DsMbjotzk/n8wCNyi+bC
896sCRTgMdTicHxPuMLNyqpV6tB9rqFynq8O8JQth1W39DY0awNZuyOTjP1kDMswyKghzzMD109D
NHwHT32XZdJjw2irjbbpuWyLtCDIGU7lLIOPitlWrTnAbPpgE+aXonKqNPynYsOQl2aCw1V2edsB
HAGQXhGrVfUdtpO07ssWXmrM24R2/5woEvAZsZHCtjr8APYS/+DOOLrDiObqX7m99LCG7gMM97vG
jSgjD1T0cFi+4MLT5ypyTqRAl69G7HIEVIueM0htpZTAPzc85yCV3T39WxV8NWoJbwo2KAt8uOQG
ciLd9y7X/chuaH+TM0Z1Cr0UIiWnWsiZXh8FWp9B7dDAQqKxMQCVmIRpLy2JexYWnzGfOnjgjTXQ
1FMK16kWRUWj0xcpOOsyzgHOldMgOGWTQcW8bCaENMcU66dYnoRUhM8JJZP1gV+abSzqzow48NiR
jL+L6GRI8lDbLQ8DLSL8zwjEKTADrv7ojfXHryMreTBJgMODMN/hAXKGZoCfv5XpNSW9y4nH61p6
mE2PpqZEnw2UGnb3bGSbPkYuiXdCy/F5ny0LlHW2Y1O9wXOrv5DaLzKUaoL4IZf4bI5aRkDOg/Jc
kdAIpmVQv9HFdq1tNiBbaSxgMyxPw4l/qXMpXklzIyEAR1fQXDdJZaU5JlhfOP+PlKyX6aCqKOhW
Lxj4gH92wy6MqyTkqxKknnUsM6UvgOAIdG35x6U6N6pJ8t5EM9jRUEuZxkhgriiuS9rk8jsedO+H
8WnXdmWLdVbCn2FxWQl5EF47RjWlTNgpzwUAZUHnGLyzubn30wTL6Ml11qSj8IBC3/1ED+L5RVaX
yP+dY4CPTF5npMqpbGwNoJh+LkhrTmeonBLv269G59YwyFa/qPrm5TQ5CvEAzFgbGRM3GsJprtsa
r45UJA/ZnkeHA5KqczzaFWSQzwUz7Kqh5+Yu0oFzUxKvA+4XpXDHp55lvsYM5g0JakHgmGBBeEyw
AOQlOx0H8KiiyDl+JHFga/G6oCbde+ZnD2NLXyuFLk1YKcugpk5svwKNd7VKCECDlcCD3YbWaWOt
FS5NwYdXog6pm/IjpWTzt5MibskhCJny2cMHtCvM3RXtyOFe+eF9oXn3W+WpLX3/VbrvjKpvWE3g
cFpdiaG5JkkHDD8YRTctMFYzIfgpSej91sDQDQ2Ri+lbToqqtHvN2eh6rlxRoXL5/O++SUVK/B0J
TmS+zdEHhekX00ZNApyxZ7kdrYQJL0igDsYE9FC+Pcd95wVf+XXD4yOK+CqIvaLaujVNClCZpncp
DyD13kqxTCpmH6g/J4Unk8GIO95Dw9QnO9TviaLAine+PKXWKc6VF279S0csB/NCB8FT1MAKt4pG
CEd5UC2JKU57peWYbIEiBqlXq0/Z+3H/eWfNis1uWwlMxqMGZx0+Fi5bAeJKty6ncdkRr8tWZGYg
uk6GXG2vogA4241JnZUTs3AiUv/7v4x71W2JL/867pPnCjseeBml6tE89pTcKrVv6zbCcens46+s
0z9FLOXTielDAXUXI/PXz8htsI/hKXHFFpp4XDwKSfiScbBEsCooo/CrXad79f1bHdA6y4jfVQ7M
4f6zVNd5PhqXwADAluQhJQYzUZIiiKgK4LaeeVxIq0IEGnFB1F9+EBpItGOMQmvTm0dMSOL07iSh
OHg4WWE1I8T3Ik6AH6ok2kNgZEiOG0YUr9UxPjHo6JrX973Q2+e3097wQvn/nBy85m6FLH8c4frz
Yx2iBBBQ0aZ/Xxzt+gIz2qB/eSA5IXBejvcLgIEjfOoQwa5vEdIA8Ra4Tr/APzu/o8ZXBqhSKJiY
dSObBswNQdPuKtlrEixL0LPcOG+zG8NzlAYGyBypM7OQU3grzOtSVpaGmQVB5IZOIWfv/7VVl4Q9
edgAj9mVOS+vZEZ7JUSlnsqE0pVRLk4UH3PymZGboOkyDNcXwtLbfyrsaVcbRXuaD4kpk9RHD41H
vqHudNVp0mT7opIWMerbTlKsKGS1Q2vzPlk/LBdQy2CTedfCPYa1Uct1dn5/dvTVcq3E/eTsPL/g
8irJoI0pyz60Rxs0l76Q0BZ3bAxg2N3m7I1xfPltbNg2Dw44guF80unf8XvBmijGFuVu1uEtAHrq
FpX/uencYNG2Z++jp/KRe1ZYxNCxxxjxgGwvQfzlRK1f3HtSYgYKlYqcmVoJ86dMdikPJZ4qiOGc
eSss+QO2awneeyXqkrC7WG5jZugbvLQw9F6ex8jSXv7BJfRo7rFEumepD6duYZ7Veh6W94pB9Yl6
+9zff4iBY3ead7Yq/TasswGwTrIwHT3cWvjG7xjvHvk5/gDdgTbka20WVer4Dot4SS7fsiKY9Qq6
U63EzVneq/4VSI3e0QesUxzYXs2kquwWIz0I391zCi54qhH8XTIyHQzZRXq3am8zqa8QlWodHju9
HX4rYIAuFYcRxssJAIXTkvbVto7wMscXJERoU3u0gQUcXiIEkToCyqSgGnp143PlAdTbQWrUSdkD
2SuuLxcEgcc6KcqfWlzPskCZBQvpcJ0IaylMkfU8oEiaWvg+6vnTi8Ue4Dq134bVgnlVg1gv/NFf
lfI6KfZ0tj/cmIMC5SHjajVGUt3wyscLa7nM2KXhwmXcl0FXKKjevBBG5grndpoY6W4Cr2aaqEHl
V+YKEahzxpZq1tP3NF0pjrjINxhriTfC1hexkzttixYvbEv47yPyoj4pSuvHGjOh4OMSykL/EbTQ
86dSpgl58/DjWqbDKGvgpIi88Pnx/vwOPw/sspmc3gDRpUGLPQ6MCL6fZC5SEmHRThlPqc1LOurS
a0tOFCaSVIXIDEuh9x4SvBNduoMJ0TEyKkbQ7mm9LFRdVOg0R7GMnwoNh0YoQ1idEghFN+E9+PCe
DBiVcqNYVuVB5svi4thpyvY9ei/5s+PjJQAQPcgmSXsMkA6Im7DjRY4qxe+PCS2vViepM6c3zb/n
44/mkGJqLLeou1HTSWoqrHJ1M4aRvFQbBHbSwTgipFS1VCelQFmmLGbcXFK+hqDlXQ/uLIJA1WhW
w7LISWtMFsOBYaANwgmxOfCIG8QnC0R92NgmIKGXGHv0iFP85sxV7dsQ4y/pRHvlM9pf06vfpj6a
ONaHmpZhDrvkd+P10syZyF42ERWLa0aGdx4WHdFy4Z8UQyC6/73cWUH+pr0lUA+hOGymnRRFSU1H
zNlazgngB0+7zOVcsvGwsGEx7aHxRfz4LQOpetd3TyDztn1Ew8vIhcmPRNL5TRwxL3hkzC8TUGtX
354c9ide4QKu+ZfTd262kdJg1b2I4QvD5m0/SPFP3Yn6OkA+5e6yi8ah22TzIyt0QPsWKvnqFmON
ZmTU7Z0ylPP2rnb6qRoy2cM/iWpslHAEzcw0CU53NhREeIAKJkHHfB88odHoUxYs/4CUfS7eDhTZ
wkTD2cjAiQW17HGo/36cyJnrfHsHz4L1klRcvg79txx6wOqdDsC7hBm+Fqys/8MHiF6XD9p3A4dR
831eC5eCF237bKLAbqdHGyluTYqi4qmO7hlmB/8aOPHUikoyj8ZKlFB8v4auZTdxu/3D2sa67MBF
tFTv4zxIT7v7vgBqbqljEfuAeLIWxZY1jkTevmwGaeTqE7O2WUK3vlYpavpP3OEG/Hu+Og4ggsFc
ZZ1lsnnr+VYaltIbxCMR3ZWjEJTVIZmGBtqg39Il8GAyC7EDEwmydQSFVJu26KAj3ZtW+q6Ge9zY
jDT+VB5RKCtssfxlW66Nk/4pI9bdeUiL7rLkva+c65qx04dZXJYaGh9UUCNqUL0Sd8dgv3aHvVd3
QWWJug8zVZfdTdDyIpghz7yPddjRZo1cz/2DXau/RLZq14i/dUtw88ghPqh5JJMllXNEPVLUA5DS
7Q2ZfZrTwjzUJoMBWayzQ7mKopytiVBGf/Ui0xYP7VU5bHQfIYoZHPe70ovcRM94ShV2EpX91mGm
9aqDFZa2946xXMrClUNtbzCMFSKLrpclgZm+bjPY1CF4Drg+DJUgUHYnmqizBRCEW7FbFbuSpYWN
QxYAAb5vi3S7LJ9PGY/OXpGugfz0M7GvIiML5krnyZwMFkTMr/qFMPdCaHUo9TVTCTtmogkd+fle
dv6SJSlqgg661nWxxyZirKhnNrNtq29KBLP8RcWdRHvhft6/SY4WMasvAouCo4pcAs2R6lZuGv64
G1EAnxyeSx8TkaaqiqK7qd9DX8DKq4tPEGhAPD7DQm+wmskxiXN04hG8zIAG0j/3Okhx6qr1Tgyb
2EZ/FHmDg7+oG/WXRnruF2XDW3TGbQhShMDwrij1CT8SpFDMAzLzGkeb2RtPaV/wUbT1u5SndeDm
hM+EWGd2o2AdMYjdR0nUmBrnna8jbQfc78HQgPl/p2ReF/FafjZBtcw+HiQJgIjsNR0ysTlBbbe7
VpV4Z/y+NG9mohut+mdNt2vgtbB8Jt5NRof1oI0qYtWHdWpv2YGto8sNkIs66PrOHHCsnLXO//JX
6q2nA0UEq+Y2NblfCFywq+n4rybsV3z+svh0lOoWBypV4H7zVVcBkeoEyYPNlnePCYLaMmdkQIXL
mq4a7YNThwJ4JPrWWqrMcG4f1J9NQ3bIgdFIT8qWDMl2Yi92cVK2ZYMBR/YJ4dkj+bqxRoW5RnB+
0VHafOcZeXBeiblY/vtP2pOiJTsU3kPz5mSW54EyZok6dWzrqFjOcO6wbxRAdbKGMQcgUZ0UoHMs
AT2Kw0oX61RIn7Y4xaMty51KKKjxS7dgXYp+3PW5HedjuIOyZOClG7IarWiRypId1583FPQU8xac
pwDGRT33QtX4GpkyJA4hNbD59YKrQLDLEGBllu+VZw34QNwoBDTLln5aoHWsewlpic3+q60zGGFm
0bYuApYQSWgFTF4854wAELOkOvylfj0SkkZx79izpiUqRjgziWzOQvNtLWALIGQ42cdpPxvFOBCm
LsOG8OEodrG79po8fiH5Yh4qbGUrLCDEdq06hE5pT6T+94XPkFC/TFsPRXVXt8UMdfx8XvvPEodx
bMNueFKrCXymXBotKGs+z5CmVDCC58rbfxPFK7XOYg4r9FfVN53XJ5b5UjqWM1Opua5VH+Y7/1We
pu2UfHySQWbJ4yGwCuRnonaSR/owEkDzVYxB2HbQgDGj3+Rqce4czNJBmqy0AMMgrCU9M4q11HXG
9DHk4ZlyhGuMGwSQqFxaI6W+syKQBxT+vrExhSBLFgh+mEMuWrF8YG5wyvccujRu9d4vF17ayabh
xRlrogvB2b8E/m8/lSHQC3P0+vJKXhgUtw9GA04NFvZDpZTksDvl0fDNvVgZ0FvT3GSm9z5Q/jF9
/8rlfU+PBr2g+zakqeJKNYmb+xxAxJh7nZ9YTSqDpFtTJqv11C63DBkukrdr+TwFCCCZQhX8iVzp
0CNGXc8MxmsjrtZKBbs+DbKBQO3pVvMQTseHcLFc3G8JHrTr5UPOhNij4PFMLmR8US+ltxumep2R
duoKZzhBx9KKB/G4P7y/LZTmkMbSCZfLozKFPnt2aPq4vX6rDJ067/BUK9Vt5EQ4ziEB6DLtZ+8c
oo9+x1lzqYaD7IiLepaWHelGILBbstR01eeAzsg/OxYI/M3Xo8Sm7wzqgrCkttWdCVNEr/ItnhEh
KS4eK1kjWbuDAeyViDlPQ07ehSPCIm+Zyn4tCJHG8CJhnRZQQuKSDoTqkTvba4h5aDKlaJxMNz0u
Nk0tqm9Zn3frSVaNTbD3A/45l6clzmtSbchM6Fc8ChLbk05ksywrpwv11aTywvZdCOF40yumUAh/
rJWPtvG+0F1ycZtsrPDiNItERHPluyPrvGaGnHSb7SXpLm1yy44O4HtMjWiMu9f8U1cilABVKHSN
5a9vedXZouT3D4ENrd+4RE3A2Ck7Krdlps2G+5Xiz+x9zeHES16ntKSRJsc8p0zXgz32tysSvMZ0
DnZR99+KyBvjH2fQ8pR+E2xtTLa4OCT0MYN+cwGdHNI6Nw6poDV/Em1a3Asb/KL582NI1REbNo2p
flkg4fzsO4WZJBjkz4876Jfy5YZzPHOE1joj7HbEBJpMD6DXmPwkU1AMj8ZKhlCLesuawfPpK3ex
2H8dNvIArs+aShPfpNlJimjPdb7fGqEzxEpYW+nWuSKTwxScUSd1tgVsY7Fryq8p0Dh9m2PP4WdX
yAp7QlHeFJU5Be2QQxHP4aIBzzAwprGO5WYlph3B+9TCvv53EjF33TdWrJVxpz49spbFiAxzkrTh
npHftSoOSlBRPQUl/rTfuiuMpMP3FkABXXgGjexmfPll1t2O+l/4b4y0Zc5BdgLXsH9ffZs3qYCb
7ZlERZzyIW7IrZRwXe9WOll1ick3MVfuUEhoMfGSzWSE5MX3fKyx5WwFATE8FjeIw3g6OL8H+K8t
QiAhNSzp4CRgC1JfoNKcbeVpxsdMmqkKLmCPBq79Jrq4GViEMwnYUaE2JKsSw0c/+BPcf6pXIaGy
e//zkYJswuqeTT8/YupUiasdzCIPOomv63HDEHfjU+P/dHWcpE50q19BdnuWX9fFt5qHCluiSegt
6XyM2K2DpOp73FRl1UcoPda9zkLDcRFFu7PhscKfnSRv5dYcDsPGe9xcioLEM5ru3mlTI6ekvxw4
9G8g+UXUkFnoC9Ql1Ux5XJ56BqurOBc+WpM02Bv9NsNFk84RjxLKMoTT8oA1SyXbxdVD2jPWbiY8
68ji7+XrIM0hKV/ZPnbgJBcbSOTHkMsDUeeRqa0b7C+WM4N9fREK8xtThrC21z+7PVKKfTlg0Q33
ZzBJsSIj6nbLeA6jlcKKClKKcxrZTa91fzOm4B1FOz8BvXjK2PluGHAkVItPjkwZHB9KFwPaKWc3
nCWmXjo+zFCvp5l5WatZYaV1+WZ9Cq1/N6U/NajVp6ZA6tSSRznG5qLsNaAXENiz2N6vAAcA0juE
7nMLpMvYwvU2Q4l+AAlC6LhBozzqBDEcXzrKSaIQYVL747D4G022uOtNevoHyM6Mmg4k6Y/CN1ek
E6/fH/JFR6+WAQ+HT7rxX2YgL6BoRZbS713p0qmPDwuIvXayPN4JUrbI45JWv7clBXDKxikJ29fp
SjS7PPW8uRYKhBIp4AG2pXdpDYmmYxzkIKlP13GKt7Dyyp+QBEuAbIlm94iW8ed7g+jL0a/UgZEy
AMZOHxQLueOIuOge7E0LFsZBDaIaq8RkkfBrdrLr1PNnGm6pPvtRHHB1iDQ+cTJiLPqdg/+cuS9v
nDLc1llD8//YQv9T/zVFwOa1cZUf0cYR8A4Bw3060bXQfTeZkWZDniBhlb/ZUM/2qKkYFt3zOmHa
LnYDjB1/A630+h8ebLIIpVNNPwbVHKqoTqcd9GzVtObPjAoLTDDg/jUXrDTm/gPo4qd/sF6BCXjv
TSmfL2Xko4krgb/XC2BlyE89ADjKGlY0/zD4cRbSZiGVQyXcIoc/wUUy1CKX+HRao+4PnfNORlNS
iudVhEqZH1Fmo9T963Ad8rJL6Hh8RPsyQ4UGtL9TlhOa7l/zOlwJ06U3H99CD4tvwhK7kq7ZbuS3
tXfFm8RguJGzC4KXoQxzmjA9VTV7BwAdyVsZSJcfiAv9z35QCsvRXrTEtznu79Fx1qnA9QnFFGJi
+1QOsaQGpvhnKxOAJSxojdkR2jaGUqMsq6w3zaUYLF/enILeK5uVes0OJMsTbKm7SeZvZVQ8YluM
qSMBRg0eqLtwEnaTj0zdIQJvVK8nceFAMd9S4OoBwWBDw/g0gUNLEkV0FdutnMhgg/9NOcCba+e9
vZQvOG2/f7kANdHihqe8rucN/7H4wOJSqo5jsL14JUMPpOFV4XU9NVVubvjMNs4CqPPv9WuGJ7Eq
sjA2Ag5uC8PW4+cS3Waxb3fWQ/B1AJ8445qwBQ7XcsHgbxqf9VXfbw02alaTZ3dvwzJT9meqF3ZY
YhhsPxOZN32ji/NtcNQJReo7cXBz+Z/aAnFPrzM5Ao0yYx+ICD+wmKMz15qAI+5ocWJHtwwu7Mq/
M5KdkwAqzc8DbbWbhOghmkegB6KI7b8J1M1RMTGfR7fhnyQLSU/5gCHCNGguF376AolWIMByzssq
564XX/5tt1VbU17srPfftcSkpJrrDo9M5xXj49CU2XfvXRJKgqD+33ckVo6EFLW7H99l3/qrS833
PiQVTpgrgWxYEntSQc5rELjqmnXKNeBEL/jEMw6P5Ii/M5M8tHIDfsCvmTNA9otq6wy/uY5XgNbY
8oOfnVlSLPH5CEuX91hA3udE58QxdFn+0xa/4VHkqDprbYuvWcNEc9WdWQN4AW1R2N3oM4aGSI9u
tz3LTlYIQjbfRMkMJKeUVafsI5uoX7ygX0c90luZhlx8bG1Vaw6yr1ia7+DZ9KsU+OkbYCz9BPqp
alt4fwdNxSHk+BtiskdL9iOzR3YMYEBUQcdDIDskt8qfxtqXuST/IA1wgkK20h7eVNidEEJif3yU
qE1JLJKiczFUkyrfmUDYaq60wJxCkAXH9pW8ja0kpaqVwuLN90isIP/4ArKZ+EDkgNllAG6Ps25r
PH5bPusVgrJqU0Bf5GYSMwr4lC9a8M9tmDKjp3P4/Jl0ggbOU1l5o5JahxHg58YC8O0uRhYrs77r
L6J+T/lEh73kwYNz5tVxSinTBiz12K5HdiOip/c4ARyBwwrNuGV1MveBi4OSwQ86CAt7lHZ0oUeK
NCRvJ2UE6i9TmSK+5yheBOqZgnh96xs6+1wr65qto7pccv32OH0yamx+hYzgiSZ8QdfCOHRkBsp7
lsd7mTTApTEDmqE5aio+vM9D271WjJZsCg+XVXeUgim+BQpQtjAm0vWWUXGiEv+GbPyaKAu8UFBx
5eg/fqfVslohDWEweCVm6vFZnz0RakfRTlcNFh+h52OdW0X+FGaLsHutwFuqZ7BY+gZcGGQ9GoSc
TG3JMuAhewZWXIWtSiUXsiyhrXIs+jSMzzgYMfnjFZ4ZsW6yiwOvLNy3Fv2IToTxvjkyShkw6ubm
gMmkkccPESSXn0gO7X+0RiUbBhOe0omPnc4ql+YptwVz4GveiYUI1RApB7K96SHc/UWmT/UK5Zvr
EbLN76mTqqRTSjIX1WgovToLMVWYPpxMN6Gt51q1YG3odVvSDjTeKn18fxrnehljEQAKj2L19t/6
jayoHXTBfXg7OF1sntXO/qm/L9eRaotcUpxLi9jfdGqI48JwWJ3HicMZrH+bgcFE/KbSsCzYcxLz
5WMewKbV45NKtRlO+31ssH4/ZSYFQ2jLwyqTaHFzObRicCawpaovUqiobvFDwE20nWd0XVizifvU
3VbLh59HTlNKOubGXeWdAHQ16K9MtdcU29huhdrbZ8Fd3qLPA44Di6SovfGC5h9SWciyJGf7RjVR
JyS48LYDQ41h9JiQW52gMHaXqknzS/JoD9QvbzwOVINzMz7H4ESmA0SjioeTLrjbHhYVHiCsT1p4
4pONcfm+dDccHqSNn9FImSE3HysYphjvQosdAz0q3eN0WVoOJJNRk6wZZPlI79oPH4OH5QEVkp31
fT71qdFYrvar2np1CUgdIdR9E7z+mcSPhxVcTwCO6hC6hGYULUUhfydOBabIv52mzefGLLPusiKt
VOavvjfwtPZjO0y7jNSCmu2VqnNpL8yQzh8Ok3cbwwUcYmm+vs9Mn7HfrP+UERNmdCMfjVpsoNbO
w+6vMeSM3iYtHao1PnFAIQo+u9BE7ZBvLv8lIMufWdKoBvnYQ9SSRf/ukEch6sEYYR7+3DmYyaPY
Y+mpzWs+Ff4orrMonOYq/Qax6qTI6HwF36nnhyqObadwSq+0hipJna5HRfMioAnLRrl6kDIncdrZ
q16ad/mexJOwVDdDqX+fUSFs9gm13O6oZ/6ENYFX2u9xQQX2Gqi34eWFSAEQpMj6PmRsk0zXn/Vg
9Vt7MyxCbWJ0UuDOBfCkb5oOKEVPdsDlt5PlTjt+ArjToyD3DYSkLVF0cikohZgZyGUNuZBgRxi8
yFzc+g5lQlnR3Fz/c0CD0/bsD9ZlE61yZDI3zPhUh3hLR5SH7BqOYMoopSHMRrPiWCyE+BJMb12R
zQpqd4FZLrEXGAS3uRPxvjw7vKyZGBw54FnU51eaue8+h0Avqsj26s/Gnc7XICNr3DYiYlvIWkrZ
PQBff0dqa+/b0ZGOc2q476OtC1BKCw5kJKkWDtQ3P6jUKo4KamDp/DmHwmzAfH7eYFcd4KBx0cOl
8PA8vel1BUb2mbmJ8eHTp7aMUJyhmEMnlccIDiEqpM62x2d3ty07L1UZuX6NO8EZwXDzdHyWOeFa
QgR26mfnnNpCMnIwvbRPzvw0kO7sNl+ngwylO4+3AwwCXWRmYYYjLwk8W/wUXULLgyOBAOu0XSZz
qEn9fZicmqPeex34/T2ckxLnQX8/SB3g6fQJ8UuT1RK2P/MXH39I4khrMjf61r0R6aXMP0rfgrbv
BWy73jNhQrmt/0geDfrw6MBoR/DpkW+O0fT5xBd66/Frz1KGyYNlTNiT/GAkXD+fqIrSmAQYHnbj
lXvpkeijbzbW1KlMow5f/Y0VqrCbvFJxVgU6mBNLpha0WwIMUz2A2eXwzD8qIwWhWysM5L2+Uhn7
dedKPGSYJRzz2ma1uJjt2zFuQKJ4NXl2sE7FVRMv7KvVkS5nkaImD7svn21jS2WZPRs+TveMuEhr
dN7CPK+OAyfbpTRiD8ZaPLyF0qpQkqBS8NxjJzdTC7SU6iRSxVZxYabh55F4qnbEjr7ssRHsAP8U
IDM3nENuRTEKyhs9H39OiumGgHxfqhqXNLrUSfRU6DyIKJyepr13ItGF52uHw3Bxja9NYCMnktMU
9vkgn+lf2eOCcaJfAisuSGN43n8FNcqQzxpLocqygplDpYtl19faqczHBrw4flvvwe6URvf4qBpO
0gUJdTudF/1VZhxZgESWbgq7frB0KYJrppn4v9pexqlCs2kUygx3kmkQMd7Vb4dWPfhOkYCCjiBo
/SRpv3JRaCPytKCSsUKXMY+u4JbFPACDkat8fLuEJvx+hJMVIhLIzVaEajPE84bBu4PRUf8nEAAq
OENc1lwPfhfu5KU8iKVJt4Tq64ZpcNyDLRma0oyaXw/wjulsuoKP7el0TVVGYNEYXpjjElyoYwyZ
/U3pNKswa53SN1LupTBwK4t17wpzrbWVAeGCws3ZFpNIaSGCVYkj9IucC28iv6QzZq+bCUdxJfJ8
AYgid5+gw+FzT09q0qERXa7nztazuxlBYY0uB2Rzb7yia7rZaS87JKphxiznKPIc40igKR5NiGYZ
udlac4ix3XH2j4/vd9MmMxThAm0xMQsSUQF8AcYqXENBWgv8YwYZBpMvMx+/nkS6L8//FvOn4KvI
DuVTI/KunaSjd6nubcxvgXDuFDsbfX60YvwBw1+NVTMg13Pih8oVNlbJsm01iLgsTc4jcGzA3OLd
wePqc7PoQoo+a9GksS0CneC1U2LYabdEIdTrbKlVUs76V0BD2hJwmh1oRkP4PPYp6FtkvcQtcIa6
yJDraN33NF9ECBLKEcDEWBEuGROm5sNUTd6juEapG+DnLYzwv6MgHCm+SPnKTZH/MwDmw+ta3AeL
E9PHNwK891ukRzeHjR31KTbM60hjtmDZxAV9JaAqqgEHQCnZyOs42Q99qyA9yK1Gj7jyDngD6Iiw
EUBxOI/8T5b8Hms1Uz/Lk0flUMnOjxwUTZAaiZ8iVvPuPcYtjxjO61pPOtsZzdZqXN25QdBEPp58
WDTsQTYTt/DRvAj9QsUs04FCTvab1Q6+5boIP0LMnvpGojs1khtxyXmEF/JT9oLYaMQXnNeCLsJG
DgqTlTlmDHRFUPgx1TMWuU7ihLxr46LEugkh7aVm3NwnMi3C6pX+2B8lgZMsd+lnCSWzXhZoMkvy
L0Pqo26jMkC7M1hbbz20eaR7hYTU0UjwwaokUnxYSVI4LZhN4KpiyTRcTihVVjHuO3kQ+1MDoy13
b58ibYaGSnk9ujQZhiSW+sjOF8ioG00WqDVklRCaWV7vCj/imLGT8GrmeSXkOJKZ/IW5vOfHGX7Y
pqLsfTwQtgqbSAn83JnBeMdeCT9nLzKIgbBT3KHA1Tp4x1rGb2kmP9nBozh7if8MUI4W8vGGNFNx
1oDAkdX2pqWfZwaqC9N0d23QVXoR9gLYEf7zJz7LfNVli7iHH/eHSnx0OkWd4I/uJuSQbZyDG4nR
+B0ew72i4j97d1HnQJJXhvdKbhIHLjelv5Nf9jgAoKTG1UBJBHZgXE7U4Jcm2VuF95/wmtlulfA8
1Rme7L75N5w8Ycw1KDP2Xgx1CJz2Ssw6aB716jwDAcI2iKedLiOS0uMgsiYHB2PnyR9HjGmA48Ug
CToZOPihzh688R+AWYB8clBC9P5egqg7aD4IYpSHRebHOmMHz3j0uOfFeFJU/7QknyEoZXxykA9I
J5HBi7FtLe+dMDgdhx/JLKcTnlTsIKvjHLZbbFDT91jgspHq1+x7HM3KHgprHs5yw7AbmaA7ODHy
VavZq/Ms3DXr8An46EZ0R7awZOWbK/TA/LzMia8z6En0G02yXvf1v22ZWxr1o5vUJ0wGz85W4D7X
ikmZ8N6CZMpb6OOLMrwXikuyWrFX6mTwhY0WyoyGfGgstCqDuyB1SDytCb+W6tBoojiDFUFLB6X8
GnW8OnpXMsXPPKfCEjq3Nzf9jhH2pP9zjB2xf5yf95T7ewf+ym2g/vWNihUNzyFfeeZ4quS9/veQ
WI5+TDEFZyYnsMw2wJdXFhWzmzrcBrncTVlk0r54LoPYUB5eM+whvKjY2rWMKiew8DRKtfCOEMXc
4VCXMwHlZgjuZq2RUVuTNqgTPT5IYM045oxL8PnWsykvhsGRzYpw90FVQYA8cpqRfudqBVXLtNjD
ncvXW6meFWVpXRqp7wpnSEXuObtGGfBbQQvEdzbV7ugWptRk2+gNSD3ZDn0kk6NxCneZphjpPy0s
UStXuqHOi1lbC5TVyRjYSSEEahJGtbBwkS3EPCjWN141btyZ5WBJz0iH8EsU2Nn9mcq6U1QVRYw4
0MleqWVlqiwHYXpOPYVInRnXub0UvFb4gjrO4hk+Lhl3PPY92zuMtY8s+4a9fNCF4v/eUn9h+STX
I6t+jbeeuGBXMb5W+cu7HkjFUbXGcn8abRoaNwRHQL1Mrs7wvW3QuDDZIuRu/92zPqdhjFR45u65
6RjhTOCpeqN2twxb95scRKv7bvTFPp6SnBzJQ6htJl38GgDIgEqy4N2fkSlTHQgptXtQSUe6fMs4
2N416gey3T0nOnNdFd0DLf3iZ2HBDf9kHcEhmyCVkxW/pAX8YXtySpbVW6MydNNQUTrFs02BHVwQ
hQSWjWRFFn+SAjnM67CSGau9v/kTPGAbmGFnYawhG1g5FOWwofC0wryO7gsRTyOE/HBKZcw8/y//
LoAxoePZiMIler4BEpeBdCA2pAkPwwQalpvCRshNdXHpKIET1V5sXKPYayzyA/bDJFAjmLkgCSyI
Wh1Dt60glYcAu50pyhDNhU6MclRedzj99m9WX8xjjQyWYkbzwNJTiDKf85Qu8HEVZfhk0M26ZP22
v9F7k4ka28d+Ae8SWt9nLQrHjmD10VA2rXpQnWkJh8CMT9WzFA3K9mEm+CR2jY9qI/dGVn2CkPiy
7k+/2tQgFdb+7KX/AXuQ+0ZfHLniORl97Qp/JK3TNZoElbzufrFJTeb/eKLRNhMN0eUM9O0Ye0Sf
lb2Mcdv8TSyS3HAtzCuGwnbmwhVyhCXhUnHaY7bN+Aq51Zoqd2NmX1Z2k2RJPRFrY7T1f+4AlfNg
5Z03vZ4vbMsHCHtg0fsqasy/ABaPlHuw2Ysw0ZtAdXK6I/i+4K98bDDD+YRqqm4cr/84ZyLhprnE
PYDImyC+LMEuUqeqhZV8/WKa0G7Lh4e5Zo0jOlBD94f9JZOECR2i6JI03f0mBSqPyvYZoE/eLl69
HJAzLoGiutRszBrPHAlbPk0BDXIJYSmk5lPwt3gyolLLNZcZUj1UhHBiX54SHOI8YavPxnhA+N50
Mc/MJ8tOkZP5byTltZMY6EO2S3ars11kiTxhOPTgjj+7cmDEM0bjQD/RIbx1y8CbR3O35I5dllwx
0u1qQVbC/Ri2rv0wLgg71IhRHZf0uRiSTInUNYjOBU86binIx4VBLfVdNJ9s9HdM2uUrXc+HWn9G
4D1tcL39bGpv6CK4D0jK5WCYIWlYQSew3Mnqkcfwm7Zu0Ml1jA50mTqF5/scm9BzyphppbEnIXUF
pOvqnRUKJODDkPDmwbkVgE+aodcJBy+IZqdOTAJiqj+dgAa9MCcCLg42DixRXeGQa7XXVt+X8Bti
1AmO/ZIWc0P2Hcy2Er94lvU77HoaOZWeifHXHV4i+0J++KaXEpP97e83X/1O++q+o+EYMxE8OdKe
GPOtmNtDfclrDvVMs38FKx+3h2apinoZpJ2Q+AK6KrVIRsygemalMz01vkh9UGH3CoIuaQV744CU
N/wzEn6GuYPOu8JBOSkcprc9NVsXOWT48By/5VRVUtfz2rYv4EUOcP6tZcxvOBUO+iDzRFLGJC+n
3ooi2fo6Di6BfgvwDKsTWBaGvlhTi7hZ9xHzqUmQWBoJfbKaqq7bDzxIwR5AOLBvD1vfSNQzawEx
soicmfkoCOiFph2coGXIRilWeeF2aZcpgzHf4bt25ybyao3jZue2QO8uCfsz5Dr3ygspjz87FCZi
r4s0ay4DKKafeiP3ghbZZHLHrEcLUFbfxF3BbIGnCk1v7JLAmJ0q0Sy8jM3KM+d4pxntSunkaguO
tMZJ6pmK+j9g7X4KWifth/2QeBOVj6EZN7YleQplKTZjrmdhXf3AYcByfGOJJ9qceWi49DXuK4dr
kWamTRFXO7DHOcO66wEmmKpnsUeek0IrDqZ/ppH4eDeCuyyULNcOy6PNh4UtlV0551Q4s2mj0c2S
rIhcbVcOi/EmXGFdL0cl59bZAuHIduJt6UI2P4PUpQhmhL426SS3deVd7Icdq0WAU+cduzdlRuJH
FBd8DLSAYGHnKOOLBWonSKwTw9Mtwp35qJz2L63EJWsgnrHYLHMK/i8D07rMmhcdEBnMDFAu6l5/
pMAUudHSswQdFJYD9A3X+U8n8VzbpzW/YzbUiQ4179lC2nR0kIhFAfSGzMhAdqTpuRyOHdu0NxgO
xbfSiVfK9ZGm8UrHxZ9iLA+Cj6q2Jqz7ZLgWTm1TsTd00CBMgtaL8X92FVafJyqPJSsW0UTE7vOV
QKE07YOF8x0Hi+hJ4uwfmjfknbmOx7mipSS6m6ZRUk2btdyTfcN5f7ED1EBXipQkgqhw9Cp8peuA
qtWAcR7eLhloINAzUadMQNTW+ik6G/URY7s8OlcpWRKiAAgh96mpMD6lSwMkBPCHsQ9dc8nMPxKr
YL2uhZIjceOyMtdA3W3KVAQgFlPS+is0+Os58BjrpwxVd3QT5Q27Oqu5Nwjx2byi9NouKGZy+6VA
Ay4luNwAs6KjJ7aYiwHAPwdUrOLh4BAk6RmwjHlGEu+0c7dUYctx1wd6QauqVoHkqjNBLyD7aDRC
mU4JwPhT7lzFtIOQ9kq396wDe8b4RoWPZTXY6T5E7giYxK/5/kgp0H2Fp5Sb3bTzi4V8992Ufbhx
u18953JHtzEoqdgoK3UzXOuDFGWw/FwACq6gnWzAidoQRV9VA82mqDaVxobCp75SBwfkyg/nTUVS
/zbCJ2HnQ2Vz8kJckIoL/336+BM8Tsj83WCE+kQzMNo7kEPziwjgX4fza+5rC6KfsKsYi0NQxpwb
FEVfA6dXPYApHR0XH5TqHa9Zvf1qQupkjJAzhbQYiTIaE5ZCovvqyozJloUtMIt56vIsA9dQl0g3
s0PdGnvUvUetia/unRrrVXa0hZV0dJ5xcFJlhm4oFxeBn5xafRQ3KpSU2TbVt97JP6DyKHDsLh+4
yIVs/TKuXNcH1TINLECk2An9jNqkG4ah9xM/lcPmddlae1SVHfaxqea7fz9SO8DXhsBWjVRjGkjR
vLXK2Wi9LTBOFh18fzuS2KnuMYMKI0jt9VPp0u7WjRlgBg0WMevmg3n4N2TWXISmnDi5ofyVTGdE
mG3NzpxPPctCiGgoxe4xEuMhaQ+KAirRyN/XUpGEWe+jzyZZoHr4qA+n5RMNf28xZP61I9NzBsvx
OI9Tbb61sBRa/h/OBnPQlqpkKz9MjkAC7DYbUIiU+tbVz5d6IrgkhOGKx/Mx8jys/AYRnJ7e3txb
PWsQmD1YBTPpOPhAAZdUOkJjRrwcrffALSVT+qlRuN3Fuv+tHZb3AuHOitIiLZhiLjmNASR8nknF
S3XxFdudHdzvo154PqKL0zFVZMk3RWy+67l6AnNkXt3njmUZlqHmAD2OvNm7D7ZRwrf99rfFNhbO
PZAzPekx878S9S+oqCHv80CMPG7f8baQMzVKf9dheq6qyYee5ilzGqrE4II7BIMPAk6jMN65unPh
GUL9mnMwAiDZqH+c1CQG3iTHMqRLRsAHN302/0t8o8Q/SjE8sN0nI/AV//rwQ5hah3yFbcV45YG/
HhYDz4iGg267K0SNwGZNa5ZSNk/EJ+Q7ZOn/L4YeRcO9/dryfoFlk2ucm9EItxCOU0w4sm6oTPjL
+GrqhY9j36yhVmXTFzMymfUUzFcrpMxGmkszFWiVhhk9anYx2YRJp0/6DLgCNuQfhfZpMt1Xh3gv
fdZI8HdEwIwbJ0ZdeETGR7+TR0+b/j64PqmxJZ12mC3avPeDEBUSQZAMgc3PvUaAJfR1nbsjHaHo
po5UfmTiL5KZiiI7Z3tohiKS7MNVi8Yavj1Z0PipWo27CGAbiG90bHDnL0pIDyk1Aa8pPomjDRsG
YezisnZ6TzKFi1B4Hdd/i6Xaqhd14cuNl4M+4zHYTy/boOG1TNhfgdJfQge4afWs766J5Op7v9z6
+bZEmoU65rh6gHnIDNydvWN/LEW3gjoTdGeYEU9xg01XUuABZbGfwwhgBeRL7lolrjkN+yY8kPuB
6/YMROZ2hgBhAhJ7uDR6nbiAO3VbWCNBpuv7l3zqGr2427tGSnu9bKUmoyiXk8bl3ykmAbOiphW8
Q19qlVQqGDz2Eu5N+T3WWNIXrj6Gjrjk2vJw4CW3SYC7N40BJPH2D5PUeRh6SDMrFnIk8YYD0b2f
ovD5QPPCNqI34Gnr9AJ26tV50d8UxazjJ88iJ6++0Rdv2QdVMfzW7wcayWWuHDpmXPNfZKj4xGAa
i+PmebyNEHySiK7FpK3c3k9S7SLnQ2eCpbmUcnhlF8zMaXjnqLwH2JLNrL5r0yLkAIbEwNQrkkqT
UD1ZP+AxmhR5OfuXxt72KguJa5Jx9pIBs53RP/fsk+NKy1u6SpGdHrxk1valxTG4gcNRvNs4Vxq8
rNBgj7Jf/xvTvqTB7k2yh2O+NITOExJ+FCnBH3WSHYuTZ7CJw8e50NovYNP7hHZLJapy+RSIYibq
Neks65l4eSb0uM135K/q2sMwaW2zw6iIrwFn8fFoAnArLomT1gkNkdakcrKLlfm3ZGoaVzt/7b6s
f5TO+4wjtw5dSnxgsOOCH0X+uL+yIsGqbuexgisEPlRePp0jmx6d+uaaR7ygBq4cyG1XE2bflLZs
/avE9xdpdH300oYE0rnovjHNQ32uYy1yRz4d9nK/5W45EgvbfG8rltsIy/NnDNKdnR7YkcRQ12sa
IWk5pWITxNuAf1MbPiaydSSbMppwIUGtFan3V+5flP/xJK8yHZbn1HlsR51rBW/xThK32v8Qwiry
5tMmfBKysWALGJ5t4gaEoDQV7yajtTafpTsd549bzmjIWu9BbJ5/Wz7I2oqU61fEDwJrny4Oyqdz
XSSwqzEvHRWC/k7CzC8aOzQCItc0CGqBVO3syBJulyhYES0fo8kJ1zi475r/Qqzj6ZnLrM28NGwl
K8EMpfPO2xV1k0mNrRMAVP63G5z0HAk0Uzv6zY7PSdKCgVp99Gu1bvgsDt2FQbRXkV9Tyipg4b+t
eHqs765yaZM+niEdOAsN5k2HgjMG1OMweA7uTsy4S/7ca4/aPqV3fPGt0Ys+GGjDvYlLxrTOLUr/
vJ6q0BqThgEYxEbsNdYY/mi7iETNW+8rrVd1SfD011Rg3fMY2S654PgyFv37jJsRreHUJF88k/KT
hjBGbJnVtLSSRXb/fBdvL+qIkHVM08JeycbhJoStJjKsl+B+2AO1WRCmj72MY2G1DxUwCRdqCA4G
jOZIBX7qgUBzfM4Np7wjf3800f8jpB5qLSTt/ntB3x+eh+wVmmrklExFWOrBInwn134FEX+Z+w0G
eHqvjzWUu36nI8/6lutbSJtP8vnXhjhGd9aTOfg++qEDSkSnKIN9KFHxKMbpJVw6y7FP53L2RtTp
PGKT1dZnKoY1tZCGft5PrEpqMQUtcckLl0lT4SA91IKdET+q5VYAMbDPP+KNocQLzF3lUvyfaV8L
UNo7rEXE/+J2kcFQ3xxEp+V/kn5aamzdBq0ZjTRTkYJ3hgKyjfU1oLlNDBjK71MbHEhCFigxxbsW
Wucyj8CmfcWO9p49VUZw3riX47u8ZMmwvFiekVChHvwbLFWBRD62kiHRMw8qSnNpJaN4Y2Dg0L++
dBRf00rvPqSnozWMmG6TeqoGYoDThqgEP/hW6QajJAJXrn2WHLqNRxKbZRsDXYRSiVE7pSwc3oYd
RwFSnHB1VVbZiwDprd6L73XsxZHDqY6BDtvuvCjvqiYrEYuP0ZAtFc1vp4+IVrOvHwHFXVOzsBbR
Dl82DiqUy2c3oWIm5WQTCwosR4wPgafIQwOIAhBJy2ibcKalSarBFFa7txGWwGordxgsyP+5Nf0m
siFZ45jx12Nc8odtD8/tkWkGVE9RPqd+YC5C7pGAej4YS3JSS2mEfL0Imz23JShZhE0iUwug09/y
fGuAAluJkFQy8iDfeJfqwrCqXCp3ZOV7D4qEg4jbMveVDKq9Xy/yHNnmV0mmTjjQE8YOIhAMlyG7
zmpxOWsr/UfANFjiPdtmyd9YVmhg4fhbmwiDNrqdFbTror6b0myewesayLeQPcryodjB1fFVeuxA
AFE+c/PHobDc825W+SsYRND0mkYBv/GWfDSaKqpsG/wsANzXS/Ky/+Bl8epHHpDMR3TrMKkz1WHQ
zwXwiKnSxqD9XDR7vPqvHeoDMVK+g3XJtRTCtEak/UjuuasqpH7/Q+DeYzOLsQBoh8pc0jkV/nxr
4KQG5DDvrUtgyV57hcC8RV1xXyp7a72uWHyfG9ir4W//8DC7GuP+HfLmndw9BXfbpgIFmeoKVRv+
DC3RXmCD7b0NavVSXDXvsVrQ26yQ33tYeWrZwa1xXi8RXU0uRZ/KeT+K6RVG2ude9LN0Onj3PPcA
HUQe3rWVE/klXoU21z0d11x3eqKAkSFFY0s4l3e/ccn+o3hy9nmtQ95n7YwJRjSLXj2wg+nslouP
23iV9q10tos0OfAtbqN1Me/DJyz5km5fEykFU8IIW+TcTegJCSCUCocm93c6By8+cQSPJ3BDVKPG
BU80mBXINpuBCGNkyv/agqmxnlE7r7xL4zdrSYRtTaBelwdPTIBT1s4/9Q6TJfHj1R2WnSUAWQ0K
p0BWw3QpifA5BQ4X1USb6vlJSk0Zs5xXjytXYSED9FFmPgFvlGGgHerysBuOsli+iN41qfB+bHBO
jH5S8FvJaSSmWX6XQW4MhctW6Fq5Kvh0H0H8Wdow/HYyFEnjJA49qNznujVCmz4C5lLFSKp4sqfw
GCZYlsnoVVlAhNbNkVQo6gFdnbAw8LKMXkUwqJFxFBEp/o2dg8Pq3YdnOwpiTDNGkN1Vso17JXvJ
OQBzkb+6fsCxx7PdBuJ1FvgXZfQCS0N/3gqZ53VqrGp1QbpSW+DwWf/KFPYQbqS0cxi9hrO+eS9p
A6LgZ7QjAlKyR7dXN/PqGGSi+4XKHex/5vg/SqViK57ugHnoxni7ijGIMIQ9YKuMU0rgkL1TDM8I
Klyeuqga5BWUJMVmbgc5nWNnlB4IXA/Yb3l3jkGSMTiBAnL1pSSmEXghOVNWbKhdXBm3eok2tz3Y
vXmyoQxh0yfBoe/qgvWSSErpYvzvmgcGnjijG4AffjfEdEG6KlpzLjt1klrR+GyBcg0Ri0ILJc/f
Ix51nDBCC8FvHlPOy4PHenN2BpECss4j1DQYJsXzVL+ay8X5R3nJl9xd1L8L3QDqQsA3M2CiBeqf
n2gDTDdDPOQN/QqtKwkRksXod1OlLoZO+HYcH7unlqsIsX+KRXcmC4XGKNr8EbhfyV9hzXQaZ47B
oknhTsUaH3SX4Z2QSOahEtIL9ga/5lvYE8QqBT5oV8G4xWGpPuYp2ASG0LIot1EdWCK495f7wGX9
MDVj/yj2CJ8rN0GLufZHwcLCUOYg5gvd+SJVfqFPrPuVrIuRzd4TL0Z7KbrCD4/oUDw+kz3wpPYo
eE2eR512gRvfc+wqOKMtZneRxEgaO/tbmP+hEm+CJcYI1OU0JDkeFifb4RIX4a8ZfMnFAqOSra3G
tO9aY+XOKJxwwPO8ceTqq8UEtWmBTfNWdnUD5IltClnh/EAtqGSa/4xsdNuUDCFf66hCWbxxpCRC
dnAT3fbLHApXoca85LD1KdCnwU0TSotyh8NOvYf+QDcVYDDv7LJRy9M2H97xMjx8QJM2eeG2dbe6
U7H+K6+Osa5h3UQp8H7NnmHZzDO2QvaELmDAgoap6eeja57vsrSxZOewzkp5+/T2dGDdsBM7dX1+
98mXAW9ncjsNZ8+4+vBEmIlcqf7s1bnUTFOO9q7qYsNlYMTtdli/XiZy5Ej6Wh3sHzK/niftRpmP
s0tDZRx5kMOp0+SjGod0i21F56lUY6UfpRFMaCSQB4m2rJ3P+QA0a11lolVHhmzxGkaFoXLp245A
/QHmjqHGPxmbtyDs+K9EpYXmuZq0Wjg+JTvwq3e/G02htuz8Vm/z6+hmGel+n2ZoxgMPhvliWg3W
fA3dBnXvesR1S3nUV57itfkvzTDV5014n+uUZkjy7sx6XHz3M5+Wltlg7h5Z+7/nZiZwMtqCWyWZ
ZHqTAjUdMkpH9vTjt/gvz5KQhKkf1W0FFHk++I8N2eMwfPfUxyV9urGlQK/jrRDA5eNyQpRBbaA2
QkhEBg4rhSmoxgeYhjUvsnmfG6WPhzdAGLKJu47GJyk6slluIBnjnxkVa5JjVsGwhgi3BltEFrUu
Op1ofq47QHF7Eb9rK7cMTCfYXCtUo4t1cEXkhjiAVcB1JK666F0b81ux94t7s40HF/iF4Nv6906I
xcFlIdreoY8oKTzw1HdaBMJ6sqhkcgw7q0aV/NyKF9+X/o2LYaT4+dI9ykTYwzPn6/YFfecSt1kA
3GthXAaZZumcrBzZjkfaEMThDDXWQXEybzH3e1n4BIym+dw2LmYVmH7V+eaVBo8pveBiDLuBeNSG
g8VPYnPeFae8FzSFnRf+vUC+FFh2S/bGZGU+/I6+GH1KEVzsaHHJAjzbiPdW29Uhr4fzB1pLzEn9
AlBWxBtttCnrxgG6qOnTm6vl60I0m2BZNXw+cqyxi+RPzhuk8R2kF1TAAmUPjqo60flTnmih71Wh
YDEc+DBpPZZo0Gog+gdznIj+7Mv9Nkm0udYI3W1uQSo+JBfOkbKfVptkEn4Kndse+wb7/LAJ8UYQ
y0SxH2hu0k4x5jeyz/t6P4h/ourvFnTIJhdX4++v6tR7/CZr4so3fzi+dAn4qN+2dy0suR8MRivz
3p5pgKLVs70G+3g2qTWuGbt+OF7NXsWdrkMkTbL66+vrN7o774U+DD4qGAz+HVmlE5SIwlTOFMrd
jhKCl0KFAug+vMJPJNdvHE93t4aK3SiJ5pvqXLQveOFqrKKS2qUUzK6HagVcKJHzxEHhZWMORMt4
0trf7j/wDRnZ4ughvDJHwxWRY9PF18G3NN+TQTsuPFX3ujnV5GxHWeOzvRXZ8ReHpy7UGthGk2Ek
10uSF7+1fBMiZ1PVvCP/Q43RF8D4kue7OGswPfVHL3uKOx9gOrZARUA/JUrqIHKAL2uqsWLUe12M
KQAHJ9lIVsme8HcNy70Y51JUlp31D92myOzqi++Xaui+8aV5AEnppI6dOCwsuM4SSBRCpFmGD8I7
J6SmR6uQtNfbvIbrDPl9Mv5oDhNQNPbBkLX4M3umDEn98E9sprJZleXJQAv9/5W5e0ZXAOQ7ME4b
VKab6eud38AJj+QtzHr8NYQPwZTKscE51cS+/9VsFcC/7lo/zpN7wet/2aMF7gDCFzNpkLzwrdWz
WPPVQn3+ZOmBLzzqzejeCVyUtim2XJt3a20k8mQsg61dxNE4L2o0zZNue3RKnj1854QS6EJ5RaY6
3E2XRupaMfQR4vkwHkEhOV7M2WeFWNyCNHfK0r4WwC3DrzFFn4bmAEQDU544kXMugg/bz4DT05rD
vsqWECmcc1pg1lsKIJ3qiRunGbFJaizzfwohri2RYZ34LhOH28ypXmeKrBNGnm8+cQUmRsAPVjVf
gTQscbyogV92xVmIGcL5HJs/3UZmosPOBcknK3fkZ6aDTnGPVmKjrRnmphvkB8C9g+UOej7yn1wA
SSdZ8az2JHgSDYSd8rD31IOOI88RBl2bpLbZyFmLaJ6c6CEf8ZNuDL0tQq27aM/wk/6PggPucjRX
fYDRhA3LLSyy1lWyB0UJDpQSsCxu1AYO1j3cCJEkuSBHDRctvUCxI3vVQlAx3u89fq4yqfPUjbMk
BGNgaTVeeteXg92UtJPq/S0erUkCAG++0j3OxN4ZtTBilk3golHK8c+YXkkx+V87laEs9XjV0+Jv
LKtWDX96pPjEO+1E06NvRgd2xeidNi5OZF1bJvgu9Gzi4utGidCCPe+lhwC2NU9mMDzQ27dyk24i
GmGCOQ4fyRklCWQDfdGGivVH23BfGZHkD3shMU3ppRap1iN8vVC70PlMDbN9wIAvM0ilr5tc0zSm
EkyXjck9QqRJQllcNWblNp/vcvPD2OxodOthX8phPYsEUoWG+hMrMS6ECDWTpp09hIP69qvgPn+s
4me596d5Oj3tGyxWQQ/n74bQ+dkH+4KfyrEBvJncVco8n71A+Hc2tsaygEUuIZWRbR9JrtSKSkKj
+oVj0AOJMYIUKrhyv2y2gSF5EXTIeFRntvGxgAGgBTCMCirUMOft+/6lFPHV+L1ReSZtHWpy+l5R
C/nb0YSqLRJP1AgWJVcdblmcQ166eACDn5nKvPFve13ET9kWrS21cN7vFb+0R5AqTexBOWXKXdYW
lHObMIVO9Q4wr0NZGUzEdGHvPxR1AR53TQv5dyPdQ7fWl9/ktSq6gBpKxaeolLujw5JsynRHYxEm
H8AJDvOgcpGSLQ6VPvYDP0n8CVpDhPcFsJDRbhPNdGQYO0bUyEHkCoaOsb29GI8kSJdEfC0SRHYs
hGvCMgmfMMY/yhOZN96/iNphrPs62xFURNTU2pTn4ow3+3C7cQfFam+EBrbEFJuW4rVelJM5pRtI
3zsu2py7eA3dJD1B5x+kmDuz2xBBoiOhF8a2tKXW8KqxB9PoDhYIPuo9mvUhahfhaUUTcuIa32Yw
BlJUuk0YKV6hOalh4CX5CtA9YwZua6kp743z0qkrR8lWL8zMYVpbRLaDJc4ggtBzj0CLrCJxz81B
kN10F7MZrxZAwjqqnNFEOusT+T/bVavHDi8449GLcBBRutLnr7s/H/+MJJtbZTHO41mrMvhzWRDL
kKvR+OcIjauHTqTAP2IRk96P2KM1l/n+/kM4ov/KKZDTewi96jZTohDl3v0SFccG1FuhkRgbsiUg
C+HJ93JBVa2phfP5K8MICevam5WLpvCxlRdigMJInb4iLTjpzvU6AK77qiWLth5LYHrOPzZPJFUj
WhPSl/UJbzEpYOUHQFofHanaj5TcX6/7k0TOyAI1Vbqh5oeraT1ThG+IrJk+PeqBNgV4iwm8BgU6
tK3Eqt1BIvEPGMhBnSOM0dy0+kpAke6SpB61OELofPecczv/t3Dd0F/abShwYntFV52kkTaGIuaH
+FHSLcIMAGMa1LWcAAAB02H2xOEIiJ57pGdVT+wfut1aKE2AMfB6NyrRAUVD8i1vh9RHw2nj4aii
5rFiYJZmHeUwZpOEAlNUv61BIXGUbK65o1f4xvaD6Zd6ooApFkdaKWcPIFVkmbPHnuWKLUxJ6MOh
HimHliHBk0ndGeRmzK9kxaDJcG+sAiamlYIxUvAiLG2SqxMS7ECBq9uGf93LHdLkQTLNJBWuhCkB
l1082MTjhUwD7WuU4xws7erxA8sJniQncLns8qCOagW3Umc+nAxKDwsHlVBzfYbEKxiAkAMBbXi8
c+T4yMb/QyUh6qDhm6jpGDB/gB8etLgFyGWxgtkthPgZizaOTVlWarjWF1nk0UvJDX3gVDgb80Up
KbrWuK9mmMwcSh+Xd1IPzw004PTq6UmRRNfs6FMuC08jQb86iKs27Onm4yjNEKGygXGYhjNfDmYm
hH8xRTcrA20LqEcDCvAX2NFMmCplrRonAVguvXxTTEGPGPmrwolJhK5Evm6yMb482sDfqANaNUKX
m+gpBPMa7llCbq8+2toIJ1Bdz6s79PtxDTbHLiQ8ErtG5ectY8/6ntQrn/KPax69ZXgGNVbbrUG7
uhZ2L9IjhgQwxA/ioaiXItIliX3VJVPyyYQVIf9GepjdMU1oXXaAoTdoLmPOA9VKVVw21DZIbOYi
PZa7ZvItcKsASOmHcKKNH7iGEQsiFbMrE+4hSi586m69jFDB0rs1TYBPzlETBRZzL2JlvgzByrCm
MfB38M/xBdf5F/7N07Xf+KhRgbp9kRgq4sRh/aP2xlFf1WA4lG9OMrq8zvgZF0uRQu+UK24gQmAr
4X8vG61nBmnXk6r75MtOEUvvzfAyrt6vsMRnP5eHCQdONWLP/xkAx+qtUoVfudeyflz21dzsmRPF
aIG24/SHQvsE1nbAWtWFq1MLaL64BGVZGLMBvgYKr1y6L+l916Yfc4h0ni/XQi+uEOme54fdXibn
HjaXAjgldZ4DckMch56RQp/T6w7RGRrVfgF6m6TiMkmlmvO+YSoYSdcDLL/SRvPuTqsSWsXYk3q6
4JAKINOKeksc+FNeMSFWUBsVTHsFn0JUfKJVFSqxvJlYn24h16k1zFjcF+ZoVsAcgHPRQ9rc7OOO
mDKUJ+x5Su1wksCIn4qNJpuxMMxwnWqwcbL/nSwHJwLUKs4MW5kWOqARgE7by/uhQHlkdOyWEPKs
ccDrVlJ295eATvDmSIMRo/n0mJs2bJn5kZjTuXHA3RaujzmoFAtdsPid1qt/lSzmPiMMj6ZmtZHY
sfGLiTIodFOby9yH/ev+KUvCUshMbeuT/NkUEZaoJ+vr73+83C8FoRRBqXWFjqj6ZGaje78wpfMd
8pgIrBmKdmm/ilOsah7PU4wenrsLTxIHgTQdrm4mbkD0cMIbUrBo4kopc8EHJWtifXudCK+rqzyM
YjkzSWfDIiVvur12WocQNLHcky/Os3iyK+KdAc8z71aT7iqMNQyRCON4lDa1uWS6pAtonSlS98Sc
5Df7vwj/XNWyzZsv93RXF0/N+4CO5cCgjoSVXnzACyUuM2pB9ysLL/yie8iVJcTiYnSysL0VRIJA
2pYNPZFE+Str4D+bVFWzEtnm3N4q9UYFh295guDfp5UpJVJXWWK5vyBr0YttSm76l+doZnnJQ5wP
kqiNek6qMYYygf4r+xwOs/2TGEy74sG6Y0foTsLOM4buVQ2ZhJj3I9ZDvCGX8AAWopZ8PO3EUvH1
JX1WkACmc1z4cwUb1ndnWxgTwIFtE8o3cSfkjjsiSX0PBgDFUpXN7FzYHA3WWaB12Zr9V/BIlGeG
EJfvJBG8eCtVMWdx8Np9w/p1zoMdrtIRBtPXuExUC5NBNibVGDWCX+aPXvGprj+hDigDYn+4woq+
ykCT+mDhZYba5pbGBE5PYWHNE5xPMldEfqyuEnoLXzLaYde1B0WYN/klVM22HcdsIx3leVct+A3U
ltkWbFpNRofkh3JW6XOsnCHoTs8hO4SwTV4S55qFZ9YwIugrlRJ3IcenbpkgdRZZQZk3M4HuRlx0
QzB9PTlwYZVIBDKpysy65/84ZQmkacy8d400xqCNegLRguo+puZHYJhZ/USJjIIah1kCJSXANfDR
BV0pwFdbg8FlUZE2fht0+pgiqiysu/JH9sM7nrDULh3gQuIujiXsILmI4jBFmWa5yg001wYjaECu
HflegrfJRWjEfbl6uoJyj10+jgBHu8Jnn996vSd/5fJf3lPUdv0mUF3+ZU3b3NjaiUhvQxwQ81in
xer4AA22KSQa0seTd6aa/SRUOIqgjwblDKS3RoE0VLmWhDTeyChru9FzNFezdP3AskoAcuTOGjTG
b4/HAd1bNIIJdEXGk2BiUllfipMgwtYGV37Z/6HWuog5zunjzHbQcHXjgnvroqwAlORE7bxQ8Fak
MPxr51CNdCI5lDhuIUf9fjUPQwx/5BgezRAH4XvqlbtTaxLNpgQHLGdBybZiJlnP7QoMoI5L4I/z
6WCCAb5eXgMb3vQXQv6XgTRz6wWvqXQgT2TTUtpHvDTDcxqHYap90jBLZdi+pfkYdCTskl5Bp19O
s6UidqFN0IZriUO07c6Tk0tZWxyrWTkcVoYsmi+XOYDTFFfhBbDOBleftlgePw6CfuIiIi4knGP5
ymVhdnw/V8ULFtQ9PidVkF0BhWJRR50wwktkERAR7Kd8rUG8ZYKbIlYG2bNBYzWD80Bxc+MBMz+M
LVpPyFcgGN7SqN9zdS++HmWiJ8EKfVRpFSJc1ZDNEeq3Otmb2PfLWb9d8dna/tgy0WMEwf8c//pH
LY7Vnhe2vKf69toZsEojU20bSmtUchdy1vcrSr6uebM2oE3hi7HTrci0qzCW8g7qjR4QjTwFYVpJ
pDOiAAxm7eNTuv9lQbvJFOfkSpqYjLMS0g3TDYMvZVszUcUW3O+vO/S+Wka86TDRV9qr0CapzVws
K+fquVGuLhhGNO0f5B+TA3HgG9ympusVPctX0X4A/nxo3ywuDmvbfs30UMP/PdXRTXEqGUiDTtbZ
JEtzUR2EqTeuKeO+Iglxz75yUDq30YGFflKPGzVYW1Mz61gmLdpC9UvPJTbu+yAA68U8tEXF8VWH
fXXl1Mx679isWXFbIBeibfd7kkdM5qLKJfNwr2GLGR2NZl4s+qStXieaPdCj++nkoimywqhhwLth
CDEtfmITO0VIS+KFgOt83V0UBuy0APVJyfK83d3lEBgxT4kHLZITgy4Xa1iQoF9Lb92u3TDaZuKP
aNgi5DZ1RAwYglyg+1/Gs+l0GihBqkMPbcxJVNN5YykQptiFvhBoE7JxeZQmISk/HBBnul6u+er0
1ChGkoB/1A4M18PDSeuGE6dC/JMzSAqPV1M8fkQvS9C5lpP0WcwLAYXykfYazw0Y2+hviocvJPvm
i349OnKLGlzuFPj/OmuLQxJ3hH49IL4oaEKCNyIqMscdcjfU/UAB1rx7kdGjbSPEQQxBgjZOOo+s
5YGUYv4W0ENLwQiHNTsoor5eHJfjVoGduR+d/ImDT3HEchwr0s38CJDEbKCJIG2cMGaJ41BNTt2B
3j48NhSnp1Lqr553s8t97RofBN5x85PY49aGjxDeNSCyd0PG18p83ENfomJ2C5sFgvIYLefLzxs/
dRlcWgPhqA8ilighKkgBklkJVHUdD8fQa1UDT62CNEmT/+src38UQ60vWT6kFxoxa7B/2U6xCDgZ
ggnjFtuH8TZ19C/76/HaWqvhX7OHCBM12qSOz1egQ2DPgD15j+VWXVT9GqSPAubbWEpXv/9dDN75
LlR87S9umIaEMlHIc3pwB2WwMo2Ur0uKCpW47zRoTp8mcZ9WLB+PuWB5o5tTqqAPD0gOp67MX4JM
2ymK2M8Kn9BIoOUcU2qggLX+pSe0D4KNzs2/Igpr0Y2NkLklrL6UWEukM2nHogDNjAmFJWKW9hQu
YWszKgXr5wozo8lf8Sy0rIGhVO4mxY14Hx2NMUhiFFdR8zLYMvczgP505Vxqg3JxPrmUMqgml3AA
za8pi/FY1Vyf3pKnEEbYPRpavQHNswtI55u0eWc8rdybp2x16117gyEAVI4o5R6B+eo6mipsiEqp
J1tDDZsSpbMxUV5HfKL9f7yXxUWfIK3v7e3qbn35RRZubByXs8344vD9XW4+0fNZLFA3hX4hLgSG
4Ylt+fv0mu6saEYouO0ivt3vAHa9p7zmynHNftJYRvouEZ2HTkchzom6pWIm0BUWqUFx2e0UPgpj
chYqfVMj3Zd52oDy22VY8uwhVJt8Tw0RN0JJoj1yYQuShknOvouYn12xZFSSrdieAihbZbihFKAL
pBhKCZxXa3xYyUkkp5bL62Xs53mA8aFkzX/SdmZNe1geHYrqqdoINESRroeaJX2FTdTnZ1Zr5GR3
J8GrBJ0tEF8UOE4bITPJ8e2xDli1MQAK3lLphE5+phgpQn6m93P8ZVJIK9yVEEZsXCMsiNfoiqYj
1v8pFPo4MD1Tpiv0Cwsqkc7ks2RshooljHK7lO9WSZJim/CXx3P15EBQirTAvBn9mtsjjwbgTOLd
2o7qxnXoqDgq1Oaxfv6er9Itp0uzsu92SWTpdyFME1qZxELVtsrWm+K7FzS4/BtkW/5jKtpKTl0G
tWrrd1SjDY0rMEFJ/JSowdWJXyo/ghHroW80GhsUW9Pc06TOumtU28HiP25e3VDIJtROkqusntn6
pl6cX67Zn4nTdivSjopQUG4z+uehZmEoDc0Vduc/YYhd1KQ4ePcX8ZzdtXGxPuC6Vni73jPkH0PV
oMKkSUSRFuDK0LrhlvCtp+0f8UuWXBECL46suZSJJhRAAsFHmfsTd6aiqqoO6XMk+aMhoMAXiIcX
oxYUBMbFIAxG1Jg3ECP+gTMeKBS+3K+TLfs4WGzjhlocDaAj0AzzJQ/ngxmG+J167/OJwPBp9P9u
OXJ9YOvSw1gqNhjb6FASITsi9CckY4qfJ1uEhExze6ECbdK+Szxe5/ZdZZesbDuuVVNxctnARRQ7
6LyfSEE8zvLnW/qDTnV0SOTPeaTyTuLJit04FWdSS0QxBozB1b44QKouugTRjtJ7EQrkQ3MSJd+M
Ib0cc2hlGIrwH4oWV15Na4WtPzeDNBQAJIlhKnCZxtrK+4sehGLrAbtjqCWTOIsu9hp8OT4mZiFq
smTErjKDw2dA2uTf6mn/ahW8WIBlbxCPd4BrlS5ltB28ksV4Os6bW3sAn485vra9lr0pEz0Ey3Mu
hECUfaKcINiIxC1VXEhbgAw0V1SDsK3cxQR49EYqszkOE3f0fTrYfM3F2OJlG42Bx63m5bOzp8IV
bL2YkdjCJpPshEKkreRBK4n/elSJzuVmFJZ8C+Xu0OQZWiIpvnYyGXBF7kGiew3CHoduRgRjDvCZ
l0BQF6MZJmGdhKAYK7KO5QwmE8stsqnOjsefKuYWUx+UAHQLjBgB4BCswWIusYiYBW/9mRvvFpxj
maM9dFyrRX5ucpXyfn4ymB7stN2+szkspOJ603UXZ4JD6mCmDpX+ae/q+8oydzwM+W4NQN47B3dt
N+ncY1NfdEs6UGqprF5bZvCz/zpX5lkJX7t9KUfWOOppRYs4fvCNa7v32tSchQSt/KT4IUW+kuUo
7YwlTqXq6BflUHhls+fA5xJKsqzm6PZ2xYIbuquF2eHVe3KyVjgqO3EM1dJ9+6vqnjNDBSWI1WBI
KsJogZ1lJkFfTgmCWiVmJlwhrE5YR4AGTCkQyaQ7LJr7It2ch9UHEr2X9xn2M0cHcthsRVtr48Xh
7xtYd6rDoDlJRoTYADJojr1rR45tSeiweGfepUnhLTVnUF0OTnVKKycXvuY98P8JbkKbDICXK27P
Mi8rnk1aeN7YVQ8ruUBiiC5IyWxUussBgAy0wYkQ26ap802ZLF5eN8HS1msFwkhgPNVJYeeiy3+4
5l5hTwNRmCIf4rz/2XDo34SdN9xIsGcoirvEV9eeYjaZTjb/FxRElX31BjPOiH2nE6JQymANqvbn
ZP/hVb/6gX70TNQV02+6jvSezZa/RcwiblNAysubSG1alh0VGNaNA7FA7YHiCPPbovVZH9U9hOdH
IndR2/LtgPiNRGN0M/r384XElRbYidC8dLC2tGsz2Q7r4n4ia+QNgTwbB2Ll21uw+5gtsQ8qWYrB
rcZDHAVCv6v5SjzGEyklGjSoewv5n1T2pr0UqSNZC9MdzOGPE/HjGmEEaqcgsReqE036H7V2MLb5
YjJiubOx7Y1X1gYJmnJMWVBJCscSLukiI4AFUwicyCLN2WxgjSjBYOPxZWbOL2ja9/RqfRTvopiC
WO1lUwD36Otg3a+No5pOVfoiO6gfb7r/Cu67FY1KdNQIPKHS2M2ohvZuVfZobvjUbKqoT0ON3MBy
gmg4R9CkIXeaPPO48xJkEvJGd1AwO/WRg1hGpQQwbDGQJ2FyUjkrQpBMPSiO6JAMn9a1cIFedwtU
hftDc6ifuWy+azecyKAXK8C00TK1MfKDY9eIHmerqzoo99bilEtAspmqtaIubjTZLPgmXfoLeKKS
qI7A9p8xmdyVuwflK8QWlwb2hNnQMPCV5kI1X1E176Ql8iSvKWrdwgwIejOiNGfpPzx56RTNi8lD
OkVS7pUY6x29WWPZT/QtvWkOQbhrpF4Gxq7/ZkFiesCIgNQbJN+/lN5Fk+N3MQ/9V81UeX1YIaCb
M/14H/C0h26u/22rxMxUSLnC3RD52S3x+4XG95h3q+EPXpZBTXhLnyHwjeWvICg8oUoKALFsFA0v
KfM2H4G5DbWQL2disFkEZ2+sZio4BHopd0AzPm1qDtzjyGQv8q3YQw7xqE+FwzIgnatCcjpPBMfn
VVZabrWFcD7UWwCP9w9z4fUfWxqHA0ZT75Hrwf5A4HoEt4LxHCDay7N+vqDDkqNNGupHmSFSCCqa
n1uF6KMiFGAL0m3FuDX7FAsEFBuSth2lp4UP1W9mqbl3Yue3cS+8qnkb/J19TNrhbk9LDC4Uo1/K
GA37TX8UBtcZEjKDkZpfDTh53oofPzLdbsAMmBrJfqTdTeosTQLLfLlCW7RDgiEByEu3SzMW9lOv
+mk0hRefbtfHS1fxwM+L0eiydW9Q8KbizNhhuB/Bjn1trg5lV9cKR4HAxkmHn+p7d1tln3+5b5cW
GWrpDiyX3skUmr/RYR2iH/4GRtybyrLGXdwUF5qfJFbDN+YPALb1yKgSvOFnFLTGJrlkEffwuYEW
iWHl8oTKNaf47BOaHhqx6Zi7Sjt5eTeBDk6TgzYsfy8p+plC9qfZBfitOVHZ4HhuFVYt8/o8HLr2
GhWVagnkMj3kl9kPrX70Au6Fmbc9rPfVyPFQhB6xp7A/wkthLp23+DryPvgP2UTF3cOAV8Ssj0SR
vusdiWJ+SOKoRXwQ97FSGxbKlx22Fby+auTZvKKhOxgNtzLhOVABMKcvKNxG90IgOvpkNB6xO8jU
xcY0w0huLCXZxvFbX8BBAegvAr2fgrFsQ1oZjr2OFL+qN009HZSobn/UyfTJaq2slbBrfCnqJ0ax
gBAg3jcrYdoLrhio7enLws2rc2PiwO0idf19UKRddp8yk+lIqOqABnHt4T0/+TB3Atsdh6knrGuL
hKR2Rf+7iYuR2UkiEW75Z1yct7cjL/qd+T6UOSgo4MrwkeTYveX2OKaYSDD9teTZv3k6YGdTqlwy
YQRqVS8FsjlG4vFeUxcY2aoM+DsNzbUwdPs4bGJ9tzJcxJuz+9Pj76L26l9DFazJ0bIQlJHTH2tm
rnDxjlFVVtw5ohkbljxO8DS+jpwYGv7tZpJ9jKlrY8ONytGrd2GeAZhPlkZvbGjzNC/AFYbn9TfI
JF7/a7MGHfuMxYSSNBJlRukrgpqGWpaa42k8zFLWVUec++XxjlFtfYtUCPMkCWX918S/wC0SazhV
NMs7YjigcHlVibs46+yBsnvGhgMzm8yFBZZ2HZ0aIgIwBolUQ6c/x45BkYxb20+fzICLCcvi3az/
n7TD7aiwUvRYjoEkgUBIIZD/x7uA2i7cmq7NY9KFmqHFht/dP/nsHo9sCzOmugzv8MiV/0Etv1Ij
u/yxkvtdKtyvWVaHoj9H76QYTlYB7g4LHmwqnpeb03wCPru9xkksSHVo+IQAwL4xP/G3UxhYy3Ww
lh8KxHWPf8m30gVGTgPVHOuNwreJ6vYWYgQwTqYVjXosMNcWKb07myI3vAVwK+q+Idd5V0tF/0F1
Rl1emR6n6XjpL5zKlAkrd59SI83kcWZIslqJGbke0QM5tjfXn+kXG5Kj+cMloFrja3YODZ+LnC9R
1/6Bqyvd1EFdonIlEp8uSVN3YL6xhuWKi97QHCspYcG9zD485ardRW0oC8KEdqXvNbjfD/EZdaiu
P7fe11nHYDD6eFIuKzhxtJZzSRWKtwlfMbOtT1zfV+XxUMYg8IrlobfyLL57kqG43kEhCRaDB6mE
Su6B9VUq9NAwiSslX17qRHG6UsmCJRXjU6pBnuCrJg9u3BuRsUrhz8F2Xp1KD1JdCwckHFOnKjbB
JwRm20k1YGlu/U0+SWn331se6HXfmFaM0AnxpGz0CWgIhFpNweMkavw43AQmX7bZoOU49nO4KyTR
pP/+kFX02K/dpwZUcP5FHv6K5K4VuzYEwkdbNORlN/0CKAp+XR2PmzOOlIK1sD5dq87gjcBMWAXl
QJ/JLcdZ4R7ek3EX7Y3yzR4fBP8ZVNJB2UTMP+0nRsfURYgM8+hDyXbUe2cQZWnXfNUmKf1akKh+
nj5+vOphTz4zIrD2ARX8Uw/L3Kwjni+iiODGcW1/Dd+D+50xZsY2M1RDZgWs3ZcrEWLGwZlGTwyv
s54w/IfHmMJu7HgbHSq9ED8yeF8t2xauolN8wN+V0mlDlpzSRMy9+y9Tt+XjkpB0PT+BiyByy3Zo
ebrSkYFdOj9WTVOSykgAAWwbix+6Qm6bxdPtbGgcfvd+gXWdWLYT9evGsiatPWEX1IY5EwVIoHCU
ewGYNkqFt63UhiIs14o1JAbGOAhZy/vVl3i/XtyciiOyvGjV7oLMw/bbGYR8d7AvuHzdCYAM8lTa
wwUBk7AMWTivTHxPG97FsjYzgr4eGTowqWWFaHHZjSctaDn6H8sfbKWwkGmTdSNEB2ztxzH8MnU8
IqbP93ZuePr5qaDY9G8YmBl3nVqmAldUyrzWXfxlJAdbNa4FFYIa2uBlq7bn4RzjCkOgId0CdlOr
nbKRIraqRfsyLsIU178LsEAmHgzu9xS4LYgR9yEeBbyQGzBxqAHWKxslIxq6VQ1GWXU4N9VIcV/R
AiV1weJNfOWMbwK/TIC4mQ0OwY2xVjTM013jImwcCTYoS3dELrb0bXJTzofhAzBADQQ0WCMj+vHk
2NJkqaZ6DGM6Jqg7ashuaqKAPYgRpCGM/hDpFRF9yPC1Os055MV0fInpX8QmlktpXGrLnpNj3DGz
IhDqSKDQRXClDcoimkVZheyrbQH3prEL1NeMqno9aa8uXTL3SR6+0gcIjqoKRN04/Qf0Ii62N9a2
qPI8UL0CppmOKv3ucW3lBBrvJ9AfyS6uIAM5z0FtmkvDs6G7oJ5tVBOF69ULhPeeFblrRtc2zNB+
SK5E5K4zF0naPMFOLySI8RdtkKiPaXzayF1Ryy5chNXywBufyyjjG6AbkeEbKNd4vyGg6HwaziB7
iCYhvurZct1Jpj9l3ch7S2sv7PfqtbBSafeSpfhwtY2ke9o5E40X19sUujNOONqO5V2smbIfgZcX
KFzRC3i6yPkrpS2Sp37Z2mE2CJqK1btmIbxHB+JJnJQ8GPKCWZRrZtHQw9GiVDSL0/aIivaXgtZa
TfXz5/oJ6Wyrg/TD6uDiPcgR5QLSkIiE0WO33BBcdu6U4N/MHpuRYL0xNAR4sOJSzONyXdeNJ6Eo
N3ZTS3QO/lHcGk3/G4IeyGimjJfdZQOAj9zx8zlgXod40paK1OetY5cnRYxgQovPYsE/6/TYoZag
QS5co52Dacq3I8ACZPnLoCCNsVEheKXsWXQvMZjzE8hm3TafbZyOC99e0/ZIwN5HptmoM4Nf9MEt
9+YoLa/wdV7uvtKOPco1VBLYezWHnVRM9ZeLSyemfFwWRZWuWW12Kjl9eLQR0fh5sZ6s3I6woRpx
TMqK0Bw6jAduUzgYtjZpKYB/4p6qJ/4hgIB1vkgb4KyBYBGabdWlzCYLpJTp1hByui5NFgmJFl45
AdjBdyCLCRX/DykdTfn7jorPyOPCrm7eSS6OkEMcJOXouPKzYdX9RDwY2zlMmPoXwPPsUMu34i3d
yjTXEPN8ZBHGee3N6d7Ac8IuUPSdlCGDVEac7ZOpuTK9wzmUB634AaLf0pZCULO/2ffRwitcqdGM
C2bUHgp3lYIFobd2LDNSeV9Ns6VG3xq8/0c3PDHNnDRDBV4ym9tMloJ5DsNulH1hBJnnVigqfzrg
EP3Yg+/JI10oOb4OsC8rPIN1aam/tQtCzG8lIVkYohIWs4yktefK2Xso1jyiCqW/VGInmBQBfv9r
vXE75iDdM31TAJFG8h4hLG/cJHkMbm+ePuHYUD31MIXpdq1u+kVbhcJ03DBkwV++SmJQlDTeDrl0
M7baI/RxfWcqFt4C/AYtu2Zf2rkHJzBEcSFfOw0JtzW6x5CvWqKzIxFZp229JFv7FvvzpSb5cjn5
R/vXBwJESXS0KB4cMCz/j95EsHjTXh3e2Vr2CJmHBqWT9bzCMC3+m1fpdnqyyM72NS5yhYEHacJ2
smGCuY7DtmWuK9tsVv5kcfS+9jyo7KOc0vXAfji7ORNX+2gRx1f7jq4uSxxpuVdUZYDGPVa1sK78
WVCrZBKV2oJnWnzCdbxhEw5usE2njj0BCD1Rc73p/XYTm3L9XyCKhk7+hnPUa8aclxpMZ7oTcUVO
ENxCCZDNr9Z+yY4kZUyPGNrtWVHGkMtOmotg+81tvHrW8NjWuoJiQXiShmP0kX+0notuATIPo7D2
fS8P3Eomj01UTG3mXMDK9deBdveQUqNZ90aHphjmh0KX/K5H+UkPZ7so5MRrbDDc+MRwb63uUjWG
xBhTSHF7cUyjXPAIWL6dP7XigSyDSmuvBHOyTl2m3sC6aa/cTFDVdTSa54/8G+ZHlBasazHELTEH
LiibgI03jQLtr+SwOoIa6QGy2uBCNVd5BHdgvR/XcehOYfM9o/bKjMVMKF/eD2mDV4VAj/Q51dMU
PUiA7C9yoLg4rx1VBTDFVwV7HOOUltrlfUvNAKgaVvPqaTRPKk3H4/KHoVizSEOv2Cpvc9/y0y53
H2RXKNHzwszj3TmolSs4OyqbiD8O7rE9MNu66uudrtmp0et6o6n4nHFIbjCg78NPkd81NYoWoWIW
e/VuB2Ivh6b6Kxa3M+M8bMN9ZdMtPxHLbCJkWxHMVV9cuB/2sCird2RTt9IwRekwdxJEMD/XG8+0
Gmij/SIdNJzgoA6mL2gZm2GHVrjEjFX3uPR9UitwB1siX2yXfB3RciD/PyQkoyuZN71Freop0BnH
ckNEQZ4H5yPbn6jQvaLNHtxK4/Ym6ESRWwZK73P6W0pjAyKN/VUpkdzs2YCtdMA67+BC9aE8Wq9x
YvB/WRV1nh9RTobNZ+Wetnsno7vIAVN3S3B73Qu8Krc7wIr7t0chirkKcrFjN0SxbJ2HtOO2Pvni
AmApbv0E+4lc7GpS+G39Sul9AyQZzQInDw1wJ+jXTB9EGHjRyLCCGox3p9+Y4SxHaRNIEC38g8jO
px0L+/eEtO0x0JRaYYW3/60Wt1ybrnyq+KqLpDtYO4FaY2BCKNBELw8Sfqz8Xy8ZSqf2ASrnkElI
efgRzYjGATjcsYdBOljI5SPjbq5UsPzpz/Khb5DSik2Sk53vBvSMGryCFqq+pbH/7okQgrCMmYX+
4Wb+7PeUOaM7bL4OlrkdmYuekVSlgOdqFkIsVGxL/4uIVYVy2I5fBdvHCH4zwrhMllS0pzKs/+Fl
xBp68hTkZ0UvAUM3m+XOyYZNqsF2t1ufwdW1H408YbDlUmRe9QR4IIvyLVc7u6nF+Z8kjKyMiqNP
OBHMZa1uYWXvVtLcOcrKee0CmNk8D/Twnq1KaVX7JJwe61zdDrLSfmqkwFVgq5eGXh4kG2Z3szYT
dzagAoJVrOpAvyBn4fZhNEXfUMKzU+Ia3liEmaV/D15RH1Qt9d260PfVetmWDHmQXN6SO8LZ90f8
byCmPN7nKi2313AY75mozUQU94wyL98haXnz/fAjj8ntSnm2GhqrzAep/MjY2luV1yZPwNW9iNx3
Y1km1dVAzlewgAGanHbKUShb2d5D2Dq2pDelurpeqkpTSh0UnMSL49uVOQHc9T4pv+7cjCNArpzb
gNy4FLJsC+KEyB70CCsvaIZwrhDRg+QI+dpoq7eW9GQeZAyXVXgWFZknwgO2OZPcB8TPQ6GMLgPr
HNgfkL/3/Qo42HnTQb/vZcfle6RMtUWLOfinJxK9Sx89xw+7gpT9Bb0NLKubQEzZwN+THhKJL7tx
tFqeoTMnRb9YglR1an9JnKbB9NvwKEROcbL1Qw6TtACSILsq6crMmrWFRqexQ9enXa5r71vwBiit
p5yO7D24hlcHO4nUtmlh9Xd8TZMwLvAcwI4JLXlsXH4D2UWTMMHnaz2+RSkzraIh2kP5i4LnuVjR
TuS0qMuXRmad5zuqiAV58+zCelc+d49JF1SF3tvKcJgjWV7WJsVCKA7JmsrVEtduQHEyQYrtja/u
3MPktbbFfzKtxTmrq67VT3/Nz4c6HEhw6zPnAiVm/8uKKQYkA5WR1NqbL2ZQ+ogBIycXTpTv2wW4
c1wcxlWIYqRLcXhtv+wwqpmxghLh6Hjnea8QthW6XZ5J2Sv2i+FUDmfSwZBXMBWUIofEboEQLfkK
W5Aj6oOrXC/jK1xwXKJ/ACMbrUSue6l9Ww5njliilyhwpyKnLYhQJfaJ2G1zatR54ahf5G71xviC
SOe9Gcd8eN5TXgMH08ZwVlkCKGRsjS0D2YnJh3+x8lZ3m20Dm8LbLa+aHsV79C3BbvuIKy/2XxWl
/Btfl3MofSHYXaQ1+DzQyNVscOXo9i39tx9F2gQbZqse94PQk1zxidxLnlk/OM+hOAFbg9pW8Ra6
iHNXLSOQTTYLc6HWHNkTuG/JHvuow2RfCwPgXy0Wfc+88rO7Bt01YCl6fLNCoROPTSDDMoR84CZ6
o/ura7r40Y9LYsBpnmyPNaHBXcqr4dUzW6gLnEVn2Vg/glTgIAxYrjneySFziXHFy0Wep2UNj8Qj
tI6pjINVHIwZL/4G/YIvQQ70fXKz6ZIwz2tLtz9rx+l/q89Jzj+pjUDQeTscqUOdzgF6Lyx8+gLz
ZJOmXkHE88Glm89qWx9Ax5C5jnzE+kFZLfw1ZTa1QpoKbwRoMq7aAJOxdqnimfPrPo4w4BfQY7mB
6973MADw3c7u7mduAFO4EhthLLJEj8IC0+8s1Pu3eOFb8KA196fuRgxuOENdlry2ZqMwVBslqsWy
uCFcE38reLlebURDk5zx/NqPfivd9HTJdsOV66dnEMcrv+eLe6W8aIoTEKNyVdOej73Iedc53E3G
8eDQ5DOfgm72UlRVvUgdII1CYrDUA+Jqq2JwRDeviRaUvBL2fWVyuQX3tnvNhSmlRYoX+7d6ABaN
kGyGGZqnbmqt4kyUs1CC/SiYbivDXNB5q2acfdm64JRXSntDShFfnk9IFNlZxtMZjLuPxGyFlits
8ZRyoRjQD87v57Ubf9dE+0XRrsFVbgQQM/03L3+J1G9Y2UCywEvYkbiWx1zET92zcgEM5q9PAOi+
FbF2a98/EoyDJ0kLe4xd/GR5+tMb5QSVUGhed+77A2PdAK5jL1GSVK18tBh3fyn5Z5OBXdsHSZxE
ZTor7e7g+/MEy73l2J35Kn0cVljfZ8iiRZkPtq13Nh4MQKPJ5yMj/i0v4auw0fPahWQgpqBb+Scz
5EG6iEPwQeOHdEDWHO9KUb+/X7F79KEW3yKfuhtMWH9lx/Yz4P5+k5vU4B2en/I22+/psYR7dVca
56/qrqJRmqBwa9bhq1/uf2YXi4OzVsuuncHex20koS3+HQl71KNO3aXi9XC/GthPZcw/iXhKKOBj
ITnNnkXKdEdfcip6qf8SjUF6FWR5KKIodpDGvPZ7s+roDPV4pjlEXql7z9Jf9+z+Ywo//4kLkd+e
sosE9fsWFUF1Eg0Tmz1WIHgo0VuEQXUMat5b65kZEeWCDyCEd/Yxgs90MR9wVQtscNXMWp7CZDlF
lhiOskZ6VNUJRPzw9aveduhDeLPmdO0feYh7vOHA4HNw3OHzjOFl4mHFfrXleJod/e4hCSJ0Ii7k
ajqwfBiRCGv+Jdn/I4AWpX4jfAZc2ZpiOoa7IIdJSFpnJrdWes20F16qV2k8NQ/Lj0kCG5AnX34k
JMjw6BAeE5ViwpNfZEhPOn365ilsIkcqkFEONXVfQHBEf+UpMpiEtZBeBf8yehvOKuwI1cK5CC0l
TDW6TZAst0KvoDkdlQRTr+uIDZpC5OnqAPCzYhrV9iySHlFhzyXfDMtoxKleVtgaBcgexHmlSkBb
IA2B0bi4azi4zREnprpveGhJ7zDqjJfrZe0fklVVxuDj+CVxporHNFVL2z6iebP0/DUlH/h4EO1S
JT5jELCP8g+9sSVKbYp+4Ml0f9UPcPgkP18rkZ9l8/L6KxrZ8pt9zjdSj8ryzGu+J8GsadIb3JwU
o1ZeV5z9b0QTeRkOGwRCX54VbavmFKcyhkOVfNuyGM9y9OTrQEqYGjD33+wxPzHHzX3xy5o2ZmP1
vEpru2yDAa7Puth6kfW5dtmpvbUk+ZxvB7Ua+LH66pcZvbf4uRd/XMuqGTMAClnozNwL1s25Jh/7
1XuuPaCEEDdiAEcLXRpCVW1kw3t5+HZTalzpMQWnH2cbxuf7YTIJ3Y/tkxqKEajVo8CofC76EMuM
BwJHLF0i2zTpCUigLK2yEpDnxFNhtuEquxoT0cmg577WcnlJXfDUH819L+1zfwAqKCVPHbKIhAlF
OIPDKwUATZJpVfzjbwjwyVLya0P0WWiANAf2G2OSjXy8bbqVC2bpQf6yGyzmbXgZlXCVy08Di2vy
Hzyy9hqn7xVZ5ReA0ILqnQrEBmFdMtox6xjBep7Yw++A36amFYmc7wTGCvAvxwiheLRCja427D7s
cePW8BWdHonk6u5+8SmWkKBvDHBi3Y2tUET5oTopwrJ6zvHabqfV36EsSs1IeyWE9ngvNGaUbMPV
HJiuJ5M4xzD9YkVeuBtTRH3W+TunhqpjgUVu2iHRqPW6w6P3YBUjKjRrTUSvyWu/sSbcFZwLUz2A
WWj7Ap3P0TZ+m+qlyT8g/zr/r4sdXHetaPvCc7+uokEYoqJi8eocigtVq/QEsHD1DRZvr+QeZ5FA
Do+GG1ebQM5pGwnG75unVLqsG3rhFwrSAofqqkx6hxaQDGhUnmR+3KnPNl8FqAusZNxO4xYbpaNw
iToeV7rH5+ynZu7Lzom5JqsqONdofkeegHlXIyjQE+tSSxHHOOpraRUO2PJqx2VLq2ZsDAkKfg/P
L9Qwv5SHhfVrk4v38sPZSM0HERVLLKzru4Mkbv6HplfB1GDx4kH6VTKsH0aeC8tkG+Q+JLjTJzOd
K5JE/XRDcfTGSGjwsLAbwRUKeTWUs71RL3u9l8xNwQteESt8Zp1C72m+g5AjGoOOQCHVcynmpPC7
x4Vlb72RMMaOYTTi7++oasMAWWG5f0TwOg03vx2O2sXfTaxAHi7z+5lna9YosSFPudRvd8uvfj/z
MTbCEkTpGkwH65RmHczqQZcu8mBQcB5XpESIBVJlz9vV79onpyNuKRKp44uz3HTv3jxtVoc4m4om
XHBgHfoO2RYtqcDctuA7G8wGD56JIhTphm+w0u9UkLl9EshK/El1aNDaDffmbr7sKr2QLcd+xbjC
0kN5SttaWy64qJHueAzSe+WvcZkWvQUlrSMbZIoo3nbEt08CSquFizITjyZ04a9AO1dhu9JyK3ow
a9eUDXh+yoxDOVU92iquFJaAG28JN0ezRtDT2uahYSMeE1O3Mi5CI6KZxl6rGTR6HNFhBOKFJyTO
i8+UMbsv1wLtt7dLc/D2mkDPJJTL/ndJiEhcpmbSXlZ71MK31VlokkO1ULLnSiWYXoOUOqPcP9wM
PaYBIzEDGXVgNmZrJwsHXMZ/V8toGfCZXUBYzCT6I1OH6roP+WMvjm2TiAb3Hyw5uX5cCFQHB5lz
KRDTSlWFjWWCC5pDNDEUpPcGStIHcajdNrI3L44SMbPgfS0zODE9FFjKEywvQ19cMJgexBEAVGyT
nQtBrVIaywpyBImvde1GrJSzeIZ6Nj2b/Mp6OAyAfHRzhfKw5eUDyO3H5uKoZhuPnL+CaZA9iziO
nZX6ywVBS8TcqUkYq7Yb0Yy+/foUqUlEaZpKHoT01O/lQtHNXRgCHWxD0Ub/MzsZlgfryJYzJd6a
a0rQ2XcFgFjsiKD+MSP3WwSXH9fliczU6uvT+qN8gua3P4g9dIN/Pj/1jBpcXN4vdt9uvNO8OYsw
PFn9ThNspbVWRW0K7vboMZp4UWh19rhzT1ZbB2MGMp3IwtQ2AnsJWqKXB3ZhWaoTl/D/O7SibnR6
CLHD6mcGNB2r6Fnrh2HRXQewzmrApcOzx7ule1XWshBQgh36IqMPJb438z/W/6eyOe3vArAWCc2y
De1u7sc7uH4zj6ndpGjXJ3LPeFi2wMxfmCVbBeVPFCc3huvhjqeBC3sKE6YJ9JJ5q89pw9NMTuKH
wTlhyQeIW7AVsAeSuAfI5Sm8mClpvhzHUYNnE73XMHlKMKtgjZs4J8Vi116fyzoZaKkylhmSWgkd
/30o5+wMtVdMHfYFZZSrpindhxBKwvQJSBQR8yASScYGdbTcOS9mDLnrDKv9xOvkuhdJT0F9Axg9
lzpzBp2D67suFt70RlwDx9xvaR6qrgmCI5O53O/Awa0eU+EaBZpLawbhrQMj0u/C8X3VZUU1JWqZ
pp1a3oc76JjO/mq0T+RmHGzb7niXoia5iTDfG5YgSmzMVA18bj0H95iSLVc0EOS/REkDNIMHIUJJ
2EkaW4GiUUAx/Grd5r3lFUL+jIe+UuYRnapVXJJEphH70/WLKABjwhO+d32ydgMk1Duh0z69pKwH
HMDvUbB/L4038mXDYfDLUsTXmsBpvEeJADKvkVYEz6FQA3aEmAwHzff8deWyY1cRHiWGURIFDjlz
coToYWRPbGSqygJyAjFL3QnZgxJ9jIDFQ2Y6YIUhiJwUl5UGxZJlJtxNVvV2GIslrete+CA7RUcz
/aiSMasRq0EPUzZO33o1RfBDtZZj5mEiq1+Ayqhx2UgVdiuhKdYGJUwQ3eQCasl2OfItwDpWLXFZ
/NJjOkqHu3gT/PV471IX5XQ3Tgd8uS9W+Qno8XdfD3cXQtQPF+jGZfz6nGO2Opc1wHvz+OwdIqgD
87xy9vey7vCKZB3E6AAP8GMACFM8UDKb1SO6bm+o2gheG6CeO2iab+V+9dDAHKjalrBEkSWThqhs
sUNIDQfzTA8KVGn0ivoXzvY3kUihxs2vcWW7w8vV0k1OZEyNC3X+mwOhEK6ZiO61JytvvF5cuo45
AvcaTdWjZSUewjw3a7T8XB4S2liGz+7Ly4xATfaSBtFtm0Qr89nZczLLbjw2FV9OAb7DrdJxoI6N
z3t2CS/n0z/vyQy6HprQmjDlqnfSpB/U2fSNF9jryKGuPsKFkO6QxZZLoV26duDbo2mQ9TxA2SiT
NCjUxbfowdDMNAvBWPP5rFZ3UOj/nG2mQUaOT4Q7d0IexPvC/59VUavlq2igLzFpke+dPN76tKMf
WXpLllYa1bPESY3eUL02VzCecNAKsFnVbXnREYTdB70hwBHSy7cm8wDgzmwyZjwwKt/3c/5NRTAd
4Oj1O24TOvs4mLS0VzW+s6t0uzFR898mYjUquSVwgNilc9h+Yv1C3GOi7OSlPhcFmgT/4gUomeyQ
hnQ1P+LjJAPFe8SDP1J0lb0qMLRmhoyp28pBj/qFarIu/TOthxlQ6RSfVBm+Q1yavgnzleSgR+I2
67FvGAQtg5oGoXMbd8h/iBh5xd3DDgzPDblAg0XlMFUmlEskAfWgv38Ldrb2hL/fV5lXSkmNguO4
2HdcCwt8uQlvEv0B/zcD8Vl0GtiApH/V3dMevmhhG/qnRN0P44Obxmy9OgrS1EJ/G1yb2zqTzuwG
zCjTu/Lv2I2dljvTEwqrlA7gM7cwszraeclvUxbxNOPROzXeitlCjBOZlOZtibrlhRd6rXd7/2rT
r0SLqcb0oPLOCQXQrhXJbrbXrx4xOnfPxPmuUMgzXRb9YNC8rClVhlyNK7A3CxzOPgDZ//dYl9nB
yWUlkG/HmTZJd7y36rgl9qromk6zCuU30SuSpC2WD3tMkVAIKdzdwT1EmQbis9PhaLIitmuA4+EL
9/rkBR4ktlpQ/UzLlq7HRjaC+2ldSpm5hVSTH7eR1LqmK3u38caq90NOwGnF7T1Cn3lIlH3U5Ile
nzYLR9CO21YgDU8jiwzV5TDJyVB9Y3938+RVzE82+MmxTnMxc80J6FqwFJYat4SqWrn/ml9Zb9jM
6SEMReDkaSaB+UzZgcUYzc6luqesra7DFdAggAXvbE99gRIx1t2RajI7n1DdYRnJtzy6Itspi0+E
8wLG19finvu4r62WmzlqFbSRBEbd9zdnQuBUhH/nDOxAFJAD4glpSh9WbOhN86lrcYy3LxjJZ5wE
edYfaIZ6GlRUilBNs1eCg8lF/bpDJk9iGnbqE0P3yJASjGMO7av0+AdMIlaaUiuNjONhifNSbv/d
edsMCfLC2lGBv6SmdlLU5TXgo+C0nTrTw8h3jlcMwMncv8uOED/OU5ChqtQ4lWCGndjsNwbi+ZW2
cKg1T54fo8aaCcJzBC/5EOdXPP23SwLAw/D3HZuV6ucxlYwsSrKYM2ba1OnLTHFcr2fGJm2nLpn6
X/CzLuxgzxhqGvoBPQHuGtCHpgHY3Um2W/vHvcxghI/8s+dKVOob8O8r/ucURxgkT7jqq4+BXo5X
6+SQW9K8h2Ze9+B9wtxGFaBg+tpKdGkAGPRWgswSqvjKvaIl8jXfNn9w0U1q0TS/H8t+/A4CZ64H
phcFViZEu1CRJiQU3mV0XdJwBH3h6NWb6pgfwy6upV/ucmJllS6BzPtJS/pmb2Zkaoz4FK7sVjGn
Puu/mcIDHdceyqdOpIqp2RiqFETDGEEyUkcJSPKbycpfATTpJDA4zMnzQfFLfPMABTnby0ILab/M
NDQORYo21XYa/tCw4zwpbbwTU2pAW2FTJCczAx0GyfZOwLi9FVlKv3UjBpxwu+LTE7rsNNsYUefg
qtiLt/tssZLnJuFxwyuuCmOb4FHjJ5VJUh2kmbn3lQa5QdBABw/KjRm7qsz9gzsC4frtUkw9vwyE
cjpbJNdGtBnJdJ2N40ObCUGdz0K+vIcL9p2VjGaNVD6PrJkFR/pB1IqipDcy0UrBxAphPLMXRtIb
9Z9x5miaToGXVLUzrpK+ek1mSOyDd4plNlrRJxVrI4m8P0vALuh0DXNperLSpoGb0xIVa5aXltzz
5IckeqgJhwy2jD7gf9CMxJQWs9WYVtTl7Wi8sD4Tz4czJR289hHT3Tp40RRi1ozzlGXgFac4miVb
mnflBgYwDcWK4QekHqB5bM48/fkTXtEmSjg4jvBqzAVg64Mdun0Y2FqjPfoJmPLM43ccMjuXZJa6
+tjvnM3R9EmOOTtmBzA1ll0m1NdMU61Kli9xMqdE+/eseC7Z24seU7b9KhH5GbxZbhYx0qoKfJan
k3RJ3hV2KsGq8KKebNPLQJ9pC6zTrgFZkgAC4eThqgnOCJbIklA7/ONqM/QWLdxRXaruB/ZQ+dw+
2VEvwUPzadgKbITqgMllRU6GGisRcR/3EuhsSpKags9JMtMIDoLNHYsWLEqK3zYdkkso2sqpflkF
rOAtoaBrnOKh1tuCUOP1QMJ9Yps7BngCiDA5LOXjPx97XcgtSFcQiNsS7HbWFDf7qwhipU6Tzam7
bJZ3AMJnxHYLglhdKUM91b+Hx2tIGWlfnCSy7QGZEgburJ9+2fOXnTsAUAhRqfDO9XTfcx69d0w2
SGAQdcLwVVdyF8kocJX1ZX5BfriR/4FI1hEav/dtjqx6qKb8YTRmCzVMx3IfhMd/dZup6E4enCIO
vA+3YtlQK5pQe7w6Tgv8o2gumlOxmaodZBf2twc3Ira9XCyuA8msRrSPtkREb0wBBAF79KRJJFnA
uI4v14T57Q1FlFAkVauYQvWHEYDmEfVFVfj5K3UZuTW6Mda3dN4uqY0PRH6ehsJ+WW/7gGGj+YmD
SoYkkUdKMVoX3VVl4nZHz6yRwJZNYNfyh3azb/RHhUq/iL2CMEBoTwY7bLBdfeCQ+RdYlPgDVipj
2AdoFjEfEakwRjmzS3ey31PS5t/2UkwaPi/CuUeUevymCGVAHGHWfParhMc7eDwPO9/JP1Sn2LZH
Pnn3/YE7i15Nx6eca2jm4yvpxCDlMEFXhczAL6fKZe6Dq/XlVU6OK4019vQbcJn5ljIBAWM+KFzy
vQl6hNdEDpxoKRK3xDTSRdQg0VKL8DXOosrcgtLDsoGMdC4n39vnXLKDhVkXl1CmcS5yskx5rRxt
O0qzRx52jC/CJBVh7TIbC6+++Wt16xq3A6ERRqXgrtsMxUqfWKYoRNSFMnAKvzcd+1wEg5Etxhoo
SakQ3FYj6SSCBLM4jXKxqEzIVPZwR4/7LzlaEJob97dzv7YxffpzwqwT+XX3Qti/mWX0U+Oefxvl
YrIQMdkm9K9HcHkOWuyVv8sXUDLBgc340CGWtmj1qIKQoyrEuESjCq7eNFjKYtVSi5vJTfamLBRA
eSjDD1JptZpk3HMSuzXlLuWljP1zGjHYr56BxDPB/2ffievXewm0HFppdWiypWK9vmoSjMMDxVr5
sN+SdRLKYK+FkDPap6gvm7mOxKtbtv7b054g8GdIBO6pMfuTQWXHIIr6KSsoRmRDC82JpxcvghbN
uK5a/EZ5Z81neNu1BTn2CUt12+1AN5OOWlM7utLaf93sf0P+61MmGvVNfxt75NVvyCgxmhmu3Ivg
AZ+f+wShqaJ5WpERddcQMrAH9OHX7KJViz6XkCXLY8gzfsQZgiXuyV2Bvy2v5GL14Ek5bctRCO+i
bsJAhniPPxgtb5FIgER8FxlDYpvgjGhBoF86yBMs8Xch9Jb/oMaazC+UTCQkdmkkFLrWqyx88D0N
TaqwmHVa61AVR/2PV5c0tD5WozaQJkHTasq7JlPbqBsMQ34j2fcyBPiK+b7CxeSkwXvX6mOrn4n/
+w4XojqqmxieAL5oxkwwo6hXJ//v/WVuOxRJEQnU+lJE5iLgEw07uop4Es10s8uMtKf6DQFIQxJV
ZFrylZcIhjZOHH0mPEwl2j9xPoheH8XHr2LfDg8uA168TU/17v+U0AHPU1tamiLCMxOUGXmBhfpg
bzeB+MGlSdwaPnDyuh/OEprTisE4O00/Ym7WIDgEsK8+qvYAIU0C8IpdzaFZRcNkqhC6v/jD2wBk
Y/i98/mZ8LqQSYqqFHpuwFr5r3r62h+YdDWNaT51H2p0GolnddJqWXSV0AlgYdOVmuHu/7sHCPPz
DuaM0hgvoFHG6jY6PW3C1+j8PEeQZjKzwoeZFI1zh3hVI6HgWHBNY8OUSNnbDni8lXywMUUrWHke
oR6tVK2HG7sHH1nrV4hxXvMUZXIFjueOlBcKX4I4l+zkpjr0Pr/CKWNPl8tH1BPln31vfGSqr0GF
EDIWyzUAwVDmB112ZdQugBmAZqHkqXxVPf00kkeeybmDNrce9m8Sor/7mqK0nrHgM5QbC8lKn55H
Woko6kuRwaaeJtv64AM+E5jVW2lXVJiD7J6zYjuD1KvS5prVVOOCfEUmm1QhOQqZcJft9peCS31T
ZNp2avZxIJgMhdQfHD+qm224Dmip1x+WNA1FLlhe2/7BXfgLgx8rrUBsqzGRqh95tCkJ+faVpS/o
b1VbWd2qjeGqE9Mc0V3Z+5pjSIdYSBWNeRW6CJFmGeMDHDTgp/G1Q68/8r82X74JvND/HsGUNel1
y5CKNpJlgwK5r51a+3u59U30RPX9Sanlq9CEPhgIqfXzuha5zkQR7gB79hOzKXNpS5eWtJe+8T5z
8jZTWpnkvojLDtgrfNyn890GpFzxO69MO9xjthSifFn3d6+Wcjg6am663KJbsTqbm2hoAadyafVn
3EJk9MFkB9B4fjdLDjHPqEPEKfobQ75RVXdxLqgtGuZkjFzLFtC7ee5lMc6N4i+gvbsFmKPbXWHr
0IMWLuEVkDr46KSqHaNrXAy7VwBWe3aqojQzB8NrsnSibUvw2fSpVc5lxSxHI8Js+/Tw2gSgmB31
kCHRwIzi2XF3zIwsc4S57jz2i7yVKJOixleyPk6nYiL6A0uqSLgIKErm5h4gwnBIrbDwfo7/HMSC
nGtezyT4EAJH4i6IFE6UIzetBaWIP2GdfVIs6PJehHR0InHbgx2aRj12ZtZZ+FuoFqNa2624U+x+
y9ZmsLELat9fPTcDaBQ3dD4w+w0CAsIhr1UG3Q4h4912nARY7UZiFsJCVaPJzi7KWUltC3ZJL3Fi
YvfxN2Z2W4ZS7Syl1S6eSEiBqM2AkZ8cdXLeOvCH//r4xBqKOLU3R36XHwHTiI9VpAW9NQ6MiyAx
j36X0XyZ2KRnWCTBBWP0zGZhn0asDYwZrouVd7+ydGGKyfYF/03YVluet7HQvj3LeWox2Aq45OGQ
OJJttwe2AR0+tV4FhxbLT2VvEMfV+Q/wOqsOx3YViG7fKfvoHvB1aT3miihVYZxy5dlI4aDcINqK
YbWDROjB4PqsLCvn0BzawswvpEoASwKPaYkldZDi2E7/4YOKMuB6drKJKTEGDIXyabo6drXPxd/w
NkoPh0zNMIuFYuxxR0QtYXFpxqkAHPG7u2iVOsQnKGNhNs2XEaFIpD9M5pcp1S9xQ8UocNI61fZ+
Iw8P4dWFNCAVHW2IFTadBctPh11COBLnP2ERr9eQ4bAEOh79kBgLCTbR+LJKrACpo3X2aDbx5ZN+
RT/gQbG19/EDM0Gdej+m/Y9G5++p81297Rc10Y+bvhjVosAnjo5mu6FAGCzw4VYfJRslzo64JSAX
Jj1HJZAEbEo2ASpwvB4xC3YR0yvXTbxlwtDTy8hPbLN4lIJYM9HgomHYfwyzPh+bvQ/FnUOk67Mg
MWaCjqAhiAKL5xg4i1Opn9dsEJI0nKioThMzlIAVtdAnqd0IgvCeudO8KmGlX4nmZ5p7zm+29eS6
rD/rSrsw8hdEUqXHwz1Gqi1DpVX4udQndrgey564WiApIuopPHEzMSbzwbW/6VbVn4kxzN4sx/Gj
NkO4aMutXVgUE29pz78nwOqagKbKSP3VG0FumT67DChTqC0X6ejNgisBqQ1JyDoRe/s9/E3dAa7j
BB8P6ycL+V/l/BOxejQxlt/jzwSlhYwA6bhABaCn4k7XK6D8ZXBHTmGIiJ1lVHbpXbG1T6OZvSEL
jp+/zVwo5JiWFcpmi/ZI+YOBYw4xUWdQSsbJF+uMSQSIJJpOWbpuUI3NipVx38Zng16I+QZeSChe
+Knd41QlL0JOIWRhUC2cLhzXdc+HTzg1w9YyMohme23SiJEQVBAqGTz8bAhj7v/IE8IhEjrnjWm2
hNeZsvRWzlYPDruw/4gkKWv7mOu1smauBNRYpm1IY9xmOZrE847NOMEgivQsQhElqfeTWaDsHvli
B0Odg3LuNSUvyz7WGkrAipBdb8cYgRADL5xrZhpgzsoX1mnmB2XJGo6h3u0VVfBoSN7UvZSU3b1S
37w5xmZlIViMlfrebCyydYWInMK4D0B9SAzFYLQbmSywFqVZQ14kSj7ADKEapVwDVg3NAlwFDOlE
3fW+2Vm1uHQKQSUR4CgOh3Qlf+JFLwJlFdmbffnG9fwcCynTiDIcESK3in6uN4fuvQwsD3M43nGD
UljeiJ3I+gBtFFQyMYdVUaQZMFBb6bfW9enHtP+RuT5b7yu/wyfPWRJ4G8ulwcMl7E1mui78kCaF
5FeOvJBK60UCKhG22CdRndpbrZunTqoxxiB/qU+E31icAqwB1gGOTWlJjTAWJ9lgTlGl4f+EEQ1n
oScRZL3giJI1LQJHEKGufPUGcpfsyvbmMQAdUvxykDLTdwNEs4KIdSAvGBK3Ve+D3HiYQ06BgMUK
1o6NMg90XVbVHKVOIi3lUqWuK8oQinUOnjgdhGS/o0As1g247jhnaek365GNjxku7yMwgzlDVLjU
grAJswVZiW2t1/T1RyFtMF8yGM1yLqn88e5UfBNh7/vf8XMmT2qMp2Z6wWJa2ZelMKmDN9qdRNdg
nrw7OmQofvxYNM7o25oRhtVIs/5v38/vYN3j9/kYxEOXg25rL3Qt9weDWsfPmHrImQdCaPgTvI9x
WbX5Jqb52Z5DdsEThl7t/X+4gakC/jjL27rFnO39KPoKdqKlJR/tXAGbkagXwPNBZPnaeiWYwvxX
FFoEkzPQU+Au5T/3J+P7KDAXztvfKdRSI8q6WXZ/Dz66UVQo/B2v+kuVkT56nnfESsjdmJIubYYu
6+ENBQHl8/6AMBZ4P+ohvLqVus9QWH+mX3jqTmbe/zgLscRlFNpgFrr9rp61srzg1M7fity0xn+A
A6vYW3m9mo0kk6NsJTcgg5Ymn9iUzVA+tbdwEaztXZkPwxx84j+8oMf/Hdt+wRsdbzmm3i30o2N6
P6RG7Zs3OZUXEovF0C8qss83QVe0bRvn+K4ttpKCmS0aiOkpfMBAI+KQXDsOGwENiT5ZUPxexDml
FW1SYKQqP6gjUQi9x/m/K9tzD3OkPkc/t8AiLGRItZ0kJ8jdnH42JmuN0Q7WAMaUr53q1Eh0hld+
wkhZBiUi2tTyp/w0yFLMwzgFhFvRUwhLtSVB8gLZfMp81nUMEKTdc8tOyZ55ooYjNFVxgRoHyK0L
IMT1FnNnWc2aO7eI6qyM0haEeWYmC0QAy2CjOBhGpHB3aqaYKqHYoxHZcnm7t/VVdgJiicVIccSu
I8ZoAqiIjSK59apRo8eGC7PH/2AkVapPLsDFRNwJVKJzJ4fwM18QVcqWoJXBB4HQjrmpzJo/4nKb
F7Q52Sy1sGw2Z6oRkrY63s949HDauj2N6iPSNdNkQUfOMC6MmNRqUZhUrzTwOj40GCNoKEhmGM6m
3FOBl6cRfzDFIkrleHMeTT02hLn2YMInR2NhwwAf2FzPjn7tgNzhF+mrRvQxKIw0bY0fBFxiddxV
J8smFodRC6ZFTdrVgH9ykznIITfyNaMo1RUPbgvRsZlyAG8UEMDvwD9f4/X6mBcZHUVJGwMt2CvE
0UU6O5kXw33PUUKV5RwLT3aZxIOwlxvhEY20CUpltiVwBoLve+GiLTbU46RyUqfxgMWO63Oy5TsJ
pWrm3A9qe5vBZOKHPdCjd/vD9EtaRZEDuW2UPFJdnZsmZg3pnnPscO6Zrvq8Y3nAnZdQWkVWP4Iy
UWleCqsN3oqii1mx7LARqlH0Eg2UycxYX8p+Gi1d6lYQ6kZ1laTFaT5VzOdw1E0luNCOJo7RB/6/
8Ox357VjsVWS8TPDjFx2Hf9KiXfOd1bj2eTk4SsMwzrSM9PyK9doXaQAh4Im6+nPpUsGQ7i84xFI
mDzK6dRUopKpLuURWU/9uR0wVUsq+pWRzTPgALl13BHNqygZb1LfxYTE27YOlPP9mkQVpQCsRgKQ
fza+ujXs4R1TTLD4vcYCgMd3M/zdYCBZAAJ6civjRiqmNjmlKkYzPACk/1VJUnCHoxbqHMEzycAY
lIRHKRzzuZxx+scL7wVEu4o2pb4aW/6akaNfUahMQhq5iAwnZnj+8sc4Iy4za81IlsFzCAf4923N
CaXvugkbFim1dIc7OAGRInLuaxS/uCPKrvBr/3YG4pSay2sl2J8izeJf3H8t9xljcfkoNMCbECLm
28Xt1rVNsbyd8b7EFvRdYJxXPwXsuar+L7vh7JM6ratx9VfWVN+JP2C58Wzp4ZESBbA3Hs89fefS
eWY/XDcxe7NO2f8ZH4g6Yf3Aozb2MGbrO0Q6xU/ObADDCsLK+mt/sHNH3CwbbILWAuLrvFIGVzN5
0hQseYoDVGBRLwdtfKgeDffK2c2GJK6LqkyGb4U0wuoDEjePUBD2OgZNOQxWQZ5VlvhjabKXl5Uw
b1Pda2D6XqnDd55EYu7x1GpMFHeAViyA3CbhQDsQs+vclXdoOcTceIM/xktMXTgiv3u7352dFhQt
fIh6MjMxlxzJJh6JX9paIJ2zZ+wAnhpWfIJqWlfCCvF5cBIsk+9avaxwiuCr1fAcdFY2o3L0+YcB
ePLpZsahHjdjpbd2f6e4uLVADhE3uo0wKtkX3QsUf6lxOj9Fq7mGbaQ6K4QLXkyOyP2SO6c4fqsS
7xaiNUoENCWS10m9RHygTGBn33rngKHGzyTJGtC+7143peHPN0qz+0s9XQ8hOwwg3nFyIs5RiF3w
wIKGypoLQR7XmUyo727qgoZRK6yG9+KT/CDw23zKZ5xXcaau+WlcSJNwKgqC0r8L9Qj5SSB0UpfZ
pSAdqupZbs8anfnHbmWnpwszsqMLOm6tpef8ComLurB3KTT7e4XKYCGBInmLjOX2y9oZVn9KOnah
T9wHeo560NmRx+NJdDtz/MC9xIfp8H36m9NcCBsNToBxWIhgXu6xGwT7EiBIOJDRL4BtsYiSQE/m
RtvVjtHjnA4Q8Kpbvo6aXCReA3ZqNZQdAaAj5WrHEB5UETQvVhoHLdxtlVXAt1ULvLQ6Ta4T+T6p
gaogrmLo38lF5hVMnlhFcPEOXPT5/r1K3d/+2hLvQr4AlV6prtmOAFTzNUSNzCu+WMdaV+QQX7ay
BcZDwOc9JM2LgNUcYoU8XDPz3/AuDVM3OAFXVRuCUji7lOluLyCif7jRjlUpYDFje8yiF50zB5O9
HQoaIIdQkUxqmy0K8Wx+dWmrAwVF3WxTIiz/B/BC+nU8cGEbvHoWtQiBlaIGyioVvPac6fpKEzcc
L/RTvsQgJy9w25WE+xK/6F2+swW6K2RQqPn1hSiKNPtZQQqVKy4fPpPY6FGRj2UpkZ2nCmwm4VPX
lQnBNoGlQziF7OF8x4jYbAuZY0i0AxX7EtfO9YiR8GyPMKDcXWXWpF6ga6GWY7x01JL8du2UEJww
8FfmErNkOrF0YBg0tt4eK6xFyb2DpTazHLW+wf9iiXJEjFcFAOiDhqoNGfmUdYlXtC9MccUcZRpD
dma9bhlZUqTbwqSLllxfDpVQQtVGFTmsIjg7D17p2T+kegxgicqhgOdsVKK6t7dJhGn5wmzOecXz
6WGIWD//32Y0L6NBTWh9czkxHdRxhtNrB7nQ5xVw0keyhhi9tJ7RvkntlqeO6jKoQI+T6qaxwvH6
5+STVdcQqVU3FImmWUxlbYIvaXhhasyMb60oab+9X/pgAML9zxYqKl7ZrwNeVORVf1HNjr5uyvTS
JuSyQhDkeaO9iQsmTdjrnXO05s7gkVM7EP1dhRZUFrazmcgB2AA7g3+FZppIDBQadci4QWwmZCHs
/v0+KUTCAY3+ZjRkUlViFWYXbKdmHQ90jh1M7PfItv2kmbwRPJ3PiOP6O2vS2uYWkKh3pjrwVw9i
szVQENOcpcDPinAQB7oah8RucIsfCLjJ6qtfxiwrXdTb9YPo1zGL2b3WO5argFv8i0NaGfxmJI1u
GDE+MQAKSftBfUHUi0w9d6RAUYbWAAqfQ/Zmwp1p0wsxmoaunVHPF4J+wqFcebq9goA5XH9cAXjD
QL5n0uVJbl9GlFQsWgyMsjeJDD3DB+bmuyQU+Hrs+ENlT9/+bKiU6/UkZPNKyI832+gkqgEO+rQa
Obm+WMHRGaWM+pJ8zM4SWUpAJQor8he71dxh9sF6lKhxSM1t1VP20wg+UhSBGbUP5J+sVBiFmKlx
sFJeLywv6HfYMpwGgRQ+5Ia+qMV5vI1WBL80GKmspO3HnBdAJOo58Vn1FjDNp8qemkN+HMFIgbLQ
C+tRK6odNfrSyOaT4GF3izzkd+hlbs0uhQPgCYaJm2dVpTuwv5D8xOFJil7KUoSk4/iKjbeL+qn/
ix6Mhr6PXTXY8+yQMAyXWcEgI/BdFLFcSTc4etN8/dyPS5aHZgWBfExlgAZ5AFMyVjjZcPm7bUXd
szO07OyNw5+NkyrnDW06hpe8AwppYSlZlqznZMQECIXFnS9sTnKGUD9W3iGw35KCYbUMbS2W9T0Q
+vYRZb+ApxLhrt2UM2sO5gsZ8VHgM34caFZpt5sfk68fsy+XofoNDQayHQLqqKl0qqDp+/G6JWXt
SmrSQS+tK3RRf6hU9U/dkVolcBriCqL46TKVrn0btkUTva4m6CuKSkDEIGQuEffBlHZducPIY1Qk
XqquCdlJVLA3GQnHUJWki14E8MeQKQBkusdJmAtNCJo79VWjwDzOQQWb8umEKo5oc/uoQRNO3aTt
8Wq5lp84hPjD2m1aDHuNCwo009b33tRDVg/FMad+Cm81CAlhXVGv+wJBAo76epLPVH7AwyfON6nL
EtfbdUBpibnIONmkfRgYD0FKNMN2S5IUS/mmVSlq8xAOiiFVzWWUvgyxvOdSQ8cAJuu/jPEF8kVS
Uv8mrx31onTwDDY5uc2ggP+O/Tj8TtDmaYFxLDJtSaZrDlbtFZAHKBjnia6L/Rpd6d4UkcMJ/Zlo
txnUgxyXA5SdUlsFshCG8ukDb8I9W83RHjlnTY1vwC2bx3vO5hSwlkH+L5wxn7+S1Q9bTQVLRGTI
2608JpfNZS+MZQcWjogQCoSAt9pOrLj0yF/HkymT7Ks7GVg0azyVVY9IjiDH0MzX04Cz7y9o65+9
1P65WPlx5WLHW6omYEpwOQcY4ZovrMiICWfcZrUnyH6+kpzSvdPEwPnwMcdp3ZSJ+4V8ue4pR3tz
r0ne4bTLJaXWbzTCLsSZApjMtDkDgmirHWRCn6PCBbSgPl5B1rHYasZjJ37hAChiGgpMuC/k6dgF
vsrExI/Q9sm6ZZErgu+OdGITly1SA10DUvIiFJao9bK2PoPyxtvMqbjAitXXM2K1ZoWjNWBgTtWG
iNqujd55Y/iTp+BAY+X+LtzFg3X/9A800RJSlN4pgoa2xP9s49V3mdzVLaWgsr43V8O/Uupf91Fk
oSJ4MiEchy1J7YQW1GZdDnro+wAPzAWvCnUj7w34OqdeTEAbmo0GOjZ2KDV2VDIXj3eXPXj0lT37
JB7EvjxIwiTaA0r8l8Abdd4ef675UQkkdKBcGpHfnhdwmqRkL0R0uUzoCULaOOSBzX+VnWZLGkQY
f0oAv80SLAGuWt5QgHIJb+8DgFTZR06x0F2tA3GiU9o4yrlQTrxtMwaUQ0/wNxO+KWbARBea9bby
/ePLInmqGuOxgYLVfNLAlmN91SwI9vGjFdmc3O98+WNMV5dphEq1UqqZ0pFLJAhe6/d/kEb8hCBR
HlwdbsHNcFqjljf5psUYwOU4t6nPGJYHHVE0+USbkv1/q54CzM0yLdAqXFTlhvbskIkhm0ggkQWS
H59CULNdqN4cyInUmQmmRCsXOeffQqpXa3A9ekuX7QdPpFkaNSkPyHn7QNsaT2r1HpNFE1jI5G95
M6TDCDVg8wWdbvSBsDIED+/GRTrlmoUih+6KDiZQCEUY01VA7eiZRd/jrjamsE55SVfuS1x9XqHt
eBS1+cnL9F+DI4oOEux+htJAaYgUkMq0BASuiQkS30WW41KJDoGLscA1zDe7Mm02OsSjl/acXNd5
n/ragLgKF9C5VEHRDGKOl+h2F35NGFVCPvhdF2t/acT+hdnYVEB35jHAGymjJoIuWNXpahTwjK+H
RZQN2X9vJ6o1OK4nHNqAkV/NugkIqtYpOrE0m+A4sV9xYCm53IJhtH0yea9/278ApVjjOsAT8FX1
QNPAt2YDxldrcI5eHyVxaGyulehF2QYjm611EOmDFXV7zLfHJU4Jlka7cQmijtzqMx+J2aF13feI
DZfex82YO3YYzJAppqzRPgzFOKQd/t5Q3PoQhoH8VZQ5Kqr7roKaq5yQtO5yS6ROWSRT7lkxzWtn
m0A5R051w9/epw+QkhDZkVCxVyxzJ8oP9tMuJn/qZLvSszAMOmwk9obS7cHvqAAqmNhhV/OuT05f
amy/whVbBvwNegGP3IIIBmOgdyqXeCLkXhwmyLPsy65CRVMMp76ix/s0++IKu2MpQf2IxhZI7QE4
zMcoMyLWHAmUBaErn83+qo1cN0l5ikwmwln3dE+y0QmAdb+U3xDFQ1taaJizz758tcphc54/0x8H
OdBbDQ5ZizC0c7URHJM6FRS+gqxK906yDkqW0D7EhivoRdtl8L/DdWNYxveS9qsWYajQHCyzafNG
Jon7DPO5Flw+owMi0m0pH9jugXelDa2IqUVNbqF+Wo12vn80Ylgk29Gk8M8lRRck7GfSoqrf8CpL
2sNMS96DfY86u8Dm2d6OvXBj+Hod9QltLdlPvQ088omYymnP2GnW55mmGMu4zTuqtXfG3Ej4PQij
4/M4H/JSYTS5HPtCrkBNOrJd/7r8QRKW/Sn/sykoIBIioM7Hyx1vhnkfgcubF2N8mPUa348KWvFy
GZKEf8luPcM42s5rugZP2t4KVJkW6MlOHq91qZEz/DUjdArURb46LhGzmc201a0b5OQkp3+pkYjW
nrGpoUcepbX4KxpLVHCWVXoIWHztmgv8s7M1ZxymcLkNCjtdzDUFHv9KJapbgP0dj/WSIGIw7Gol
XgQBL5OZoDx1jrP77ineL/PvxwlgcrzSG8xdmbe7wutAbGYQ1UYyy6rmYal+U9g3QASji4WgPwvR
sngnYT8EXsfuewHanjUluFX3t5d19NG3s+3z96oMs0d3XVySoqxFDJjyjIA/wceMvZzkRBmH7BLn
GmjsfqOdVcGK1dIEg7XxzSWLuFd3/i/9dwJL/wux/rQHuP8BskeI00domotPSr3Q0OmlcEtPNuvq
vnijQiRRS+j2fghjNnTmA6K6IguTyRWxHoFYlH29zoN/4KGfNSz5+QlCrTvZKPhxZXyGjtFJxcwN
IoTPjf066dmCvkkSbfLwVXmSBEvfH65dbr1BYwr3XgZ/5WtR+LZuqldbPIGbfyYBtq3RMtz3gby7
2JbnYrKzXnAKN4zY738jLdO8uMzMg6uZvIpKEw5USGMGkBpSIkrTLvwNJIFcKhxdnFKXR9ZEmeYY
5O5n657tadKwgy9RjriyUuJ27C+YFY2FAY4akRtz1vxHDwjoZ+kik69weeSwZ4ZDA7hEBjEeNeLz
sm82WKzFtB3kNrJHw8KrkX4Z5PDhJl7Pif2ACklicarFZwc0bstuKJM6ZsxhaxOw9y+UeBWWV35P
OkOtxTCN4yU42Et1h2elFfHtT7nfHKwa+c2+dQk2m7ZIMHKy64FjmmErZOOi+Vg2GKEs7yK4YQTM
sqLsVy3/XGSCrwOscINJAoDw60F5q1xG/qaGadgK1+tapZyMAR8Xic7S5+zBcQLIf4v3QwKAiyBz
QE1VeEPJkF1BJNuukbA/wGL4LxZy0LY0JrGtvS9o6+yQu1r72lzEt/FZB+GlcIhucQwXkoZwPO3v
tVwS3v+MCRAI1MKkvfvzlvO4P4yc/saqSnCHqEWnqATFZ2c2YIMmEm0OU490Mbc3F2NEtgeYkI1c
HxkqS7gSkST62K02/Vtp+sZGBShcPE0besRXKTzrU2blFlD74t5PVZZADVs3oVOUQT2iZMk5gIJG
rdg0Rtx1wBlTx+qQJpX3B/cNEp8odcC4ZihqFRqcOco/t9oHSIJw0AOFYt8cVWSdNZMgketVLNOr
PjfHlAxGCXVD7VG7pSd0lLEY6jUsKa9YT1lmecQ0VojxQBurUwxaptcRNh6G+SNY3Y2U1xXpVcvZ
11zJhDyzVq9a7y+KSi7022xmHDzCBAZjx6qVA4MDy4UeFlwg9qQj6gXR70Wr1Ftnnp96UmyP+qiY
KhHlHG8GVzoOvelyPYuS2M27g3bk9GMKo+mGWTd0INDuIhMDK/xX04hfOeZ/R5QyXFtLxGNywVxK
3nwlstVlnZSRwLAi606VU+jzSGi/UPRcmh12iivy+B3Dp2pAUSqpgLSD/pg7QNVfSdu5LKaqhyeF
nWl8e0RTXmKPZmYZL3HXY3CRixuHOQgGALTUkekScNIbjJHOPyMJYWtIwzsw6AW8SZUqJSsn/XFd
EGGrYR2tRVN4pd3Enw4ubbYvJMK9fGTw5zkRxVjkBZATkNYYqGLCtxjvaqlgqY4r9fCFeCwpU8nm
Z5aTPRX6+5ngZ5H36oFNontwzMFR+F7N/zppa3dXer9813Q9l/GAF76meyajDKKtCW3E8ciJAW5b
sxzIeYIDVXHlsfrzOHOWBCAy13aG/h+Lu2ExoPiZuf7Az1C/gjf6XsevgznRsWeNbd8BBM8aL+GX
PoIObZL0epf3qHdVCI1UD3z73xzmzWEF2z+egtIepQbN/vfq+tLoptnQbuiXg2RbNKwCtPH6paBB
8knUpALJ4QMgtdJELLtQCDIn11xiEkyApmyOeSjyD4lduqzkaDLEpZdlav8CGUqEVSMUr8+7qCJC
RESivIte6b4Sn7gr9hfg9CBDTWjbunV0BgcdvdttwGJlmrUkn+2Cz6Uq261O9ilW9qtB4bqJ5mW4
rJ7YPFwzdSaCZ9blWU+GemH7Q+XgjuhqqIHuUbYqq0hIzsg/C0JC7BOFV9d2eWWgU7iToexpB5Lu
kj9SMUtNS3CCVP6687aLAWCbwDX2eUNT9FM3wWxCKUyAjhwtccnw/jo2JzneZIxPhATA6ILVpStd
8wqr+dT4DLHwZlnaYuQ+SgY8OnWxHNz7IMe9LLNdkCrxxX3dDDm8eZpceInKLCytzW5S7+fzPL6P
rPD7pc8h9X18u9Anhc7DJwjBXBtzFunLFzieebjiajiSItS5C5gLtsBtSHgIDq0CyO64jKJTcEY4
oHz5C7JBWSgEaNLem/8o90Hzlp9/F7WTYG/KyZxVaEZ/HaYRnOJGZSM+++EJhKeq8YyD9EM+sqPa
l6GzFC6VhEFGqBO+pNYoduiLJG/G3YlFeHhcAOr2hfD8jqQQ/747Hn1hy1OnaQzY/MRumFDiE26G
z2ZtTi1ITY/qdWVX/VvY06zdbgBv3UGy0wiKtYNYTPKeelw17xOa7F9VQ+UG6UtPwtfCk/elO1mg
knl4vFfqGu+2pv6ZfH4Ccy6bBmHsX9TauZLodyPlRtVkt46sjYOdQxURCZE8Ii50XCIjePeu1+zk
vQY1zujehh9LOERfpvAaA4FNR5GnuK4CVLB7hCRqPEEbebSsqpP/5pjm6cZlu9Q0InEgYeGs5ico
7IvNhqQE0qMYbH4eZ0np75omhgQk6WXJzY+idWLWgf9actOMaoB4v9J901tccsrzzDUI4BPL3LOy
3UWXlXiB/2pN5MLO9ok9xYILMbgdOqYo6NH1tEnVvG5XjSjb4gaL46ot2q22/akmrxxDb/qZlVy3
cqd/9d+1qfHoVMaQgREauJ4de+iJtat+YgGswYKkSPs5VOGtLHurRMxClya+vBbVp537KGCmgQBt
vxwgZjpYANotGIk9XB2nYjFkW18ZfYwWrKoWSVJlnWez0H6CfjwH7Ru7hb+mtCrtD6LR1XZfhkRH
210ZehZSKLIYkMbAOP8wRiFI3tOPgpeSefKNdM080R1+ObxKCdpE7ih73Gmlod7tVftAu4jutRPj
0w7ys3qYemO0U5dA1r4EQm7xOZQIKy9RZjmobYoV8B+2Ued2VQaEVLKyhChKlfG+2Fr0awpdqFSW
6CgGFpC/3qkKiLA4/7Q9itkEOkUXjc8+f2KPRld+ElyX0hWD/Rbbph4/Wn+rj/Fk+H1JJH2fSwXP
PdyUgGndqwq1AAsebrNpAOno8z7f8aGD8jN0ZW5qnltxr3KYl6CB/3DD1yE1c3Sq9WpJ4UtiMvnZ
3FXXsJEOAcHH45cGs2nb9lHftu9SlZy2jFFyPg5pkwuez49ESnB1DeG7DC8Xnrv3Mukmm+0fCxMZ
eFS0PMGVSAZZSL8M22roYE101ssD5nt6GzAcakOPzVbS1KjgqmkqAZ8qTeG5algiwUuL+HOgW/pj
34HnGwxyYHTmihPle9K3d2xCYO0i6l/n0EizRATaXUO6TfsGDKh/7d4SpM9jVr3WklfgUqKfKCGe
KESGiaIUhvUv7YpiscAEccH/7uQT5qQTbHldtGeFYsyjnn66Cjsrx4k+CnH0O1l1MsSTo1VklKTG
/bAo+Zr6rWZCTgA55is/7kFy8GOYnvT3cOPWVnbfM9rL57CuRilPZR5MaF5gOreQo/v6dpgEOxXa
kHKIB+jQcoP5YqXgiW22A+Cbog/dsVuijMiKqhBj9wflVaOA/hw/ovlp3GXtGBehO36JWph82IRb
yHg2gGkIVn4XLxXKVbiH/6mkscVFWkSk990IoSCMNxkeFV5K/9Ovj7VztFDc3f/GiOwmIQx17Jzv
vdMpKsSRl0I7jTLoYew8NcMi4Yo8eWcx/hp8WViIRLXwftIkvG9unJKuB3BpGa03EQrCuiN6ITEc
rt3QvxB+3UAMWzOPZa2S9i+MG7EFccabIv3YRWIcq4CKrJnPa2mLJPypD21XRG35A9US7UX/nRZk
hE0dryUrnIFyrqt8zn7sNeKoTHa0ERAvKmSAWjfTxjIYDw30m1KeSo1Gd1x/KmXvOSXTKBW6Y/k1
xDq0LiSk77svVn5COtC67g2bCywbzIsypuZyP2fxhJNXmeGDMbGkoxK3YSqAD8kPBms2AVOHQjOE
PTuBrETlym9EVZ+RHF+mLz/8INx444x6MIkW8Ddokinw+sY6e0hCRDbyffjh5yOISq4anteSCDly
yDO+puEHOVijwhJ8pP0yb5VV4dhGFIAbNiyugFjMJa/tlqbolj+GZghrPrI28f/akR7euEYSoMDe
wkhNVDwjHfljhg+TfvvDe6sZL/bucyhoD/MGskIoINcpgVc6nsWGjnmV+8BwUbMKjiJ1rU6Bd5DZ
lT5OQNxZyhGIZemiwvwRtIi3bkLUKM7wF2eiJ0t2idCw5QQ1E3kZT3ii7HqRtm83mhHohVAHcDHq
sB8/UHVIDY3/16VIbtappLIRgaRr1fOBOIJipiG92c8+5nthR5QJWEtXpgiGuPTuh2p+dT22lyLp
FoMuy5ZZ7aW4uWfYkU7EKVuvVqKo770Y+mRxDPXrcZNO1T8zBnvNV7taGZPQ/QRoHQYkb93yGy9e
9oX0CmGRncbt50Plg2LdIuJMZb1rh0bV4HvCIbsxEwSadUSlqcpwc2/9XFhFbBlKODcbaQSw6/u+
5Q+FvvWUPU1n6pTWZTxBBXxUOaNsH90/svK7MKgrj8UAScskBHBR2Nd/FWlNfzJBNCCGOgHaF350
VT64RiBzFRkAveoEBDgiKNxsPoGmBY8jUbM3moreLf0CzFQA9jZzl2lsbeTTmAOqWqLPOUybHA13
PdX18Lw4wHeeHuK8ihHkxHAPN1EkWjz00zVfQc3e1iOJC7FMWqnwZJMCFqoAe+TBLEZuDM4F7eDc
rxShNJGffP1t8jpnb604kivnlFlaxgP5sDrtSvzmxQYklXcwUIG7u8Q3uoWAburnaskDYOMOXh/Q
Wlaj7oN3NEp4BCeb4gGyqNcjfgZDrYvKRcZbk93/qlqLRxuN+wsHQF6MLlfKL9pouJBheoDwJOnr
uRo4sQTDJ4BwFM04ebeI4HIh99XuJwIG+9jWsWyd9J8BVM76u48kkt/SOb+9ONy8KXC5h0bZXXhq
xATpQpfki3nVR0o06W1lP9yRsgMpWKtU4zcUmvu73Hq26WeLLStFP8BZKkpLYh6xgxm2cKUTquQu
E7zLLidIdUV0pWY11Tc9AntQ+UOdx6U+YCLNq03pr4lw7NKIL+aOymKSfXpXHZpInuCR8MhtJbjV
P0Y4EJfbjsa0pYQ/xwWoiJjISQHTj/vfvuia4aqCEcHpXDZtEjW+fjUrcRyeV41GtmR7WwcYppVm
IvJRaiSVn15f465JS4Q6pTGa0PtBfN16nAgIACGRXASQieyTdwwY43o5ofes45Qi6cZpXeuJf8Rp
ThCBI2r7u3odZbbi275bmyLYFgN/fYo/pLJ716PfrgxR9nVuz4nRsb4aR+bNorqVG2iz6HpyFjgP
j36+v5BOMXKFudAvovi7zkaNne7+qZzw5/crC3tRu88r/m+KvyOFHmNd3arvddJgpMx8A3+uIOPZ
cNn3ulImvM9vNkHmRSPF1nugZ3/xXLXTvspdsISorFxwZQTXFKXibvO/IgzhOB+jJAyyfPpMo4+9
3/Z/zZ/dQJepXJ92cgkWoK9Vj1I10wXRHGFDtr7nGY/t6yyMhG2zqBNY3UArIGkb8pDutkbc28hg
Xj1o0S9HO/Q0LtB/OqHwQogD11JTYKBUI1JCXNn/7c/BKSTmhyICG+ukRytaA1sNdi3QANEYau13
x/R6BmE2DFtX+yiPrOodHL50RBjRg3gsKCzxh7y0Okayvy/TFyRC9tgBgZeZb2eUjiPywTdghEsd
/L3/Bz0089gKJgSOVlEYSvFa0d62B7W+HF/LfDIUxd+KEcbMF7hZD8/Dd+GYWDSp2BP99ljROS36
AvVPn8/2cXl+5nSE7VhSTlH2JSnoIkqfXdmaMipvsN8jKMYFuxIfs83ybJ8o1AFML9Z9fd1Utt1n
2EO76loAbg3kEYqqePMsO7kF9kJ4DrlTvToDxuxY6voWGjFHRaq62hCyr1TnV93HjTWr1WcNAL2j
CkJUrOTTh5qNlYWSwdQHqHIsUcg8ldliWSDSvqk2i8atyubJe9fx/fipKZxOvvRWYcLgUmgheLkR
zn4Y9zSXHHRrdhCZpN5cOzgqJBM7fPLdkid4idy93OAuNHtkYyNljWFbAo/eAvBnUpzYgxr0pMvI
FCHXZumwmQ4wTda0dNsQZBJXfooCVbUCyqTGnetNB31NrRDYls0XuhetelMnRVaV+gwhs2Xz5ESS
7RgUMbXagfa/tFtwo4bnGblIR+IvybrQZMyaFYvfiPlo2aZDB2ZWsafFsrS3N7UuzrtjZv9ulbFd
ZvA2V7rJP3AYkGrJsJTTGroHhNETtA7f7HYHwXztFP3E+0HfWEnkMoYZEL/47c2ttMO2ztGtJ4jT
ylZb4ldbsMp7AzsbIdanJIsTmtdyYATEJHVZDWa2Lr+72+hoFAJH89woobCFL/s71DJ/W2gKz52O
LRH6MfT7bHWWZeyzwUu5Xb3nLifTOhcn3GbPOXIrT1WWJmF9WPCHNAaQQJ76lNKojz9MwdueUKeg
J21eZ/5Ndn96N8jcKhZvd08hPna5CjFjUNdJBoLSNxoT1O9LXEDyuQYHmz0rRMCOfu2bSyzyPcYK
/eYJPRQv32n6w5iBQdYklyxhAU4ztWTBJ8fTJgQYP7rcspHciRYlDqX4Y3hhBgtU9NChrqSQnWGx
i00FUcRWeInP/FM6VmZVg8bnLUqzu6SqZa6z9+JI363AHd8+r2Cmy/Kjc2+cDRykjkpwYnDjcsRo
Gp/wO3aTZFw6dkHy8wjpIBoO42Vvc2uMRhxMThnMWddMO5UzqwgngyXidaUAUzX8d39xN7xWKZnG
/73Q+Ud4Orbzx2P4YA0q9WBS9XPspOuZAINKP/K9mAm/NUoNOeKpQIwH7TZsop4UDbmFdlECDhqb
W740VW7UOWV2MSdO9wr1vTAdMHL63IdldYWaYt23D4qg5D7LlIfkbA2mspiz3F3zeAbH5BhKVwLi
2+sfoqmvAVNx/4qSUa8TpA+/pKKIclKBzAavwluljz+A8PNrR/QXVnZhfoCLCc3lNBwj+Ed57M1w
v/MnQYGM1l6JiiFULLOWNqklX1WTr1id4Gk5aNmAAGFRNLk6Txz9wRkp2VVZGIepfQmS4ScZ+EvC
9pTu17eWWJ6F9pwD4KuCVbRqlGVF8oIpztLgQuswHtDeYc14WG/sEbQ/uDi904DPkI03AkN+Ddud
ZVlE0i0XnFF2GbEoOpokpuUwRjl7umX9HGLRbxFktLFkIUHLp6jB6n6ElSouE7acO4/bpwz0bLIl
rLYf0Ev9ohL/Fb+OswCccKmLu2oi3+W//ct30oKzaeuIDPb570m9cFtJ35UFPma8PBdM83NqHIR9
KqKx3S8HsoP8eTyh13y79DeWLV/etG9X4GPTVxR0ZdAQAe41Kx7dnhy61I896rjaINxVqrC3AxjU
UBmAHMb4rGU92LHp43bezMfKWJKi6BcruORkyY4zgZYqVvOkRZ0WugubyKY0EXuTCI2HT3u8pEU/
u2WvOmF/CNKuCdYNLqeuvNWWqJoHHprxEAAYSxI1xm8X8IxPIbgOxroAkGj/hOjTB4SGwcm/20Po
85xvzCG94iFvPeP/XioU7zPAxEMQwak44bJP8mqXmuQ3IwY9ohA2mgLVJnv5PlnmxAsTEUBBEEXV
91L401C85tkUoKO487SQUD7KYOLKV2MjIN7kT4i6lIL9P2STHGoKhp5lonJt62EaIc31+NHqnhcK
k73Mam67VtMzvWtZK9mo49cSC/nZwA0BeizXzXZfKxlFrcWawI4gocro/E9cJuT0ySNeiya+pnFb
TmGTgShx2oYn/UBRpXiWDRf9/F8UbVFaIofgf5BRe5/b0emPj0fbwhlpTu8F3HuZ93uAh/xUeTmq
ne911e5P1VHYeaoYGpBIDkjiDT4Zg7iGeUZ/mU+kUb/tHTpeFKEMGHxR7ea06OjNxkK/UWrhOhyq
4FemIqVqk/WqpnDioScwFnk5Tb4HfEYfhPPGeZVKEYPW6DRGkjQvmwIoHHkNbAiJgKNkwo9xT4z9
0ApDRsGvjVNWvdaJDbCXwxCYAtC+ZWKspgvT+rzvIR6LsjfTQSZkZh5Nge5m7qVGsgIirrbAKDQQ
Ll+gGrMyYZAHjSCvE5HPAMLXWmTdqYoTHha4xG8XQPzEcI1jnjPtGIrVfk+qCUtbJ2j6tzEMbChx
NPR+YzB5SOPMA3KcS9u17eazBZpZqEwDuAfBK0RTsGSvpvbBFr2fE2zUbaNCgC8bat4hD09zc2Jx
lKzVPD5JHifHfWN3QQmQpww5hxGCZaeOkFePO2YkriBkOyMToAdKFGwCmOUra8ztUhTxaCN07r1t
SpCjxWvKADH1cJyyFFeoMI2+B+3+a5PrmPeKQoRAUg+K8jgDh6sNvFkfQkEFeX+A34gfTP7tvU5T
6T54LIJE4wX8DmhyuQ+fRxSayOSG81mwe0BMaAOt2b51fZ3TKL6dpSrP9NuUOsoToD8+3tphzdDG
xL9OyVZ5u1grBmsn95T1a+T/4ZCRxBFqVvKAW1bcGfn3fUCMlHCB0/pSkcvvExei3tfidClvPKtS
EKTWt8D2XOQPzGEZLxU3LX/bkt5goQ/+6e1v/iM+PQ2nT4FkH8mA0DnHuSYdguQ8qAwWSz45Dx34
FaaPHY4/uvvkAtB9a0Ns0xpJfvaux8C6LWDeG674TSWJdTR33loC4fYnFecOUOgMs0kGFMe01gsC
WWUPOlAQsRD4rNabCNjJX2fKT6dYZf+2lbq74Qcp4jmUv242xJtSZ5kvMDm6F3lq2/lqu5zKcErr
UulmtuXRPwM1p+/1qNxOTw7qLXJMIoQGhY4/cYagtfZjkUaR9U4BgDppQyEEccS+tXXdnzieb1Ig
1w2M68CJJYZXHcFofkj+GMb/ymkbUpAJ0xnv4YvikWTMcdwY1uWpbub8nRUPal1Um9pJrT0NQvpj
MVXbUN7USx1KiQcEF4euSrOq0hyxTr6ojAFFKqtidgygcvUC8QisRTkiwI8yH5VHr2v6SRmKXV4g
NISakD5//Is4QGNcInqnAlzq2mWfsz6tc4ktT5lly3zXZYwC180UpQaZNNUEN2D1LdSJ7eBVk53b
Ly7p52vMYhvCocFq3UuBDfaE+CRG3TMTAKlzjnWiydyCPHI+MSKHDULTLssO4L2Hac3SgRLE+84X
A0yYaohRIbv6gq1kc1Zqb5KvawdntIT27gtvb9DNYqxvHaKCebsJjNYvNDR99k4rZxUUi1ltnCCS
8EbED37j8xIeAmLR/Ij3XqNCrDDYjszPnBjFtN16SYL7o2TUn+I4zKEpi4vt7RV/O9mOcdd/DkHP
E4IhibJ2apAn6XQDkcdX7dPs9Lh6z7mKVxzFLjqFUASkY445+/QF4Al0Bf2PL/WpAGJGOYlAk0BR
lVztGEpEwpl02oCtUgJsrkAdZ5rK6UU4nw1MLN05tUVg6FCPZIXXwPy33eGQpMcbLdO6HJmOrG64
EqBCRtWGDX9EZbYPQ1ZK27zFBqUnlukM/s+U83BbQwcZdSg5xFWii4JOn+RzQgyJFpuQYrTyy9sm
U9PhfIUqTNjbznnahgUamJcHUIBjzqfRoETRrvUVXudzaR2RSdCF6QBxsLH86qbOhS87hp9/MlDr
L4R15wc9DPXKwtCEXZzUgWl+CqfKorvuFj6mVzkKcRQfA380fQ2fcPq0/shqWmIMqHesXkMhr+61
5p5UaTFOt6GyYnuBlqsD7gK/S/bTfljjniJmDmbmkwx9wEqzH8TzhptcqbaIS+esKi/MxCw6qQ/v
L8BWB25IqZtbnSFrVuL+Wa/CkFI1b2nNF2vzJOECA27fVUAk7lgIp28DtRDVjFL/KdS+l85gAWdG
HOHS9aByhIQRpcswgONci5/sL54FYUIzs7nOsZFkNTvNhvknsi4zAn9jQUY3OP84ZknfFKooDROD
6rAzXBMgyoyRzow6hRtYgeqGgAy1oGVK/DP1Zy+yg+D2giLxO563fX9ysn7Icp82P5JAEEETGUy0
wBaf6KD/FXxG80EOvHEXPdfsSFEc6pAcaI2Q6zIqYF1+j4zydDl2hk36AemIQw0ZQyG4lF5hL9jV
/ZJH+BsokRcxcR98+OxGvNwltFnO3piO6r7GpCgEz5fgq3bcFl6MKmPwTK+ljS5z/scGn3Ib/ugh
8Wly8gsB+MpSqePxXrn4SJjiTtsApkzkVsmPDmS+J3cr4O2XNWxAb9KhWzhgpIWktyGuW88wgksV
8sG5/inng0U3CKr3JwimXECvedfakHgGfcBqFD688xSvzYHy/4hmZM1BC3pihhEIYVTOKn0997Y2
d83+kHWgC4KqeaMeidxnArVv5YUvd3Wg2PIJpbtanFrE8713ypcfpoVZlmmKmJFz18b5EK4KLAoR
McLdwetW9Lq4IF2DR4OAkmOy3IcJnDA8kuW9MLf+qjBjKPkvZZ8wwyJWKi5Yfk6nIBGcQI5uOSFG
+2AjhTTYwIyNRuFgx1Ohtj5ZfnQiNSukAwvLnfH1CMhp01v49fyRlJO4wdIa8L5rOjoAdozGosXG
vIypI7/NmW+R7XkD7NA8kVTisLXNCz8yG1C3n6ynqdFxnLFrfQIaMplAJ4zdfxbvi2/13jjEaJLU
9tK2/m6CZo5XyBpF7Fl31Ygcmmpm2cjssAq1b5OdJdt2Os5TtPXfHvBcUs4b+1/sPz3Sh2D/lj9q
oJZ01DovQm4iPLGJ84580NFtWjM8XzhlfeNrYoOExy0zAwiPnCT1OkroVP7K5NVgx2tXjK2DmjPg
6eJJ8ZYRbuVNDILjHJabqMok7/g9aOurzD1UydCxSDQsgGJHLtWgarwT2pf9zisApyOvTQhYVWkt
3rj1pmYN9phHalznSB6e/SphmPebeGNhcnuIYYFD9dkfpr8CIg8qCyMqZfUVmsP4Z7lItDpDs5ox
bITF64sgbbRMTge0tW4ccehflwdEsYoCGkptCCN6uqtBl4/7nJJS1doLveRJnGbzYwyjRwNtODu/
z3UUT/6PJmtfo9ahGSb8Wms3VbZLg+gVOzW6B40C0kiyAYN3WPr6L8+t/TsWvvg08YAl30KjZI2J
n0NPL1ZDQG98vsuo30vrRlhQDiW7x1a3C3ibKz1FzfURaQsb7xLB4coRgqFwyKNnhssZlajE6uBF
AaplyN86LzGjSyp6uvVjxh/fM7++z7KQ34zgXcnQxDn4f5Nk+2DJEV2oPDHhlKQnHjIFnsAM969T
NAeagni/tLyssi3BAPafbJ+7GRk2OGljrPt33+LgxSEJCKKtdLbPXSHKgnV4RCpFfSUavEpx4rTD
08ti95H8aXQ/gmSYhVIjAn9XnoA8FaX2rNftVc66YgD32MKdX+TktomnjNmYkBmjtwzUcD952OGk
k/BHOoQDDrPvQOpvq1IAtTReBSu2ykXrG/YalQ2/jJLJ+v6duIHE8XsVs4j+SE9VtUbKLCPifhB7
9MGOnMTTyDB6R/X3BGCGtRaqHOMIf+hCWQc41mEHzgXncGAM2Iv9rIHrJDCO6kSw/p9hq7kK6+Ao
meHBlYdb/YqQXzdKCSSmCGtvVj+dvGX7eYKzKxT4aGwtBf0nIGhL754mhHKyvDiBcHLL+qAN4Rly
i7eBy4S18T98AAmgqnQPaeFjchk65qi7t1hhjIo1Spyw7XTfrM/Sfe5gAYq8KXIqQxxne+l65tek
VCs8auJXqOCx76lW9UK9vfyO69ixSzuLnaTboywfb0EhdskDakJ3i8yWEizDoOLJC5oIuceWzwXZ
TOiwgc+7yVbkIns0HmvvuPmwIj39iNt7p5rPTuV4px1RyEfHDIfKECZ2TDhe2HjZbY2N97btRIrQ
Gj68yv7nud9daDlHybMKpC3aN+dq1XSIWBtNZKUrcY74mrGQd6Fcl6qez8bPik1Ko4td9Cw+qnKG
rIcLsIwEJg9L5JBWSUCr+32duloy+0zn6KaF0IfTQmBqacWq+6AZhh58qMOamqzJBu2FWPSwUeHX
KJvqGM/izzdwSj30PUdiGM/UrKw4ojUs+l6dmCVFkmOnY8LMYa6Pne9QGRfk8qRFVuqN6+Xg72c1
K+2k6nk8vM6PBj7C1HefJ86WJ+i+goIpzsYSph8QaM3Atsx/iiw2wHMjgViL9dd526ol7qDLKXYJ
TAh59vfSSIN4I9/oQqUEXcs0Ftm85fJEgWyA5eMZ9FDSRz6p0XZuJur6DIYxBzHWMXsKxh5O/Ide
y9ImX0o3cWpAw30JqyPjGLuZfdEroSk6ejgfvizyBVtSvNTJtf+rMLV1hSjALJHJ1bwaaFg8s63s
fbh42vyrg5yJTmUtavSOOwQV0TKOEeRJ9YpjkLbQwy1/uHVYdD2k9Hk8Q/mOLXTClYUADQOWrMf6
IikSmsjF2ozLT6ZayVHCafJUeuPo9IOzoJ/IEoW+4vCNrILlULTtp9gwViXLfHqFhUD+aewtehv1
64qFG/a2OJjg5fxuoAfL6gvgpexYnIWuqyLaT159Aas7Gnk4q7qqDSY2cjtIw+6/4igp4sN/8jg3
CelK3rw31U+XXon86ptNdMMUk2E1uR2i98LP9sF0vnnj873/aKduhjcGvv84DkaCOgaddka1nJiv
EDz3kKmr7vzfxDJsPVMzTZlulLEMKWpnQMFyLT9Cop39qsOVjGSn56yVNBtv86BecbhlQIIio6LO
XOM8XRZ0cqexKe2ktDaBfDHV6JtZshEPRm/2eklzZ5AcYtgABjP0SJApaWpn0Z4hYzE8vuPha2dc
rEKK3OvH0Pk3LO7rZL9DkKEOTWSiIYoZYQ7ifm8Y77FiQ7AuZwkgz5TnqaBfluhIqtrUepy5sObh
uuoa3dM9Ur0EllNVfCLGGhC+G/dveirdf+/NU8hZRW0RFwuyQB5xo4yGEz1PsY6O57BQnUjdoUUH
Dw4a2lnMj7VixmEDOYtVxfnFe7SWMkDSjhjxE07dooQskP8STwciWl/7S9zVBX6nHJqX4UvVZr5i
iXD1zs+1/IzTZVyZutj2Z68eFNRZtQ1G/OwuHStAivHSy8Uefec+Xt/PvL01LY7glOe3bVli57Vm
IDH2hDjDEd9ywOKmxRmOnO+QPKgK4mpql3vDBq57GO16WYXuPLzW0CtNa6GhgEh7L1oNGJD0thaz
tXDfDzYXKfvY48p/DELju4hjhEY9lDq4056VDKS2KN5sziAUmeu0Lx1Yr40+6D4gtEOZrwSzP8uz
gaqovrlzXKpY641Mtcm4fOKMw9ulYn4V59A3pYflI72zpYs3r9ZeyVtUg5RY9anHUIwpvePtLlzA
h2JhYK8ufox2j6hFSVRL2pgHAieYzdEREvckJDSYWkeSB29Vz3UoXaKAeYBq2n1Z07ET2wiiCkZt
rUMzti5qPP/0kze/6HYvfuP7LwEjBQlxYUuEKki6cm/8W+tMTLIho57hxcFvxdsHDwq4nM8N8npH
iKpyBhtBzSmDZMx7EV9pDa/U1OHvAWpV4mHRKN6Uw3A059WO7FT7p22ME3ErVr6GuKhU0qC3uLpc
Ji4eM+4JwozZVkZ/mjDL4dYNUesKxG7UsPbGYPiBTPMXCRGheViRbMK8CSHyYvwc8cOjo1s8hnw0
63XhLFLjC3GrSTB5p1NfcCdSODG44c9Lx59Kb0cEyk3bpn5P74iq701Cde9U0YoIkiswrvNN4I5q
Cqitk+LhWeeqk5fXJOE77eBhYe/znkbft8EU+NNE0Dwtlfzdzv1VChIe+zuNv4kdBX7tQVgGGymC
gAlr9372aqtzElEzDgfJTGOOH9gID8j2QygW/Jk0vPZb8spWHYWvF47dRPt8uuzB6scMyXOhFJjN
pydmcfeM7zIXEYXmKSKkL6FTib6YLDIksJk5umJuLRItEuMaj2K3QIjgw+r6ExOIaZt5bVXLygsg
MicTcoCdvR3h2x3oVdnpXuZSK/27YNZUA3m4IG9ePCuDppFjbxB15PRXNrJe9gDKbxKvyS7es3kg
xHo/TWTX66wJ5+9lwXX3QSnJbtlmxVnpZqkvOmzHOq35Y1uZVaUyn8VquTrMaOm07oNxULHT8Lya
FJzKGcEac5+x2AZHElsvtnVNlVuIG/ckGKSFGqLXXDANh7e9nG3OEz10RzS5fHABNjDTQCXfPOOf
QxGEpuaZ460bwOL6L9UxvT5BQg+u1aH2TaOAHrmiEOPmjQ/dscqG+SkOThbl5+FOn3vVefFonraT
p2pzep7iSkmWPELffXrHlr3Yozs1AWfDAczbevN/0FuvHu7eCOHLSjL1S1RVoLFaZGXXKx7zF2AE
4EqmQbFU1XBzGt+F4rIzjfajYXFUOreH54Hl1zZoA7/Wx6guYzPP3tcc9hhfLEFla6aSjtDWBmxs
nB6KRDKapaU/wjzl5djUi8K6MpJabLKudbjV1SEYmGHedACV/P+uiIjzgRD4veRmZqywbrgeftpp
P9ibrWq083qgMlIk1WZeHKBnUASGE3CCp6s18+QSm2ezVesxFlbnRRCh9NviMuPQOdKAy5TfbAH/
uzqwCcJDyeK8oNhUKjFG/Oy0puAh3v6JT2VPWdKJ25mMocb6bbJnLnnNMinFHXKba+xuGXMXCgUS
zZoNFh/vdsRzGba25VGJU6DDGkxrewm7hgp2v7HwMB4bRM/xu/oQ5DvozwysPVJqeizIHsaxCUIk
NlKevJuu/Cyt4iRYNakiiqpexHgxZEyMMeEwYwno0gXmEpLnhyLRaX3Ji1hbmXwSdl4u/6RpxL4Y
F/76vhblkDQQ7NHVlxBcx2Bj9IzOJCp4WmzAMitC9QzcTIKycA6gy2DOk5Hf+RaHH4rjPeCRQX2v
Y5C/70ZdxxY5Hmre30tYnyRHansUv90TY4ZMQ6TozEsGdIN3ZzxVcndSyaVDKJachK4nhc8B+9Qq
NPGsA8WtQ1jNiKKyqHA0fzhCNcrT0B/Q5J8mgXp4tgbrmo53E4HBHfxPGgb1P3wB/DYlhewaeG3C
3iJ/Y6V+6kBSVWUZo5S/cFpnJyByEB7Eog+cp4hVfH7v36zbCNTpXmcN+okOKB1qzhTvK7RdGPfa
/Rgnpn/1/mONOyQ7msFrswIwTvIaCIGal8GhZlsexbNM9fTvOo5nNcl75crJE8IbU/zXtpmefsYH
/wYZkYoBvloNFspL1KjOBAD11MWZB8nAkRB9q1RISN3NHAkQV4NSw7O4m0nJwYtsEkwHrDJAZ1hh
Wrp7O3nmc3Bur+1UKay8ycFinEKvWbY0YDWxeSSXi2ffV+55/qHga6CX6F95JCgnZvpNYyWHeTkN
zSAG6/Lcqi0Qsbg6dRWS4qegrlYmqkF+4kqtLy1lfIGh7oRqEyqsMhZ8hYRmt3iz5+EN80WY+ctL
B4+8XmWbV8NNuTaPQH4GMOHejtJw7vLUyNJn2bRoyOlni/2B/W5IunCGUe78I9nqxa5NHo384P/v
1KO5aZ3cgTD09MY7YdXM7ZSmmUnw/edcvWBFftwUwYBmWLJiwd89f5YaH+eU5fIN8omV2n/Nfz0h
wS+kAkmxoGf1QyylSNcs66GYXfT8sABb95fiLeS6UPr74VJ9oh55GFEflffjo2kxC/Q7d1wyQ/Gu
kBE32++pUkeozxusNnRskQKD1wg6wuP7Aep/6khbUmKLKe05LMUYGj8fJ7xe4shNeqdT6opjLu5k
1CyTP9HXNFtnrVSIJJW4U272RMAa2d5AkjBQMpZt/kecP3V0dsPMSILtQpLSsMxlZf5JhYEH0kb/
EbJQkI5thcc5YQZ3GVve4S4Xi+2/4DComJWIQBzN3vaHd1IPdlaDxWD8cW1WaGm6xcpKEK3gKWuy
waSzpeL1U/TDxDz3L/FonjF9jCizaj25ZIS6P89H8p/ev6qkWcvmu1mV7sIR6T/1mqG6Z+ByI4ij
uTW+bmV8nUpWreAE9Y2GEfRq/J8FOpbqig2gij5K0tISMwPlKbzUcDqQmqoF6kf0oh5akS+sLoSI
Rrt2on+FNm10f/DXi48S2Me8Fj3mxwlYKM032FoHf2SGh80k8mN0b215xrslZlfFtl4uXJBh13Yh
MbFoEeYGIyAzojsa9hzSIgrNTHojwb8ffPzUrG1VsE9YJvUhz+jvSO3Dyjk2oBQ8l0a4sQnZjO62
FLUy2gEyKfbEOnxLC0UKFEfULuICEt18f29DrGrMyDoUYQI/kPwJ8Kc8TBDCfS44Ditm7d/JkfYo
BmrKwc1UWLi2CZaUk+uocU55ozj9xU1Iy3+Cy04PE0tzzTxbdys9YMMsBiCN2+4Nkodvi5Fev/V6
sFo9aBPxCR+mZrZfqptbT6ivNMLNSEAh9sANeeSuNIXFdq9F+yGo07y4mWhBLfc5V798rMEWd2ua
O5dVkswusSw9enlrbu04htSYiCKH3AbWB0I9cPXu7fnZj4hV++MiE0rmCP2ocvpLlQCyO9L0C9cu
nuIdTRUgTWeYZXvKsB4uqI22foY8XGqSsDJDujm68LD+/vkmmguKIRQ44vTKovTdINDdaC3xB7TK
qIngwCjHK7lY9v3DloUosr+K/YBW8YldpI/QUcRH5aBFCXWnmVH3HokH4UAYSWuOsHmZ5J+CHmd9
HKHijRaxysswPgs0U04DhnxpPMgnlgXJBRKH311nrequ8Focp2TlXE0AmMVAUvr62GMjMZDYXoGh
MOTcvC0/YZdq1LKfaAIHzD4IkZPO0SJeKegnAw7pXeeodePHwJ1riHmCtzRcyNa4AE6JhUGUYoQV
WF4iiyRwhGfciNKfbNQ//9fklqLPTzTLJz1Ep2fNvjnoBLS2t84HNPUVMuwlAuQ8we/aX8TLhRSS
idXrn+Nn+KL/nDBJIQjLifkmtakwTJSOcPvRLW6NJV2gcmJZC8/3YEM3D7SF9Z5/wr19UdWS9YxR
YQJl8z3gLf4XDWd97i1hP25WFRM4Lt0stoHlUWV+MB98LP7oJ/hkPci0nVJtpHJk6JYjnmRKnFgf
dyTzyicLUkm7K2oWYShp4sjEcI6mptMT/if5iN1IkQk4/izJYGiDIGJF+09StMFYo/r7VXPpbDVj
7KhFrw5RkqEKiII3SpHPKeUeeVBlOSaJG3QNqpO9rtKLQX2i659hS1L+6gaxh01O5073eKq41wr3
P5Brun0DtizroYj1sEdG6bnxzs/tjml6lY9p6qtagq18gwSCU6Ij9Dxsr5wtBPSY23wUcGQMSScA
aUwck10RPa6VLAYqZjFlufX4kSEBtN2VTTnaPhVTMLpnDcWt4F1HOVNHUiQKib8GOzM2Aj6C252w
4ri2O1ZfNPg/g5+HRfWVgX/tFHR02ta4QGkWHe3dms+Ld3hdqtcdrj2P5m6ZxrGzhe3fvz5lZx2b
D6Ft9O3AQ8l57lttIP/8rXbl7pFh9/tMAEBqdxu0ZBRdFGa5AmPJk9tNxDzDcLkIgXC8mAQk0BCk
HQZ7VE/wHbQsDqzhZWd3zB4NCkFFxuCIomHNuWwH9LmcHCTbr70PJIgCvhMPrNDTv9kO9hTIvHYd
eJBJ7U45GXDBVcwN5F4dv7w9ZwMsqoP74jN1kAZ9IDZvJ25Qc8lx5V2GBF9UxSfBt5CqfAXliQUa
tmOZHL+mzpwOxYvUbjnr10ejmP23YMZfT1ef1bpNsbpmwAeJGeNfzFBZJcaUmsPxO5YFYmaPDCh9
cqKJwUpYZdKzy7Zsn2NLLTna8D0XuyeefLUYgTl5BHocJ3NX3lZrOWT+iSl5VHFAUDzg28SaJjc/
vL50qfzw4ivXKXH03Tr8MOOmxvecS5g54UzkdWEqKRdX6PJGL5YluSXWUlDHgHQdf+R+qLRoltA5
Kg8346aHUtwVjn+kQ5BxuYqku7P2C6sZNRWaF6KGUTpWEalepdcgWDYj2DY46xz/pcmN+CPhUOCC
jlFFDOjkYhrCzLhRfcql34tJhBMsU/su1ZNDqvTpVw/Yp+JJWsWwddL3S6rnh7wuANaXGgWvETkw
AiTOkE9eG50ehDS6u43eKd5HINHW7oq7DOhET45g8zu4G8LS2jaxz2CIMKq9nEuGILlpeVM6jKKo
z8wc/KOQ71b3f/f0utKd5Ydo1+nzpXD0SewvZqKxdeJ/tQF14cJLkqHKyhnU8hFDOWWhL+lL+V1C
i9E/dQKMGx2/prhHK6RkMYrzQX2ThAtZSDehzTB0lXloux6gFvddtORTeNJox/NN/pqutbpxXhUK
Fnep/6HzdFapiZ5zXBXmtBwhomhd6+TB+Joe5VF5SyCU/7jbyMepGKyRsNrpTvAvN+xqWtmF7d2d
wVTL/RwdacBJI4ttnkP6nYgBG7UWetpCVBxBjlEQU90jBKkh8HI0dQ/lSfupXB+rH08NHnDhJWxz
CzsN/lGF9rf4AvmhrqN7MbeYphRovOd5dZ3ljGQf5/fiK2kIODxdUhHCRvog+pOEDi4XzWSDpU+3
rod50Biaw0zFSdXDDXQ1Er7z7eCtKPVduLYIFvLgt29bSV92lFG94xLi55pLp50Da0b4dUeFp5t8
/Yt0GdXDNH7a0R75gKYfeq0MyfKVU1NgWLrK1mMBRBhduEW8sfenRhy8ZgPR0y5EoTZitnd2yeaI
mWIyDazXGEzQqvIxsZvltia74FmxLpUIHXSY8gCSA+kMqRZ1qMuwblql7cD2rqWH3tj++/u/GvDj
5MHEA6GmwUoBy/mMaGmybJVNOMX88VBLj9Zh6mVSTEhNF3QvHupPsQsn5+3zuDiEzh/c33MtBhr2
4JKiIDrSFq4dsaFFOsFCEjEDud0TkyCObThrK9j2crgkRriuPOA+3Hf1rn4e059B7x68A0UQPKMX
CvlL5wtmYR76XhhlRhl+QLNpQ3vaCYatE80E4q/dntXAI5eMDUjVWhNpP0x0HkioaCRNa//rUpbq
tBsEfRi3iD/GO3F4yZ3/FYTe186o4d7nZW5EY/RkqPCJ1klaQpyDOqMSfUE+UJ2DWrwG3F5lcxMb
KWCi+h7adGoqWt9HFzl49eZ8hl2qS3eIooRODa9cscqJof8iB0/12E4Vejpn1ZYJHegGcVEfwzDT
Kf2xjhNioCrBn5D3pGrHjpjkQHyeNWCx3xSObxVFTn54qQG0/DEUqxeTBmCKiO9C7N3Ro3lNpiEP
t8ZlTsT6XCKKoipqGOh3IowDl4XbDJwbb2UECGTYZecUAyrA/0iamhxfM4xG0euvwvLElN/pUtle
3H6AsWSiLmY5hUfxXyWGRt89q9rXnkiTAPXJ1Fl+KKUwvmokjVDYB8vxLVNxECqhdiB47ezdOBFx
gNZ6gXfBHAsB8x4fc2sT7B1X+vU9GOPBFgOpaWDlSDZBdfX+n65aX1iuxZ8zLzmdNO1W5TMXyHJd
7UVeWtxD0Pe2DYly067sYNQBmR+7zIA6/6ydsXL6/4XGrh2AN1Nll+EIlq5Lxlci8h/9ShoEhttH
kHDDKxEVYmuEwfDuJXgT2EFNINK0LBDh46IHxsyZANK92IPVxJQyyP2uJkz8+aE+8BJDyyl7kErA
7DiYqlK0WpcXLRHu1g/vbITzavsZTqP36lo7EkzWXl4oVyIW7IeU961WzbJffFjynxtUv3CPhlZQ
mdUT3JyUAbVWVP22Cqtjrt5P/yLT0q/UWAI9+hoq1HE4S1HongEGv2PBF1kg1IXHkuWi74OQut2N
g/i11xxveo8MfOhn+iRltCBJqphewzsqoZETs9/tdzczj0r8/a+y+Tvceod8fby7Qv9CtBIQCCjE
FsrlxBO+i+oGjO6IFLybi3Y3mU9rjfODb0ocHsQOk9FHZEjyzUYxcgdh7L5obM5GB8nrzX2fGqBC
+f1vSDG67wxurRS3H+M4vPiA54HMH3F13PggCNkIUvRFU7DQsSptaOU1Ie1Ze24NJQrKfXvzIHTp
DwM3mmlYP6JilDIprWCtr9fCmPI5fLnlxpUKpIx3s5Uf8XCTtvLOOwKiHsaC1Z2zKO/W4MK6BdHF
OGDG5jNmbRGmI5ejfsK/wmatSUIQhddrhMEfpdpNN4R/XJfu818JG2w1hq9JU3zITFq/w3MCNEGh
RuvAQWLx8ThuPw8vLedEn4p9vaeBJIS1ADXIEl0MfS34eq0ewG3030lcnDCm56r4VrzNOQBIOkdb
o1ZK3wWQzum86hGKGCSzL+MS0+enYSxVw4H7qDOF9zfM7eR416EIkDka7N5KtvKlY831v24uTsyL
mJECqgW97V02FcUBuk5PA8mhFiLvg0gI2Ih/QaoiMAFRsfZiiuRuxD8Irbybd9NDeYz5enMljPAT
oiCjmbKYugfYlz9rdXC5wWz+IB1UMuJiOUrlixc+2hoIoSR8vBNN+T+aoQhrJ/UaxNQB5iX9xCNb
xMOn5xgc4ydNFC2s3oCcM2H5OhPVmi6e1WoDqU+l0RqxRd5eciMd3Qb8pYdkzXJeTPjB4j0pdUqB
Q+JTH/YK+jrR4/IlAZQ+H6j8BiHhuX5lc2kxLS0Md/jwP994u3hftClBHo6p/n1B6nl3jQqxvlCJ
LUWLvxQwCHfakwj6IgQqkovCLhQ3qBdRqYWsV42oj8BpErYcTVB0llt3vatLMWh+NGzR444b5yBm
nmBxF5PnTxwXC9UUCFwkvwLfSvmKr3PMpKMQAh6KGhKtAyQLmT3zc7NhKkuSAC6vdbZcjKqYNzC2
4P/LJ1gXDTUH1KS+KgjtZdhz3xDc7Ku6xRuLNLmHTR2LmOIaiAky0NLfSiN0zvS1Q7fq1+/P0go/
pM7oLcsK7/lf6hfljvi5jUX5/V3AsbQ+8qmEHnsuK6i3T/hsVrNP2NXyFOv+mFwVz701Znvt8Dld
uW9FsAfB5PUcUsZ69vWZdrfFwiK9qnDuXihMNVdUTTqO2JWpPAcHHkX7DIOQ3S3zG5pWvN0rk2f3
AZaCt4c++YHURh3nfWjb3rrCUqx/qzPX/rgtbiztjhh4xpMyVR8JyqSqlmJIUKbx4FZD9ExA9GF9
IP+M3nmttrS2gkJuwfJmWRRCDepmDK4al1V5yQhReuT8kgrHU0mGSCX4ENSaMc/aHOdX00f63T6U
BYDbTmlcTSxxe6engINW41zsyhkGpLFgT6LS3CSPtfIJ027JjPquoE9GLQJPBui3gFCdEugXE74l
HWAbMConOCZfPgx0yz7xOJOfCUe+mqYOG9d0N47MnNPLt1J6rvABd4PIyoPLOLz9OETf3+S1V8ft
8yfNOXFezi546LnSD+ff1bACAaJvkThqcKD2nxo+OwyhxXutwK+WTFJ6BO+dwLLR+a2vSG5R6ZNL
eqjm5tB8FNT9zQhoNGfvEUF9NKeT4zUtoyHRvFz8ndQNyyi5Ygwh0n7h3i/Pwnr2YzMTT055Ztvk
J2j6DxOQf5uWe/gSgu4dWtgQmbu4O3Tg4HHpXB3/nQ1Yq66D2x9B7BgijYoQ7cTDy6xgVvF/E8G2
sCPOAW7C561GAcjUSevGWbOG/Qyhq7ih0Cr5QF8B3JSeyAhmWsBpCRemcDBqMVBxaRaHNwDtUrZ8
+2f3CPeyR5DosdJpt5ne35/Q1NopZkkTMgPgOBwAhrz7sFPV5Jc68/eeg/+WjIg5d12YiUgYRz3J
a82QMhn6qr9r9sXfh/6QpvLs5ORNtAvaTAORB57iz0IaaznafH/FpFON+D2nmqXXIVFXAPCX1eJ+
1eupx9q5tjF2wOmjZic6/xUxpwYsP80pP/9j+pBrd7LnhKUwbx/GIBkJ2SbtZrB60Sm1OCkvHJ58
4TKb02dvgnyuLxc/DJ7cQPURqAAgFfHghvElPsOW5PP/cNRcmr3kyPt/YHJDLxvzY6av0Gn3vLR4
4GZE2hSYvOHVs96wQYQz9TiZ/y29NLkiXHevOEu1EsnSjOYe4k/ze5VCDO08FFtCmJSz1fjXn8sI
xqWouTtz1T5c+LSF2ypcw5CZO/aItRvaF+IOI89Ku11w0P2lq2jcf6NkQHE+dzD9LvI9hB+TNgBq
PbkVT8yj3h6nCUxAHYFU7a9Vk2a1jZaPOoxFHCT5fdsq+jhB9ZaLF/54xWdvDvm22Yzir0Iy08Qv
+nrQ6tgj/xSWvvt8HNT9IoqM+2cuej/LdhgBxTxh4hsrIIoJNJ8OAxpOB+A+NCTH6WsmibcVOT3i
Ac0eiIvj/BdLpA41FxMOjqxJWHJQFb5SZboqp8nCuQ2ja9C3HGQfKoDGMYaRvz/Ga25nNTGjqAwq
YMr2CFIuh9gOO9+YxsOfoGuQRdAeBrWEMdvbeuAcjqSlunx1gAaJ1Y4ETidTqkF+n+ERYY+eqzRE
DwP2huhGbYCTPwymoDVs42Q6yzgzZfxuaXprdG1G8Qoq3A1rz6EZC0Z4oaKMkUuH2tDXxXvYwEIc
/J+Rt+bE9aJ/BWgA7bu9e1fWg8PnNRaRS60B50UqrNWEydXDYHkYzEnCURTNjQxyNQDdbn3eIkXF
m/fNLUIUvSw5LhLF/pCfH2Gz3WIY+rXdTzF0+3NMHDWyQ+oOLq8mpWE0xZFBJrwK4HKyphjDQIMU
dbU5i03larM7wBAgShkCrqIClaCmEZsqAP1pKD116++5HhMINiusqixqiY3xs+YW+v7B7KL811cE
ZTQlx5rLz4p3ZrYXnieBGY0kUe9zRAKLJGPk7UZRytSJQ/8CVWWq0UH8fwGxDiXzlm5jcG2AvuA7
SffGXw/uJ01M7R4ofwQlbXs/9ULWbSi936FNAgGk3n8EiaCKF+DAF8xljOVXkdQ3e2A9YYEd1rSh
2KrWBXCP1uH4rfTdL5lPowNE/owgMP/io/sWqzpUj2541bX6XD4zbFjtOI1PpSi7hw9KwYvapE7y
mvGgGfKYrJ5AJRUsxRd1LZ9Pn8Aot7Ctt8wFZf7Y3taYR/ahMjuanaZDJgQ9DoYYOUMhK4G5OBDl
NpVErWaJcHQ+gU/gvqUm+RVZBRPQxyVMv7yICRPIuzWG+I7bS67LkedYAvxFuWr/xKcYT1MeFAKO
eLVwvd5Lu45NJHb/n558PqwKCO3ew2N3PLsI5ON4mqLcM+jw4DGl2CNYX+CIPeU0NMF6XJxwlEyk
HS/M0ZOYCz0rWbLfGQL5MdVgnyGNLLCwvxux+rfpy3MaUuSsH4AaFQxQR3eYsgcgitmpIHKHIobh
SiWR5ma+zYXO5z8syC1qbHAGxgWtK1HR48jYr43EkFecwYepSlJed0mm15DskJwKcg0JEKMI7S4K
dxybFxw2i7FMT8BbwnzZX//C4nbethiH4lBkr5uBbDLqOfecU6PqCdFG4PHLeXdGWXqXCr/fNflm
aMA5wOz91whuzJbIdsXMs5iXe94SIiqAItKqnhlOprUGdNrSSu2tto13qKIX4k7PxoXc0UaADg/f
NUD4EMXo5v+wcTID6yhFzfqV6fRxZCW7h6HnhpQgGy6ePwm23pc9PI/LZlQuvZ9oSq8d7P59vxWj
GMrQNqfRQnukbnqHXrs/eVlrICE4CwBcmYrF/5pN8eoCXjfvIl1Abggr+gkbzxIGQNYHhs7t6X0S
YIzwrnrdfrPuE0upawuAORHTcaDW9U0uJasA/cToqbxKZ0yPGRVRVb5beeEVkN1AhuNgNwLuKvgo
OEvJKuXADy0tSigWKU/sLze2kf3qRd8DImZTxFUQPVWwfFEAfJ842E445oz3yekq+dp2v7UIFYFi
T++nso9q8W3kyX1UTgETAQfs32a6Goa/SrGH2zOomOeiU3BGz5plX6kTWolMds4uKYu9WB5oR65d
uwS0MDLqwt5hP9aCSZUqBjfMOJQHdRQ9yIQf35McwEFHRbIygse8zMeyHxYOxgCR4yAmm6VPevJ4
VhlEbhdBwlux8x28Tv2GZaGf80POqO5+/I0D7sYFq9msM85XTRBW24Kfhf8PdQQztnj2Fk5aFR4x
x1Z2jVKNush8H7XO7Db8GgfrkUlhlJABGIcrcUnW43rtAuExEOFZ+USMv5YhmBuSCRQqblh+ok7g
BE5lO/CZvL6/17BFYycU8SBFpydE3gNtVh7G0cqn4/YmJ+VkCeTA0+GM7LWpsfgoe0vnVTcyzoet
4ufvatud7MRRidQHYy2V1FR7qWCkBkv69B982hSmy34i7oJ/VZPl/MWAGuTp6sMIpjEWrVyjNWSN
ZWndY3J4C7VR5an4NdYJrCVNQ3reH46iNUFVv1coO1E/6t5+N5bsfYd+E4xvcwDd0lX8wO1yfMPz
6MoClu3o+YQqcFxRO21HmnQjH0/SR9uXrgLJi1peOkYYlC8i79+T9zZuvapUZxlSc8r458ijpLAS
poSEmqsGer9wqPYEWcUL8+SZ0Cg83TUfy/ZXPLuB3nfqGSOQG5LEZnhDTwIizgp6+TLQEZtjTPCA
tG4J+O8l4tBRMJXdtuuMMjHxpvpyF0SSL/btg3UR2rEfFoPYHIg9m7GJBSX2k9QaQJl+PirmRWvM
u8pAz5naUY27uFM70nXUuNYYStitwhBXgj+CgzVweM7OlaAhFOWZJEOk+wOcMqgH+o9fqSXQVS//
EEAifJtJmz953T2GMfxnRTNBs6izkug/JDekuE5hg7YaH3mH2T0pwG8VFii9wDoifxFpIhbmwlec
is02Vqu5+eVbzH3bQCzEm8rdqeiSaBp0i2ukBQHAk0YYwkGZG8D44H0nHzfp0a0irqy0wdGwa5TG
aqfe9nqUk3iFA48FNL3U82JmghAyaU4UFSP2vhW9o79NKrpsYGWIa5Kk6S6kCRdJRyqDaWK3cwcB
nYiUnyqSmHRkrHkGRn11/ay0hG6IVYMz+U74Tg2cR7A7uXwZiUump3ja9zAWfef/BC1o8lm+Jldc
bEHDPDgI24pPilTIABI3VioMtxr6vOBUoVRjq2vDyrtbUWAadZwK1xtaXgIiR8baqT699kZOBeGy
uA1rMI99hEHB7mdCb44N0dujGRFTqNpONldFwXLcqfp8Dw0F3HmrdeYY/i2mJLBvxGOhWyEj2dRo
QzG2Ix6KHFjHuRdxcypy46P+vAw1H+OWGaKa08Z1467YQ4pqXkJJWlfKgHhVNvYUDl6jkdAm/h8m
tXySt5eIK7kWmMUZ+7gQeCuORhvlBHSiLcnRq8xso4xee7oRIGXQA4A9x4bOTW0HaXd4sJBF991U
ZpLMhrsTfmBXAOZIqdugUK/lsUi1r+KeDsLVvwtTs/Z2nOMHaYFDJIRojnu8mBVw+RMDzr9WQN1b
cujFY4qPsxeR8jLOteHb91xSdxwrpyNzibAJ7rp/UXGMRjXP4K1LLzsb+1I6b0XU/M2hEnfN3q+6
9i25O05TICdM99/qYoBwvg8mwPczaplkp8tYz24KgZ5mOPtUlaINHl2QMIadUUuLxT5aKkEmULE+
2TWWGXWaCsHgVUQnlDdh6IAwgSvMFutEsqbWWPeKrAlboB0ZfKKj8wrAZ1UDHZfO58lWJzvW760s
iq+eaKRTvUUvlLfkhBxZAXOsygq0t8LLOIbhAk+6QWbO9kfjgHkeqoSMcOmMyCePgxPEc5pMs5NP
bdtMiDkMnEOvAQjWLY2Bv75FBZqcXhOIBjd/qqorBNds5sm4VVjB0v+fh9L7PFpvlueVhiCvH1M6
D7RAfJRMEGclaPHeBCjVTV5mMG64l5QOjxxUTCHFTW7Hq+vNfwjW4afGhvQTMRQGwaL0g4czYrgB
JHHc/8zSfvQRgUAQ0rPCqx33u3uNzpJWf/c8ePkMmA+mnsLSlKES1P4fjQrNUzzctqdLH9LRBq1a
Hesw6i+hs3+Hon5w73IiSiJEnbBG7H50Lw0FbGdhgGePezq5nusXjS9G2kakYBOzWx5O19YwxRfI
fsYIzJ2eMKZQuw+KPkcvVhzrvKg0RKPnm5y4SbIKXlfnkOPQB0xQdFxvzyS9hdJfv/MhRKfuaSl1
RKtY+/BPLpPDi3GO8Ddp/xCWh3FfimhGi8GbMOImnEYbQKjJJ2EPgJ21U96702XNOCx9emfjW5E5
aTi7g644uiTPTu7lpitG7Kkv3Brx2NFWLHreMZM5vWV5G7y/9EOhdUXoSpWvSVzEbdb13/tM9D5C
DaPTGeHGw9CK8TkqvcX9w/YuMvIEUcXcnqQ9AZxTE6kbed23zv50AWP9WDPnK+XIv3RZnIW7iImf
5GbBUp2SxH3S/tVbdb4qmBeMu7YLjSVKXRGVf4iNsXNuVES/sEVz0bscAK+Zg6bN7QNShQHRrZtf
27I2uNkn/hS/Nyf8NkTODvMcUkIRtHK1NU/GzjhtD8aqWH7JkZNBZYOLe4bm7VOj3ruIW9mSVps9
T2NlAkmwgLuYTxCxPXkLb9uofyqikDqaYLlQSTe7r1VtQMLJcbTjO/TNIDNFNqa+WirCjsgEsffK
uWhl/uKqMNVHISuiThsfllIIyV3jYZZ7nSJSVrUN1ChFhJU4YBCFIwXpMMUzveZ2kx4bvtdMlnRC
/xjOESOtXDZZQe3bK+8k00MrUlREpMy4AUeJrkDIKDtoCzNI8m4a69nUoPAAzmAEJ+/0b3i//sLm
4W1LUTWqhIX/LQQH2c1ynnhpk+fX0B7nVeI7OUeHHgbcXGA5Hfo3Hm/Atva8JSuaufoEv3m3Ew5M
7cNQayQjawX4+jKxK3SJdJCoIol3gSM6Cs1r52fzb9RnM3geRWKd9vVHsesiEC586bzHxB8vt1pO
nIXPEj05DZZKyuTH0pm6tFYe9wDz9Ui2SqenqfB3MrjaY2su+lgjKhSjkKESCpEvkbubSgtNDY5p
3GeAKH3LH4gWYFt+JaQ8mSH/ddH/vxjQGLKBozEh3RpKlWtxrj8z5ozev+1xy9Cvfk/f7zOHfajw
rXvsi9EKryF+J97+f9SKn1hiQMvlHim3n0n1OT0SQ/hLLmB/p5+tP8CNL9yKaPDLP0GPattGBQ6K
ubrAFuP6kbUKBINtT/iqorsNiRyHlb4mZlcJTCxJNOvSdOAs3StVLTI2CdYcgoTslutwwPVA3Ewv
OccbLNjDcpGR0guuFVxmolBxdWDnoRawuPFEMOnEmXdC/Vkl6cUqKGnE7goeutUqSFIUv1G6myhu
9PTwbefSNUg3OwEkOXCB088YwWosCWLvmB0Eb54uo/UkPUsswkHV8IBl0DpN/2A3Ba3JkpTJlSKI
Y9MnnaZRbVJ3ZNkAJC9/fcpsOxmhxXZqkizhLbwX3g2bj6lk6fqwXowkmkPpgzwUlnBFYL9qbSXY
tQ4ORpX5hhqXJLOGnoyKRRMvSiPvKg6S0Z9vLoEW353V5358jCvT54cQ6qbRF8dIpUF5TqAtletV
VQ53f6lnDdyfRhVf0B4wjgtGlvCTvi/BSNN9npP9I6zg2FuR9nNs/AWMX4/smyoORQW058c9vWmu
tY3YfFAxCXNNEFiLkSCkLZHeSe302VDfiO9gAkjlf+6w51aVjOG7X8XeYbfb6qiAHtETKzLPTYix
iO3ECUHVFa9GaoRcF627IzSpYbK4xhAqehT5CaU+tgSDL7QAA8SlHlX/bYxu4qujm4yXyp8TUf9s
wL5GbeiT3QP2Bk6zOrx0Vh1jYg7E8QCmPB3B3dN8kZASmclZcgx2sFsEefOZaFLmGee47VjmDUCZ
1bpa3rlWNHIl5xLtg6Cy4GxKIiy+9T+IZzesMyqetAG2usLq9Otf+KLjqJn/lCiPlA+sGkF0ZQZH
ckTuosCYXD+1Rb7xxbKMXi6gWhyVkCp5t4rZZvE7UG4LjueDt5KvcIXADwYr7JytqkaLSuMm6yWI
5dA1gdWEY+0AayqjK+qAGDxUG85DglsPK6tEw2WIfdg+U/DllLmYSSnzK+DbJcqTluvj1n9yNR2U
gx7k2xTnFcllzkAOVSdkc1bCSTJMY98hS8PSzbhVsgnqMaFj6qA7egZmDgx2nC+YvL95umq4+GTi
2OmB3FLQqu0T1KMuV/fVTpPdnYOeAas9rhreQNMu2nx/m/GG8Q7u6n+Lmrxvir0FStqxlYnxV9Au
rXl2R8lcbs94bYDYPsDWopPqZb9nKnXbrI2YR/CNn6swlqZBJpLZJHD7VMmtnuCN3ul1MXTH6NLg
KyPKuYeFBAyrE36PbqR1E6Ch7EbBa7wz+D4IMYSVtRSeewulf+XqZ8VtPn49AnG4lR71+gXZzRyd
POXcVtNEQ6UUzmt8wAvQ2sxvrflghJhrr4LxzsFud71kAuZ6CGPxKQoO5sVQcc1NGs8NEVNEeFFB
zpNe/8AhwIPDvFJNRffSnFJYx8eN515JGpPIhgJk0B/gW2UFmQDleBVX1UV+T5PyiNN04f0CJ60t
mhAAY08It8NHJ5cPJBhDeskb8/rVvllAINtirwx2bf6ejrZbQbMcsV8VSLiLdZGlVg68ZXq2OdvE
W8mAKnFxoGb2+dYMZDwNTnVfusLxfg5z+jBMM54m9IjgFYuVKCy008ilA0IbG5FtGPR9hogjVTfV
PqYOfQaTHuecQrsl3i3IriQOlCT7CZDxrKtPHpP885jvvRnTpyCNYeTkYq3sQYvt9eah7tLCqMFM
ACNYfiggSP7eb5MKPg+vo/efGUV+fkv+hpzBOlZTp8P7PcLS7O/pU0YWOiM/GahjvOQo6M6AshWN
RlUI57+YphssI6iX72U+uZkna3rOgJ8em1e5YzYZFDXjWQh8LbK496b0Oz81OMTSCWSSUxwNoYqQ
9L5m8eaMCt49dHbEtq/rqNnF8s6cVOAdaKp8cTX1OqkSt1AITukzFCk2ZVDK8EQQcr8N+/LJ3jnc
GRDSFCnsSVHemJMCn5RnGySRrQtffxvkbcwvelCX033dJ1MRLY9bP3UJDCLGnQZMQyiqtbSRd9yN
SzTy1bzLhNAXJtnGCGBJOIl0ao2tckjXI0qi0mWylmRsyhkKcUE3sh/4uFJZH0dcuf4f45QUG73/
fZ9K0GgtKbjzro4giPv04kFD3v16sCVGKT2eher8Ikqh/a0v89Adg0oVgTh1QtvDO/4lxr54s3fx
9EjVOrcCeOOd17DdFP8NPHeV4V/QoeaXJ40nFHzoCgwqcZ4yo/9uZq7GO25oIZjIsZ6sjCJw4ahw
1vjR/9/X6l9ia7YOBydLtLxMTcS4dD0LQnX3d0XdhucrsZzwv+jzfMkUQ2qJNaJuTgM+eqCubBcn
DaAPYt4nE5Scd8Pd1hko++XAB57AP8If3nQKlVJuHvlj9j+esLxJHfYpktOocl/lLaP006p5mUMW
B20fUxTJpdPOvnkw7s7ojTlD66AiNZ+hWlBsSRRlSIFM8bEpdvBrpqUvIPHdQGxyvE9KCYtVUPfQ
9shSzHj0SHnIWn3tsG1ZrJVx6fRaQUdiRdpsLvXR9UHMpWgBLonI3Ls8y2bWkOiHglJGu5lEW9FB
DU9Qbgl1PGDSZnR/whioohIsV3KwqLq2MBFECp/QZiJNd/+2t1CnNdO2lGppgXEbOvHJ1A/M0aMV
Ie0z/+KKfUZCuHV7/6c7tKHp99zw3/HoSEVpAYFr1eVD0g9NVgBiXS4qafMAnO8jyvXuO8Jk7XZZ
DxpPdwD3a7C1wrnDfstGnyVIvY9d+n59XdcGPmeSbVmC8km/AJlJ+O17xNsLjUTmoTR+2MDrtifV
myezb3M8yFX7hn4/FzDtvWZLqR16syfWrpll1uANyhSNweewEbBE2D1+umrdC628sgMTmunoEl2/
ePrxf20h/unhZsPJAkutHEPG2EIUHKU6wK1wsxTeCigc9vlRmGVZY0/Qj+op9WP2DoIv3jaSGzP/
BbaT/7EBwrdsGHCBzIeMQyPREchU9CQrNZYUibFQo9utdW72+4VxhwSd07LLtlMoPagmrpz8PVcO
G96WQSlsLo7tNoXw08OgcxAVM6C2cTJXUfnmRoLxKzP/vcWFGxIC1gqpGHUFueYmxDPzqPuh+QCA
YDC2e/gxzpJ+22Bku02rA41RPIctLYgd7kuwP2gEPp6mIMlVrjzelYHkE9JTHDt95M8cCQoetWcO
Cf3g2jhcbsWZcV1tJUjtb6rpLTDOSa7oal8H6yqhogqj2NydvF9UAWgFus5IJch9bqiCXI2QZhcN
ZJx5UV9vzA3yX1zxCq5Ha4faS1FN9mlg3O5t7xHu5xe4zfSU4uv/w/7XTbxLkFyuqUWqIbG90mVB
tBjCtYaQ/Zfx//kM2VACvS8ZtTTuDFFiWKrUyhb+E/aS6UUZSAJ4jguDLi9QEqsezkOePNmRqWyS
JC4ht+0DkADwiT2XezuAYwKHqGMevpe1fs4FaUcwfHGlF2Ym90AEV962J2pAS3lLVCdf4BVyXXGa
LGhNDzxSAfVDguzKH5jZLge1OVN4+HtVhPztdirn89FUMcnsiBZDDJQ6Zm0ybys3vz+BfPA1h7C6
oF5Gce+nbFMq8wLskGzMrjd9HcgGKRNK1k1AW17L7kejjc2RJf8PAr6Ca2CQ8fd4gKCgG0P1xyvb
wxoArx3Lij/em2H9D0guyIFA86KOPTQgFC4hjXZrQSpUQqq2xF3FrzYv4RMmDxKy8qcpD5LUj8ds
elDCOPwUauZjdyBdwEzehevANEX39RnIBVSlz1CAJq19RjDEcGBVHUih9HvW3T3R7QxFLgyCWtC8
QIpiGPirz6U8dnf9i0TS25Zx8R+d0Jhwp+8Xv7njeTsCKVfSI13uvNAaN7JAf8ZSfs6EipW+ge6R
tvqo274feMnZz4sD81wQxtohswxgfn2+6F3M+aDoHIxQKUb7by20TucRL3rNtUhjjGPMHbFSxhRv
Ku86sR8P8lfBxjLzVrYTlisxFdQ4V8ENVzvktDqO8hsav7RzyGaEUS+5NI17xCdPpTFDhXV+XNjj
q0G4020dxDYg1dhMgdXLlGrNYODa2F+R+dgE8SDTmjm5zHglgyF07aGmeB3kA3udkGH+UCPOJ7H7
kDEScQ684FgbatcIvRfeeGK57reAuRQ1ufSx1G4qvyfnjhwdnDM73gQ8UgbPn3/SjWRjJeO57IKs
bUlTbMlviK62igDjTVpiv7OPcHOPAajvoYWKX0oL/yeWGPdGpvmwf/Qn1XrKkPP26W/UJfDRiKaf
ZqmF/xdwaX4EdB4PPEccZtZA/qpbN0Z5PdYfZApd8E4N6C9Pc3mvPvXCqDbk+7upU72Wm+rdmqV2
v9sHoNUXvi+d3gV1SiyEpkPzNY1gQH0gNV06NYJ+jUpc6tKCNo637ibtdjEXEH9MQNEEp/CheiY4
/6E5xVNkU2oRmLlgSbR8Qhx3qCEIVsKiltHI0Tpnq1qXWU8g8NVvrSd7F7H3UvVxShjIOekSXNMq
4ADea5+lZKdR8LLT+k0VMBRRyO6bMWo0ZXrPdc4VUKqSADEXiEtpcGXkCNr1Tatz0xLDu0Iff/Kq
kCTyZo3JNf/p0wJw2bOpVcwycrDBU/qtWslAl4rTC1EL9S2fnpw7jaNOQbIScV5kr0Czwp2f1dl/
Opz+DpwfRzcwj3oualjt/3mWxlXTmSCnNTTyF+leNnOEIZq/kHIt4DHVKE5HiG+LgosGVbLgkWNw
IBz/EhQarIgBAPX4tvAX+eWaNSYGQo6nV1Cf3h9WEOMWUED+qbeyEepIWanTwrOmiXatpxlWaAWe
CC3Sw4ye6r4iTlgEFcLXcv5mAbYb93VhemMaYU6BCgsaZLjRylib8qzyTNslDPwwKt0Bj5IyxBVc
++/xVLUw8kqViKHBS2vsyUMm3IImlX2OX10pXgmWo5kIfIjHhBqxzP5aeEe/eRdOIbVLNfHXdjPQ
tuuMbwPXxR/kR4075WhKQdMr9OS0I/NkI0okHBDnY6hLprITT/T7gV0Ir8SCWF5JSXDA3pZCuo7W
ckSF6RLjIYxgA0ktIVP/LLE4uFLqpXft9KOTQ7lFyzCgUAA27FeOBxxrXA1tXNSi1SS1Xi4XBXi+
P5u5RzQy5hR8ks3SyG2vBr5E9V+ooZZgMGSGjP3daQYwMESQTB+6/xPgEllGydI/k42Fa8+5UZML
1X5vIWlJB5Nq8UH7irUnuZi9ax0OJy4/k79ow21LsmXJMbqXYRRao3ReQRqo3vJzjoG/+bbj3Mub
eJGbvGmlGg5Z5C+yt1COendRXn3S7h64HxxGQYoNMPWKFsU1HBIVXNZgExtR7OwFpIQ4PuPjuvg7
iNJBV9ofhsi1n15nBMY84w3IE58Xzm+5kEAAkFeO9F+slmjRbDzGXH6ZuSzLRwjJzl2jtbq/ep7w
auOYTtb/LQn0KFS6PZq7MJoRB8FTu3T8+Oxp9SmeukquxEg5BLAL6prG2zgdSmh1nXu5Kt+xQ8Af
NFbKB26kl5u6cW2f+BAph8civdPfpdvL/EPIH8MdW41XXAkZHoYYF9OoPfZ2/oZB1rN3dEKDfWMM
utgERJ4UaRDs+YrgzISJshWFpAPOcElo69P+XPT/qDatZPnpQU0PuxbvWEGb3lsA2+Y+QTd+zH/2
yXhNF5xlmYDrJxwgpoaTHZTPM8cKft0A4NcDsjeCtAqv2oZuFE/9qYCoY++CMGh0TRDM7S353GgR
p6FDVk8x/iYCBTMmuyTBSEhenTU3oy1BpTUB64NXkpSKFqRL6EHtA/wvj5iJ9mDRmKVgNhcteerU
IFfSRjnKAwsvnCKt7YF3ebxsfBoK9ELNwqvVC16uvIpMg3pptEBpDT0ZMkxe4ETGuj5jswicF2Er
tmte3pKm24HWbIQL9pymj6suSLeT54HqVrl7jO2f9Esys5qS9N7gMLomttXwKYCVsD8Wft00D6ap
KHUq0X5oeC8KhP9QMDKEMQmzfZoMfqFl+xkX6W9PUakyr6HkXCfNP73tHLdOwU65V3cp+CHl043m
LOGY7/F6R653ZogFMbhriGGH9Pw0yYTihICbcZBoi7lUi6k7VD4/dZIgsCk6zC1A2MpP5Siu1vPZ
RHY+Esqyk+AsMtZJ8y/0xpy+FdF1PrJLNkTdZniotINiXPLWvKGjRhEgGRXMKUeMEn3kO3jbDTJW
aWiYXLnYWuLBJ96DM5C0lxbIZLarxIgm0DFb7Ips1baa7xnSQ/VvesOTN+rIMG/I5gK+mmM2Zw0c
7dYFOVMOe2S7VMpMkxawQCyaL2tRzJ+7+Ltk/Fb/25mFDZMN9HpfwvWifwE563cAGFFe/zZ+4/Rp
kQugm4p2XgbYTMELq9vsbFbW8Qmy/nvQS66yivtRS5bJf6xcQQiI8f86HU5m0IS8CSaRsA4PgWoh
hGBiD7P1NG3rHHR/b7erQxjcGy0U+S2kDGBPAoqqrGicjQe4Y/pij0cXonZxwnPagK5cAHp4Vn6P
qYHzwK92OmjFcSXO/6kNbCbLROxNu8CXvGvT2cWUQxy6Yk8n7LomF1CAYpFINRTAI6+NSSrTqCzL
5draK11+hcbsuWJ8sL9rTSUanrUNCLW0kYA9gtNI3RUg+kRG5gs3P63P+2gL0I1YgYWRsY0V8eeB
Qhs1LHtusBJj82wedMTyVHLcOga2flC/HJVMpGklj9jaFfm0IVI/V6RjO1P9ivq3kLXjhn8EaxGL
krlboWcMLQ6h8HQeKwfu6BhbK1CQfaO6amzAbyEKvHfWCqQdu3x9yGejb+aoUSaFUF7zB+7ybazN
rqZlULDXKcPc9/Na7hLrSdXE2FDDd7ZMYmgYVS6qzXlmWbFsLcKsFmCnWnZqDy9GESYQSo7j6TG9
KkqGvTBYu3QC4AXITELHWkqRTpxIDbn804unyg7NCLtao7sIbQnrlWnZEESkpTW/FVb4AyLyIW9T
AdLs6AqQ/VeXeQY/Yav4C43KbaovXqCjxcVqrLgPZhUsjj0e/iQqD9M8jV2Rp19IYXhvLTj1CoB+
ewc21k1GSoI3GDPIWFjH1Spn3+7lxxOCNWhTUyvrHJ014W/ra585+Iu6tYHi3sbWrYINiTglaY2N
fVo1gJdNRoDDdV8P2pET2Lv6wUctnoaGVB31lm76qhBMvU6tN/R5sDJapUQS5UVNWf+UJr+bKzHa
srwwS4LVZ0yFLYlfNBqvl3XgSvk/GOBEhT0KnjrA9T1jPERfKJdQaWeUDstPaZecDO5KBlVx+LQC
efio/XR5Nk8wl4RMkoRYB41bxb/TjzgiHPb3PG8x34kxB6p4EFxAxThIIJVb+4cGgPrBVjtlT5EE
ZGsuVMoCt2kqS3fKXEibRI/EV6Zk0u//vxUQOvIcb2JVRrKWxji6q5SksqOIg32ZljX2f3oGiyt8
5WrakzWqw12aGTHZEDG0nTmYetawNHshwABJpq7PQkiQOwP2MnE/hh33+ppEnx1ypJLEt9jco7ff
tizKHRq9BsFV43LE+JTPWfkSmWxNJc3L2KX+6QD0IQkd/be4eBlFA1hjhmynspyHQ7nYinWukEb4
LRypPYBFXB60/xMDJc9dOMvEC4ES836qVaTgip4AWdTHK8a3cIhzdJZwg/NKd/ttad292xv9NFxt
7It4AXBlfma8TLLNFDmqJNRro4Lcp+yG7GYAoNZwiyCV/g9/jP+jMHNAFVBaXKFpYPL1QUVh4qhi
UCToJcMhqfxuGeEJsko21iPG6N+yO3xaGOI7BLx/NHD+X8KJoQlreWcHhIeBkeiKMCXdE5Z3koOn
qZ//+eVCE4HKy9gDGc6wItNDbdVGjAKSKU0Ddww3aLoPN656aIImfTcXdfOWQG51O4VwA+ad4F5u
2tFK+NzAKG4odcL0mPfj0IXae/TDFeztLzJtdpaa6iFvg7tJnehaoUMgkQHJ7vsQrRTfJVo+PlCl
UnQzVUuB/+B8QPA1G/O69t9qgngfeVl5WwVjU7iBvMVipqbnxNoJUNhSANNT09PQO8y84ZTsdaJ9
oXo26kfpZECiUeSJBcsIEFUUriwX/XTj2skq8VTa2wSoFA9IabpnpVrKtIKkhFNQjS+CgEBnWDDc
dIEerxKKvDj2A1dVYV8Ehp6o4oE6rFmVpT4iT7x9JJvbMHuEwb9L5szBlXs/27aMgtWLUUdMMrrY
ohqwFACIkKMZQmlpHksS+Mau4uT7wJw6hxAXV1aX8PpS9cYzNiW3dk5zkQr/Z9ujS7KXJkoRBF2V
k/XRJX34ddXpnk9FlOCEUap5WuSvSvBB/hioeDpYobBi/o8NhtgVjpoffcLNisY+6veRYiy/o0BL
k+jl7GVEsk4Xs2Aj3pn5shaHPhPl1ZItbbK3H1DbcO6BZpefutcpMEb1B48h040Q3jzf65GDmF7o
N70gujTMfYHuu6F4r3UqU6Jg9xd83j8nSkfzucuzbgWtlEOzRht4BDmoZ9VXERHTw8cPhWK/mB67
bPQEpTtR+uiz5xqm1sf4vZVdfSzaAzK0VUmRbdCXdd7Z31nWlRWRz4EcZ+6y0oThSWW1PJoYL7tt
+IpbfDI7PfGpPkWXI12CGsqh8dKSTFZ52ctElG4mYk3Sbj4M23i38PzDHU7MWP+jeEcrE38XUqqX
gQjUGE5SRfUMmi/PCskttmbPb4JmPDDKHRkv/TehSAXNm7MWTE+KVafZQhPhJLw1wZJJbY5XfM2S
Bm/gIgiNTbMI4LZUmpyfYMGTvXusoAjKmdgEFNpQ4Uoexmm4L0obQ2Q8fS9cLAptIh5P2ogXQyLI
8vCfNWwCiIzQnhYpM+W+/zapoBBa3ZwPCTbgniOOaeJB/KLzHktkcd9Ucmtqi/OHy11DWhPbleIN
WAvfHh8ltV1LEN+7+ia03o0c/mP8RifP12cIAIXD22xrS5s1EikZpov8+nE2TJWtYLhbyBwtrEWE
9fPsKDcYKmgE4oPvWpNH2ywkkEhcTT+Xaq//CoO4Ur2TPQ3TTVfeQ39iHZSfLrAKr10F68ATr5vI
B1R+Mp9CrvxE1PTx9G4ACW7472QCBpSEmeE64GxXqZo2fcKvB6Tk8BGIrUJbhoZeaFgVC0+zHlOw
gqhSYKOTz/wxjmicBUe9jRiqARUcT3MTJ2worsq9O8C8XnDaMHgbKKKXqePnV91bDxsQvAzhWTg6
9+8MzJe3B+27KG3ccGOfHMCxIlFQmjr+iS6n5xTDr4lQz6Mtb6YEmThNWz/NOyepGJ7qWqDngcqj
Es66jZ0rrTkG71Pzno3+A97IIea32qfsWaCcm43EdMVVxfCdy5YcuYwjTgkXxiA0EPjPw6UXIzMy
y6aNGNa2JaNriPd7pEIW1wjkroebl80TJHtcX7NkhGwYt2IREvfVH5LFYo6N6JZ9mmUXRFqaYbuz
Y8EmMNdhYYIe+eTfyQpKUt5XCMRR//S3VhxzLfqqD0TZB7IYfjeCq977scUvCWrcNOyG0iAPW1xM
wHkN7aY8uwl43bPNnF6FTy3IxclXxT5se72JccIpCazqxDDBlMIf5DcU1qhA93Di1SZZoasUaPDn
e00d96oSvKJ0mXQB3v81c0XCWP9NpirccpKoXEZfeFmcREXyu/8lBYar4MQsL49Em6Cf5vnl46T+
ysWCEtDqYvWpOVSMYndCFlE/q5zPWwAuqQgp8gnjscWpyH/5UxL57RnDt5GYTwXVhbEOCg9iHbLD
pkp2Dg0gUQnmF5nwudWhiAkOTGA5zCwrDzD+6oSZXLYlRMKBAryDQXF+kntlKn0H3cYLNJDYwmvB
jXM3MEFMadNPnfiPlpPHSdwzppU5GEx5eG6rFZbcAUft755qUvdyps+e3YIxuf313abzc0R5ZV/4
fU75gqvQDIu1DY0RyWS47wG8F5eRoAnLWWRO+iugyOx3GHl1aW+V10UYvcC2igbzwAP8F+u3zqDg
K+XklPHhTlz4Mivl02qqO67wS8Gfyf8Q1DQmPUD1tqR0Sh+No7RZndd/IEjgdB/HEOs+c6/RIfTA
c7fYI53uqz5NrrdS1URhmlBLB1G4n0UKKOJoxOxOAm+ltN6sPf+/FKd6Nmr2BM8PGhcDkT97vqtu
miDYpE3eqUEx1dmYE1JTC65hQzOX4/ohn0A0wVkr7Aqb/rO40olT6NbsLEsBqGVjdOC4WaLxB91y
bZ4IdmL/qbA3DRf1iMdxZCA6x/jhcXqmVfvz/htoSsIRxWoxQhX2aXgtAq3Vbtil4zMGI56lw68Q
eobMWlzRJ5+H8azRmTqu7OcyfBY95LDNpuQ57zUqZtVc+IMCyBRjeqJE3uxVJ/rSBWVYBhzlFQCS
GBOBqowfy74SAiiC/j1lQZ8gc07lVUZXbnOts4/IZ1LhvZ3U3BrN4wXNlOqUk2iX2XBM65GFu6gr
Vox6DpynOi9a47aAbFQMEG/+FGGtdnfU2hOF4SGyjF2juwNw46y8LT6f62RDLOdjglJEy5gTwMkJ
JIDUiT6gkFR3o12j0572H36dfllFg4bD+huBTPuGEBxLoqxLPVtUkSz+kIAYG067cHz4uoBJlXk8
rstfWrhA8WLxaU1A6B3ppKjDb97rJY/8f53sTXbkIEcywbHGTiMC9qj4mf0LyQehLaGTHXZMkKGD
AVcbu09A0ailI3CwDwf5QjxtTXpYl6Xio9JYLQaOFf42oR1KyCe+A9LP4y3CMGyLNj9I0nUzqVDT
UD87Q7h2Q+cdll6URNQ+ZU/wy0iBFP9185KTqjXeMq2Bwcwh44fCl77PEhxphSwjcekcSk19TQEA
j8Zn5llT7pvAWG6jvL+gNN3qb64sNNmuC7HNrtsHlxyB77NdYhFqIAj8/40wRyvXK+xu6QA0GOU0
oGqoWZQx3D7J2HaahKDeHQ1yOjwZo1wcireVYxylaGS7UWG2NM3y8DMPpZoAp5L0kl/lyLHMKK+l
8zcg8p9Ia01aawDzJB7HoPCSfJs5CKndO2/ggDU+Rxal4mG8MGFDtl+HcZ62SEAoHFl0aZUB8+No
6gonPwHMIoRBx9qO4akOKe0OpBI3ldWYO5kHn+i6YL8c3mGTmy8/yF5S031yqjWCliUgwxBDF8mp
uIFsvM2QGI5UaYnS7R0It+wmwa06/W1HC6cNe+lLmGFrMDn14ESm9QG+5Cq2oLgRJrF26rHLq7Z9
tFKHsI9HcVgeaV7n7AUjqoXEztFdDBjSJ2mGlV4R+/TKUrzmcmx8tgnMXOZW4L1scwW67xO9/j2R
UsCSZOsvHoQnz/taWY1B2WoLAVSwEOHMBSiVTAp4xQg+73Xek9jpPpiYWJRkiCYckeyAuC68NtdV
19Gzm5NgfugrxFgzGSmuyFF4m1hqSrH08FXXJwcqIRIgmtocBglxz5NWFYWPilVxfgvS6fko5xor
RzTvp+KuWWlFZZgMlWX86u6CmMezDv36nTpgxHRdOcskvmAELdpYGwLYfogByNzL6QKMk8qjLi5Q
/w1Z5e9YuUDbGqRQPOuFUmqRi3x3VburwR0P5O18CgNkPdmrjjufVRdYdckf1nhyku5vNTJiQQ0Q
/hOkKDDIqJmcdRaaur3hwXBA/VTt7AUE2M9B2AN8jqC6HyhCeGpQYMlKohl1bXFLQKNBrAOAErKD
EoWmdqF09gtRt8X1yddjWZhZ+yqHluZhogiIA2PwPz+pQvBAY6jj6/TTtVkG/LURiSJfbUOGRuLB
xCpFWp8SYm8MkBQYdBvNs5x/iqbi4vMpvWP1/aBHhNbViZhM0453a0k/bcDltN8EgOu0E4zfFF5j
URCkhO+J9+3bD04AkmzN1O9awo91nJiSu206bm2h631sGeum24cgt0xV13ZweewheeK9JtYrtXu6
QqLkWvpkQys1w5HevN1P5CI7ZtJ10JJqJSNBBq1leUJQqoRkYW7UUwcO0b75OMTCb+aoGAezdKqr
WKFGPUcaqYXnb83IM5Na24mtmqJbJhBCkS9wGmzHDiIwOnXv5lTv4U16tusb8wPmdbzOpC0rSU0a
sDDwFCUVdnG0FWnxiEZW6cskdXS/Qy3XGZ4Ylf6eUJTFatjzgZAGk3S8Xzbzz/uC70EMkdHtF0kD
l2zCVAgyNCmtDitN9jxfBDN3iJWyVB6QV6PTeOntcyEewQHx89dzhQbjdVocSmCaRWxJAn99hTIg
LMdHxoHra1bZ/KCQauk/zglsqL4efwXPkTW5cAHq8yXqb9ceybfbOwU3bsJy6TqFH10uODYP4DNm
H7CPtxFJiwVvZpqangCU39JGnUioIOCitdoQ12tQ6SGCARy4emZf/O7HRsWDNbidLBZYJM+kPX7z
Lqmvv0ibLEPfy1q8igjDLyDgALIdSwkwiXPFTtjubQ6MOTqWypBRCXBQOxjxF74JaRg1YQE8l2JP
siw4PvI1HOt8RCXSI/gtVzwmkRe40FvtUfql9ay7Sudqwui2EgTMWib/qc9XuVCj2FvzNpZD+NVB
IMxjB4RyIWgjUy6Ltin8l/iF84/w9qra+y5+jmfjbwz9gh4ryObGx1JmiLL/Wm0hYVmDuYMO9fbS
9FHoyf7l3yf77y1I7utoTuzgWskeed94o5339eFBDx2cPCRBwEuHminlbBcciIN14VowrknO3pzT
WSUzJJ8btlHoFWYuBmiB42B5He4OipX9KP6yLy7gpnxNfV4c3RjxVbjcyTttJDVRWE0Wuyly72sH
5zDXjYLn3wTeZC5vNuLdMevG45unj7+Fc6a3diKsQrr2pO+VXn/GGdTbNpCP3W9t+HQXXin2QhBk
btSumAcUlDQmBWRDEoC5KjysIe0kLFirmxvvWK/aUFNNbE79Yv/Bv0d+Ffq0BwRv1AHUzFmJlV36
EZM1P3KuBCWWgaHfjDS6kSp4Ybghzbe60CX0x+IpbbaxjC4nQAnanRPR68E0waFgu1cdtS3EaaAO
5GyD1Lijom+XsZbJXww6tNXOijgNbBDWtv+CKlCvUJsnr5T2XXPTmLbM0+hKB48uMx0yXLKl+3iH
/1eiT8+nfTLE0YfZZevgpiNAefXYcEkuWA9s8MBFmtIN4fv+xQpTw3b+QUxjlFH2TP0lS1Nn7+Ch
CFHmNu7NcjDUEcKDlVW9/6JrGtyghFixM8KRvzivhaIajOXVEEewO5bJl/dJ8OBut/ov+gNr3spj
vh8lo7w8SG7zwYobADa9RdQejIEsBG6zJVdksJsBjgnmcTzO6fXU6f4/uNYxbITJ+6qECjN5Aqxt
VPBYCcKPQFxJtbBB37PQ+LlJhL8A8WySLyNb5YpRakjvCINKVRSltc8bPXb1JxqJ0f2JoyiD+JL1
AsWF4cmwCv580iDEORy8rClRbKg+z4ccC9KcXf6HKgcP/HEBq4vu0Uw8ZIOedCDnfKw/slR+5snj
cO3JVNx/25tqU1+jQ343a5Mdz7JL36Irf9b7VvZRD5IBZ/k8Q1pHPs3+5lMAobGFHSFq4fqeqk8R
z5eb4uwAeEvrSyefYZGTQ8kbyAPhs36FuW5WTWaLYRew4+15ELyccAkITinciAncSoch69TLFVSI
LIEeQ7heJ7uRXSFtBGhzftSo1GEz0q7Z1hmQP+0whUticLySARp4xjh05eXqZlrGN/sYtcr5oc/f
EjaP16Uf2g8xAoyo8TI0HXGE+7/oqu/l0gh8xj58eXnV0PeOcv0GAPiXqHkU0Iq1YNjkyQ2YErs2
Oj2ceOXYgaWUPe5EToYzLISeliGwFQAqwVNvFamhw8uxsTi5F1ZmY2W4VdzlA9L7u5gjf+5Gs0Qk
kLzM5GgQazW/yQfvOoVj2PEM4eQSxCpvisCKY8apJY2Aix1eNKlw0Wb8ba6SKFBhjIQPNIj6mH1R
lBm8cmMPUjL4QaDV8h90eELQBRvYW3oC8S36XhLki2E5a7ILBc5Cd4+njSjobu/S4dh4B6wDliAV
QHFDh+ARBg1YT+DfHfVolwnt8Oivg7ATDB44Ebz46eCKuIxMRcOstnE0UB5OcEaBFDiSeja8PBKz
tBprmVsPOFKTq10JhfzwnKpVfJetlxYU1Gdcaf+tLXmNGTI0iRJyyTtuZvq3vzO+IZthpJqbjI18
MKPNFaUWzwEgNi4a0nthGjmd7/P71LEpdtWkLoCjTVjA56dhDiikZ918feV5bZvHsCENbD8xx+NG
3YrnxIqFMvhJ7f3V3mlC55MmoJU2soWDwKZ22NMIK4NG34Xpax5ruaX+JKaD0Amzp2k4jmS5Ruii
jaFMdueLTkAJGcZ5W70T7NLuBj6wcefOFGqY9gF6iNIac4xFHoDFMSe0a35GEAmcnEh90TVKOt5X
6ziSvehnz4AkRx82nuOBHCGpd3C3RBVdtNjEyHVPv7j0eSUgTt6ac0taz1Pdxzk5S/LFLpyQdtzy
ijdFWt9P6m6gIG0R2cjtfaYzTVxCe6/iBF/NkUX1nByUUGND3H53CaSTBgnEn+UWVX4qqdBh9J6b
Oq/8KnvLRwc49e9Ps/gn38tCV98pWXCxZBr81gotcwXKSl6/X41hM+8O/x3faICJlqBEQO3l9gmf
5oAPSfhmUD9IIL0om6ZOjuvDR8ED7DbSpnVFmmLHBeT/+IXnVgkVkPUFpus2ikWxGdoRRw9A7k66
r7dN+GCOzoniqYWciAW91FaG+okwVwtK9reDEsiHplY/n2mj5R+yLTIbsjlduumqd37nAvRYCHKf
LP4nYyAGGXaYjiQBwLRrvMNCoC6RhNLGrfhOemGJQn9lrz6+A0pnTdnotTYUdkgGHJZXtQ2IkULR
z8BGnnzkTUgFeh9F+HcLL+W9yoj/WCgrzyLYvNkT3O7gynbyZ1x2fCmSnDMp4C7XLwr+FSwgs+6H
Pga6TOYUnK4F4sFZs0m8v5kKFzV8nyigxzzrKxaONVoPPZJ2chsj3qyPL4AAUGVKsgloaTyz8yW8
nsFxBdqZUJbydjemyhBUVtt8xm/uutg4ors7cqzgbGPjG0stDmD9RGCyJlbj9A0xkCJuUQbIoX4D
HRHEW3PvlnaXazseMrv3FX9FJT4i+r6D1BZtlDu3DXvJE1zzOLGjfsuZqM8kksod+Hqe5EaQTfB1
c4jvHApDglfcXw6IWqPChp2v7CDO6H615A/0w/bzQN8GEuErxMU2zs7Pik1COjon5xpS9ZeDZNei
K3SBP4YK2g/sCKbj4zPoIgYNLtvtYfdmlFdy2rE0CZWdoQ5VDMZNa/TjVNZoqs2F0auukV3dMOaT
ZPlhtyytzFQP+IUIlTKMb0rAltzeFrh5dkYV+e5034WPJSUJ6VnmhTKo2lsewOyajH4hxP0MsjlM
3x6gxf2U9HcBx3jtJ4BksJ4UPW12X/ZFcrMTvp7cn5zRW5Bcj4thOXIoD/WPlVNfzKt7CiNQryER
Gf9Sm46CFjxgzTioRRtCoZNW7/cQrjCR0gSGF7s/XV/ayJ38zeEuXLG8dgaXvTzkZEIWmobzD3um
ASg6uEiPsGNE8gBcQBHOCgnUyuFEmjQwC2iup8Cxn5AjpXncmGscjLBiBavh2Ah81NJEaIwv5lr7
s9aykMjYOFqJqXIJhnJPF9hW/GanVYTU0pfsVrPamBKqBiTfWJXUoAQriE9tUeOUcgCiDPuShp6E
T8/sr3sjnBZSA1eeHyHqiVrnvg/PjZME+m0ENlmHrLfdSy6X+bk/16ZlRAmEXYCesqiUT9d3YCw8
sFZogrVw1lWakT+n9KUXpBnlrgRzfuz/3kleANVz1+ZLYEeA6gmlef64egQtLKArHt0hLW1UWhi5
9hM3hmuts7Msdemsgk9b/SuCbUmGgcuwycgh3Rt4z+DLt65hnKTfCgE6SwDFwnTfF3laTonXP340
O3dtc7Vnhv7CiYNSlxEwzKVZG6a83HoRAY/Leo2dBTy1XMyuX1696zrE6cEBtM8AVsEtoQZ7GvEj
eVnEeuhN+Ddc4WYtLOmYyIGPxj/sIHeVg+0L9jYlOZBB97uZzhVVjFh0WJxsY0N0Ig9EVvPv2pvc
jSfXF8gFeFw/RSmUOd5cBnfr2kRgDWJaJ0vPH+vu3azKozprYbUfeyBILK5QIKcbq9u2XIYAdE6M
37Vg2y6gxEJQfMm4k0Jix+7FpugDB3D6E7TyVslD7VZhxB7MlQ8dkx2peGXumE/mFfuZlz3fet3t
FTBai60oeTTugqBdkoZANT2tFwmgXgwmOk35UbqRxMmyBA5n0Eb03S34vqlhnIrud3EoRHCDZQQI
tfj2s5mNiL5p+WH8ZF9gCDdeBGzO9NamVoc7z9dBfLFclxS2hpZbpeYujBDs/DXBtfbIXWbvlbU/
TR+8XvUOLnbfMe6fXk32VTHawGw/1szq9lOOZXfNr7Qd+/3I4hwouxiw6hqz8bFbipJGpGbFxCO+
wqGUd6MNyH83RNlDPS2bTpmFWm8NCrT/7fs2NW07xxdyr3dfTq7qMjN2dj5Y3pX8i9dkfQyAyJZN
CS56X/xTR6etam0ENynT58r3BJoShkMhOWtmlyng+k3dJiZpXLZorH/5IDNo6IrfywyMLJrzYQiF
IrSq4dgavIlQR4iu2dnDVAyBHl8JrOht+86Q+A543fZEVdc2WYiXfxSFSoIda373Yf9v2MZls6EU
LziaxGajL9cu1DYnkM3s3Bn54JiklyoeWzKoP5xMscT++cJMFeNibqY0/ECmaKzvDy4cVwd7lgkM
3MEsjyahv/a4GrO0f2ftWzwuvRm2R9XbJ3+MTWdICIR14C4aOwLTcUt6x17NVaNs/zzByyFuq2bz
9wOP40F8IYQYPrDKImil6pyLGUqIub2adjscn/F7aiarJA2wqrQlsybNiGBDdRsd8ZHHWSGa5TC5
4piisjUVeVyfb3L5jbfAhesxL6iykM+LnDOh2XbiSewcw/+f+IQbvZWQXp45aTjWWkwLKPArNd0x
eUG9oJ2sFMRUrOYd6jX9N9Bv67TOXBTAL+kkOOqdWD4FRgw3s0xaEGIBAAsW5jCHBkUABEYNefpN
GduNc90l4gBKDnXwlGBMGUfPYRlucSCr0p0Xkyt9NA1Bo1tHjR1ecqL7r/jyMtXGfWoBV335nHKj
Arycqlc7H0Lf03mxBY1hYDfTE1Jn0HH/XRWSx1DnIuwJMuNcp1s8qy+QJJX24wwkwEsrnE90Qe2E
zKVLbflmjPmKGrVaNL71gmAh/emTrlPdN6Ym7UFgXh53IBITE5LJM83Y2hz4cFUqkuvTU6mhSplH
aCoNzG5vQtob+iqlpTheC5Rk0HuRkccqRGK718xxSQwngHEtiTaZD8M6Yjo6e0N9CHSOBVCfu2Z0
pwfZamagAoRTz29Rw9XSIDUQMqQ8SaAAhh1ZdHp2cHCsHjzIcaS3n82YzK7plXeyDjEsL/djYZ/2
9i3S1TRNmY7J9VCs/CyrvsMTbbsgcYj29Q5/yx/w0dXy1uD3JUZznWKvRdRugrXzjGPnd4bvpYna
pf0X2OnJ/fLTp1JwEqVHehkxTBp663tdvwn7One5aCS06syTufgM1ytPamdWnFQCr7F4+3cX6nEW
x8c3LqbcRoyHTXup6x2wIfEXVy+m2oSAi6xPM4nr0d5bB80ydJOz1MIRcF+f4WEqNlea7hqpzEwH
3l+1Db5PDCk+nWLTJgbYb29SbYhRF5l8YmRrxnCwUYIY8sQCf5ObiG+SaWDSeQxHab/npFHRGdz9
wZ4/4B8Rn+zCrMdEyc0jt/XN/1tOGaVK+Vcl6GLa5V4MGXhkBIdnDu2+/jrhffm/mdK8UMbJzuSY
zoTHPGyjvlYFlnAk6m0LSWB/gukMtL/ahyXdO+5jmnXuF3Wb9eNhL13w1BjcfPq/DF/bqOk1BQmK
yyzbnbyGmTO6SemvPFqoF0wa91QHrlmKKNcXsJFDdNImKYV/hpges10YYcO9WxPGLZQ0FzhI+pyp
MRmqGIc9OzxlMlsWEv22qpTXSly9nMQZQTozUnD0bOa3OARPso2pos/2wMKZ3J22sHkJDveFVHJz
xbK66rJgHOqusqdjz3/6I9D130qOZtZI8q8gmfMMztWc+ncQoA227fdWCvUF+gSBJ3Plaq7QcHsR
mO05jDDRVNUZ8wf3mM5mlFNUxcbghpXQqVDv2scBAw+Fa5e1diNkBcxiZIlhGzf+Iwn7SYuvwTfQ
jCyfLV/Njnxms+tbVY0MLN6E8UlnTjo7R3DVaK9ngIG6vy7vbk9eMYLOOXNtJJAbdbaKm35aLMzQ
rP9c1KIDFQ8rIqXD4e+I2oBmEMjo9fs/01YVTqF7TZAUSp8wFKKRJeifVi2mnMHMrlTEKeBD5oYU
7xPkrYI55YCKzymbrih2hu8+Dvkf0BHOSubLWOUNNA8VOuYDxafuYtYr8PIKdc6tLA5A0AZUJO64
tx1+YM4xqhqBH/Ge9SSmqkc/cUO+WDSiYi6XqK4HfK25SLTh73v0ePYm6TO4Si1ni+0ZQwTkuahb
e0KeYgXWNKYY3xvp8GLFxCOYcspWOKH88B9P5W3P62Iv7DVv1shrgEMh2Fku38oQPhx7oruS7Qdz
ARdzT48F0cnTpLGl+cZhJq2m3Q02/3q7k/TKpJ2/6rHUxOxEqbkJaiQ4V4qcC1DLm5USGSugVisC
sCoLWkia/VcG5eqS/GQmEeiON1hulK2XPRx+qZ+qYDTgYXRpSjVMVD158OtMHnyhJB1df0jH4NXC
I3J8vFBfpgWjeaka4lQrtagv6A8Atyc1rXg4Pn0zrO2Esg1nkK9uWKlhqBUh/RmdpBVlRtLnBqyt
6vDJEfroyMzQp/TOoXoUcQjr7EYCK6nLnHliOJZZuDcYQ4eijO24p7AULQELplIhVe329HIOOFMZ
MHuDKOS2So5TZPHng1IZ5GHshyR/BRHEFhNvKvjbIHXaraxVcuJ0eoSu1CuqVq4ngAY9+LyjG3hA
OLWKNVX/XZMtjVB7nwRV2SqbW2k7ULbhYZCZsYD45nyBVLfPx2qe1vnHTx9m5CLKOVUUBKzF7Wls
hO4Kc8QNTF7jE41pHt42nJTTF8DOMtZDQVFA7tclNNPVIusNHSnCaGyL5cs9JE7qioBdyX5J9ZN2
5aFBuBRRpg0mEjSIQZHQKvCZD0FI4FUXK6kSMFJoSONr/WZPmSQmwtH2nZPuCdltLozFc6F+Bcs5
9TMtTvGpGUQsKYsOVlPajeU+h4RE6afUb4wwTpc9b9Ec0VwRlYppo1PNE1PHvyMNM4a4GiXuuCQi
ndSElP01Odap46aT6kZG5JOziS9PUV4jC4x0d2sD4n06//izAkvEKn3dt6QJO5dbHlAbRX0EgMD7
i9XhcvQMhdEFa0KGTWbdsdwebFLXloD4hJtCgkTqsNBk6q2k+6HbDrWBjd582mZd+SwGFaRpKP45
36Z90T0L9rDxpVln/U+8f2dYyepXCLjDOF/e+/7Vl4LWFDWawJ4wNvaNy30WLGNKlpTjmRywqZaT
52PvqLdtXunhoUJEFKBCLojrzcYqQoWAHql8JMuyzQ880/9JxTJt8V/byDqWlpBA1U4rr/cRuoGQ
U15ZeTY3/ZFYtkxAWRhPFCsWLJ/EgMQ8m1Pa2kh/t1EL1/xblArJ8pnFi/B8eICNVgjUqZHyDO5X
76lK6kIhz/p9o+Rdc+0XWctsUlzVNakqP2mTZfW52F5FuYxFKZbc6L4logS4gdNRMERTxSN9UmJ5
a16GdLb7vxLgUa7hXp+mn62Mm6VwzcM49+ls/Qt89OWtedalUMyYz7MnxVU1bccGUxRVPHEzjOh0
jXFCeSOOqO75UPYhjk+fvyv+Vx59a+C3V4euAs3ZB1kmeSqEEubZPPeD3mr7XneMIoZ1cZK3KlIQ
MK1NIxUXH2F7yDEvk/qo7PV4gIY9FeDMs+5wDh2g47A6K4K8WgWD1ndqnuTjlpy0MSvbmprLmV+M
ZPRVOqzHZh446YdIQD7+nKZ5Txhi7cRVu7e2AfPo7TzQeD21HEhpz3Np0DC7Fzks1AP2ppUBHFzC
PBvK6LiSpMximUyzQS+6593DeTlREDCgE8M5ku+WWzYlSLvn8ThJVUytK3A8Rnm2ESjcLQqywbI+
SVqBLwMw9E7qwcocy3pqWxVNBHFAIVH+0RMhnR3HFM7WxGCt2vsHzQFWGUk30bK7Tun/do/r5M1q
YLIVcYs+YEyCrcC9Pr0voG+6peA69xadwY6brMgy6c5PVuND7EdgoOuwp+h1pvGrlx7qPwJKd0gR
hee8E6T97IrZFHGJ2neFc298BMklIKlDxntDTQdbqQcKzZsXZf77WlvHj96E92WBvmvuBS5XCtDs
FAVLVGkKXvFfnKjG1jn21mx1JXXRYmrVUKFw4hb9qWWzck8RuNIoY71qMamO0WWf8D+AqRnA6QQp
mN2I3os/Oxbg86dRD0OK4yiFUz9zXs359lgUi72EQNQ+92K0yVLcts5zkfvwfI88O+9RPR6awN+x
dk/2IUjao9riLxiczn1wS6kbOzkcZXhrCm7ytvqkznSCWvzoEa02U52vhVJVo8IeuwtvrrzEkACe
kU53Zi02s2MUxj45vFcCgaXzULojem5NEuGo/p8kqTe5czAnxsSAbAQRHEabkRlnOB4gqWPG5Nc7
W0k+oVBZb9rQZDYkYR8SmRVbWyBAQ0tQAVmbnF0oMpjsnDFuD4SWA6cc+VKxgi9C89mUpdGG/Dq2
/DyUe2m6oNXRlz6LFLgr8gt1fA8+f0YgyjMKu6EwXZcAHfYe4eAINhbjEQfm3B5QSTfYSOCpmTBy
hT1AwgmMpM4Xu23V4z3U0cBVPhN6cMpCFlQ5gKLwU1FaKjVqwPNHM3OhaouaqBP7MHpO1JNBDBO4
CWGudlCKXqFNE7hitj3+cGHJyLCz6No8RDjRUpxnaMYCWjTHL2LALm73OmRVcrrTGsNwdJsKByGi
qBeGID1SeMG0XZ7I3hUX/rH8NvVjOo5A2yjbR6F1zfkNCNRg2xFfaRqL8Xjw/8iT4AqZySUcB2Md
5Kr5xueFRdNu3OkATHdhZfgPh4wsNGB+4c8UIT3yRrYOp2m+XRXDVLyTXEMzhQFkDYsRYNFUr5Tk
LLB9h6W6+DoOYPwCBCI5SUZwwf5kP9nBNvpEa0YuGK5xXh0wRXhve4RUmrgAqWg3V3BbyNQ1YhFl
ATdoZk/J5DclBENMcpqK+x4vYUAXwA2WAJHkIuvwRmctc6uQi1NxSfhcyryI0lmyGrK//Jz/vXpl
mb3F24edZHL0H2Xd24gNm9k/oRqy7wwCzQfXos9LwMDT/MFBR6Vq+YuTeq/1USRcgfhefQJQ5L3H
raoFMIyvkZ1QECImE2uMjdiT2Gv7RzFaIaLae1JOkev22lav9+Qol+cPypVEHDBItqhzT4C7KZrs
RzbAjJWsXtUsLQE7DGJ//8SZ8hbKRN1u525068c8Rn3opjAuFma8yrxAAddPj3tReHSNW/GO6yeh
oZpfdl5Hh/FomqamiX/WNoZVQ1rdg14B6U5GXCffqSYpYq29hZJk3GCiBZqdmwLPDaVZzR+YFZzA
bY/scozmR2rW2S/dLrdp2w3s58Us1vpMsODFWtmZ8lQ0MOjmTZINYyXVSmEv99h5Oy4XQkFVzlAJ
INvnjsbYFtCYQmdQtq0IWNIF3aMEmWAa9DFwxk1bUza+pGpECkidEHv5ftjBmLTPFnY1IozASZiY
lpcl1sJc83d7x6jeZYdIr/OtM9i9pZ54d6dnzcuOBrm41dVW+/VZDFlQqRG4WKrFGizYwrc7RltZ
vtazdSx66DUR6N+5UxnwhLyVKFpJ7bEUaVOYzd1BZ3/dMb1vnLWWHw4CXavhpv2fyTrq08q4E8Nt
/GkfYu5X/3SRIaxYUlWxEK1qKEDl9vFO4dTsHsOjkHWgMXYXTXhrvGgL83Atdznyf2cNiNWdhmyT
Bk2gAknK7/oy0sF2QtIryaGeGPDa1hbHKAKUXVI5rYVdJ331pDkRcnmaE2iWvrqm+GYTqGgbgC4t
Z2Z9wb2FYZsofMPm680218v4qND44tA0GvEQvmvi6XsLEKIlhu7uNxojk52+ILiDLUQoQwmK+TFZ
l5XOk7fvYASfBKCm6cMZjjxbiTFr/sA4qlhAQ2MqBSbFcYpVNEtZCmA7kzq6DLGjeXQvlrtDteqS
tK+9e2Nmn+AoYUD0ANL5MwYWNLwVFLd4OrUGK3hNBmhQk0krv76YRPk7gwE72PSupaZhoyB91QYj
ecRmXFyCrid/2z5uJySSoK2nrzl9GFbCsQAiBopDz3t2pTD8z3Idv1pDzJ4YH5IZZvb99i7jVSKv
N8uu5OXLN94GHKHhJaoRz/bw3nKnsqTF/Zexy70nbvwoMMr9J/Y17580SiGaePSAMUujjEz5Mpmg
PvgTnGf4iRH/QHq9YNzlYMNwnUBQJrn1ukNJ8kiXVA32dYipzvUCf9mcTsN5ZcK/N4r2dPN6VUUi
j+OvVP50aD4Vz4uAwUQ/8IB7HzsODscV33ncFS71xP/KhfLS8u+DeHkMoXCTIKfXrbgmAzLktPDH
ghZRXS/uQP+wBbCrzQ1XUlnGs81IQSJb707hQ0ueZV8EmTGWcHy9MKIX3p/YUUnp/Zs6xfs0snRP
dei/xAu2BMttDInZDSRizHG2nkz3ogHGtucL+QKTOeXOfVHYf8xra7yNzVwl42/hEbjPawihvlOV
+75uoMrgV23X02lcbq0mh3G70gdHKZISGgiuWNTU9feRvYk2z5i3DrOkvHkdgMl0sq5SsmWo2thR
LERpY66eRy4AwJQXTKu4LBfm2fp1HEki/oTOr4B2dpC/FdeUcEVTRdx9I8QR1RA2Ve3pPnzN070J
h0uqqGk7ia9JzJtop/CpAI2gFQs8/1HV6ZFviN24Vv7pGVIqEsPWHw7TXxblnKnHZDvA2ZOjxDos
gAVIXIJxEQnJKVIPZjno/in7H6pIk1CGWEasxu4weBJw5iiKRPVupUH/vw3eRwI0vVe6YF2REhAc
/Oayh1ifiteaeryoulCFmYckCS9dbiSmnXP+ec6nY3HGB/BxcXeGxI//+j/yJe1LLRMn7uLPd8nr
daXf18HuShXSQTXiTYWgRbJ106EH2DOclD007Z4hLxS6BKEkFVMSrZ8OXHuKjmyQUwNfIPYXuPzF
93+DEr4wzcvR34z8Xw5V3plJqLNlZI4cTv/kVKbmO/SlXRoYs7J3x0ObJ2WXdsSaSfbnkTv1unWP
QJbDF9S1EfjbL+SEMkRUX8hpUbxKYy99otVUceI3ZBzSIEFcK4sNKLLWw/cTtVsENhYBTytLHmWr
sYRnsaMyFWXawly8/AT6F9imr7Bc6gOQyLN1V2v+G/utXijQpvb99pHmQaNHA80WwNqrvgP0wGpW
XtIJsbP0/jY+lqaCmCUXjVqGNBgfC8NfTJ7LHVQOsTxk9z4p3pA0EO7j2uYkbSm1OzloqoK0LNr6
7eajZyy9/34YPcSVbF8r23y++txzQXBdH1veSHFjt4VxI5MW6z8S069AyUwIMBOTB+lMW88wPVHK
iLKiqmUZUezSxPcSKI4c6SMIivLfaPa2kX5IezVTUMtDDTgNwOpBWRH8KjDvDPJRec7/H09IhpTv
ZF3MUmQ32g/Z61mpoxfZk1YFSJOwi7RIfNP0a1NtCqiAYJQD5df+pEhgF2MgS01X48B4nbiYfQ0s
xMsNy2AFjV0Qt752xiIsrLCk78BQvNw+r9fJuBrLDQyLgw9KN7P1OiJWWAYQ4MVL5q5hRyHhZfUI
K2aX/Zl6dMXhFNM4K0+7AMBb92dMkoWFBMnd3mUhvT2Kmki9KnJlsnw14VAkS6fqY0IQFcimcxi9
qqkQ8d4qD+VRSIA34r+22UezxpfI49EHPclMa+YRq630GRgzwdjeXiYIkyuEmImrFDnw8ccBCsx+
ML+V6OHQAiA/P0vW6E7ADg48QcqiaILVcLZWzr857yjzGhiY5CNW1EXUnBmOzHKPbG3l1OiSOxTS
aWOu3A8mgT7FzwsppASFgR1K4zCX5rEW2Ujdgh+gsnBD4sdFroiwGv2j/KrS/Dkt7+SnhIq5jOcG
JncHfRwsW/BfGJPOOeLQJvdPCiuukk2euJeghpxAEk3V2/E43TzatbxSGcRHxRKCJEkQiXKqW71C
FNhABl61FqLQgfbwQwwnSAK4Ge6Lfd2hx50FCNB5fZDMpiLwhss9D4NvX1061is3pSDGxfRPKTvg
bWdXMy0fSXD+s1ACHgc5+CNjEq8PsBcO4wl6W2v4zaGa15O6s0IUYhYuWV409/qFE1R8mYfdBUEy
JBIScsvwZU8giIOLY8si56cyoaIgF7J/voCJt66Ym+Ky4gJZ3Tx3a8Sw0wblfZD4FFvO7FGIaWX2
rZFojQfOYTMwIcI2ZYBONwxUVunI6P+2pT3bvl7cCZOEyqbrwyVGy1NbhFm3lWv8A2OYkyumXW4s
J+0pLt9PF06qLibgLeNO6kP8Ci1lazIBpx49N+7fW51tSHBYbfVLYJ82lJiCjaHQV9ClyO0vI+dN
Al6jcedRKp+2DdVKJYDJErtXeliJy1pU3+oiUOYoojOWPositXzvIBKeiIgYuYqpSm2sVPFWuBhE
fokBalyfZcgdN9yheryYafSke5mE4kG9ryQhhU9d4N6E+rEb6qK7K+wILUJ5bMD2CdG56DXUFjvT
0mRULSzUr5zVCM5Pm+dbn1mPX+V09pACLJ/wPOEAss39WqI6nZsas5dWhhQTxl8OvwIpua80rWVx
Q42M64j85ikaitCrzbd4VEtFFAr/YOUJByFYVsHcZl6zzZhf2+UVQZNRGjECHeDDsDULcn/DD9QZ
pjA7kuSWCakZMSFqi+5RQdmluSAdSgKAdsOMiOw9woDbdT4n5VtSbfaClxO+Ik5hsXj4GkkmrS4a
6MtwKfKLufWT49a42XR1baqSsB4oaqKG+ZP9sT7PZSnHYNU3XuOLR6RCyg3UGaYMbjA0B+sPPTps
s90lT4aafNs3gxWqKyqfVqE/gKjSBcSEEY+eZa4I5Zu1BPw33kDN47j0Mh43ewNz4RF1ZjqkQn5Z
uBdZa2s1AqgRFuahT+2CQ2DF9fEhRNRsGh+FAeDCM/Xmve7bJc9KA01pY5XG4G+cNM4WzNufks21
vV4bOnJkkiMe0PUGFIIO3ulAjHvMHXzRa3x+0At1j6kAZdajNejxhFcYLdqEIG+d2NSoMOmRJLid
ehbyQMU8svQNh5TrynRzcQX6SH0waV9Mxj3M9DO6mFar28p1XZcWDtL+AxAYBCiaw+ozuazf7Dmu
hVwXwxU4VmV3vg0u4MUh2wNrnJGPSgdRLhfc1WvrDvlp4y0cGnYMLriWvykyJH8+Vjv6EvOvi+gg
1djKEmNMlyejYRZzB/p4cPl/labDVT0O/+9Yz3LwTjXvw7eZfKfPCIXWoCM3a9aIRI6xwaXri2cK
LtY0Xp5ZFqLfRPA28gqkNJ5PbE0AR9O5Hd5eGxE2Y+tgo3XCb0C0Xzz7xnBDMqh1/qC8ZCh4hoJV
txskhFGQ14z+ITP+yqFxOnJsiIxVFxBgvN35DLNdkFDsDSJd2BK8bho0/riVlkZTP7P4eFYdUWsx
SF8TBGPYIiiB61wkt2lsrokoe5d9Q8mIs/QnDFBOpMM3RZS9p1KWE5/Uer3lofrFlzXZ9dLfysF5
J2j+T4IAhEtsL7kAa67NuIT+egnlVryHGVjEKtShwrN+gHrdpqWYNpI4XWFeqPuR/Ax2HYVcFe2w
Khc9ipcm1DUMCimrU0SCu2uciTiS+VYv+i6FnMJXL375UzkguhbBwUhnCDOh3kEuRufgAgTbkPts
ZRneTESoAMI8apuMYKiv3rzj6SWIuqap3uJOaQhuW5a9UZQpt9G0rF6iAEpqtrLDNBt165RAgznf
bKCeAng/313r4Uj20euLl6R9/HvigH8XZQKWuf0Mzm6YToS/VO9RfbPoElGoJhtv+RdVtqOI9FX0
zsgd5htrJBzuQeWqnLvxyolljer6HXJYKYRKgundJmt2VCLJu9n91+rmP2md1drMFHAZGMCSYMJ7
03Cz+v6UslNjBINs9zd4wFhUX+XNeFTgCamlRrBbWMGzYmx/6xjnS5C59fy7bwWDtfh485udtmCh
o4LC8qSSaz7FSzGQPKF5ge/9RrgMEm543UflXrc6HYr31bvDx4ItMOCW2RjOXwWuyIG8spwmZfV+
mR/B29VwgRXF6e7mfEG81KHUsKHnfAD4ufi+NjkAWRERkKfBmaKdcp8YWl5NV0AvMI3iruRIWGM3
4NNrWSlUWzKHzB5cB/5hPkjMec1MPvG4bjdQSK70GLl9JPGV10QaJ695LqqP1SO0xSFC/4WpNYGY
gL3MrtVT6rNg6LbcNANElBIgKIWy/icMXhqndMvJ2zyJ6+ZVPyQXh+KLJU59iSE4CiuRfmrqa2YT
FqSUgK3R6npmDcnxlfjERgtlYNFuYoIwhyrMxBJL5QFksMIyadGjzCy4NRhbply1Q9BNYxG14AKY
7sbehMXvbvF1NHJpMec/d3QqThwHjIB2ElIo8S3QTg1zlXaQBtyL3luy/omzZf6mblzh5zMfpHUp
+MUxC5SmO/B1O3Csaqn0wVc8zG4fbGkChP+Up4KcPeJMt+6F6VhELdHZI7MHJS9wcVHeIZqAXTTJ
tLS9XqL1v1VvdpH1qJRfUE8J3vWGqOn+W4TEBA2VLP1E54vkkcFd4bzZQY/SdnavI2PxJmiPMj3B
WR0mhyEHi1J3E7kpUKBD07KuuH3aibWZVuIef6bKbFbdp4ya9x9vff/qY+Ks8Af3KJGnT61khamc
teKzTiXks0g427eX92d93rOSNTODpw2qv5iGbO5fJWvQw/wIvNhCuWQo5OdhNJbdMh8pNNJbFu5P
CHhdrhy9YCIriBuiqBUfMWmjkstrYnOasC44V+XA7FbzbOtm2BWP/wphQIHYQKmZCH4O1TGaDsel
AwGmTlUDN+0GHuEh3i09L7DHjgKIxqLlpQAFBgLuDIZC1pkRw6LK2YF0LMDbWKHifiNr1oHq6RVx
FOz95TDaC58HEh1xO9phCzag0bVh9h2HTax86eqAQ5rP+Yp0J6LK8tvHW5dw3vwDSqriIgJq0h02
XltR3akEj/9v9V+nQDWYIdy466+W2nnAIVa3JMB92RUUt5NbigtC/HQuRivLjgNf/0qoYnlrVIAd
zOxXvtvXxawXNnva0Snc/kAY6/GKGXwdx/EHdxn2fcP7/ZGFtysN3qbN1Y6uVDIRkQbU5C4AhcCc
LP/zXYYfQ4Idpl7u1EOTe9z5Z+JeJzlz4iAGs1bAvH+5ngxJ9IqaH/GX3VyoKKN7yaT3Qqm96BYJ
ykRDnYiQQv97nc/reCtVxkwHhKH5gacVnt1gJlVZwMxP7SJ7ZA0nrHu2paDkTDEPUjq4pR/eqfXK
GJrsD9zsNmk6JEG6VIczh08Ao7C2vXMxCZiJzVT2nxuNSTZbHGV8VzdxcJ34uzIASPAALLfp/m4H
WSuqsHYUvD+uQ2+jGSTXV9EqYD0gM9Q3qQn5RSB2tMOxs/HcunXs64CyUgBzV2Yp1PlXa/sriTae
a7nJ7ZYOCcRSQrgYGUz/xetvt8WWu3yP9yCpFJ8RR4cm4XqQylcGLvTxdMfztddxVlvZnQ3Hh2eP
L7HTV1sW0VZHfxJWi2lmks2ji23ycQ0yCZGde/QDT2SiAuOOesDhAFYiBckYU6WcR6BQdfuhyOrK
+eDjZ7hKn9QWA5TTHNkXHxA7mOhq0R8fVagmR2L+6SYT6lp9mzJb+m0Pd7w0G++8SFPcZmxpjibD
i80SWmsWOiQkts0jEEMr5U3r71R+UF3bbYfpeRJ8W4zfZMzv+FoGiaKjr8C6FqOsDj/uFbJsZXCa
re8NdcBCqUKuKWgqbwZlve4wcwbIe0yndReVrMvxYsjpMQAjvbxyni2CZFQHEEpN5Qn4ZfHcA8TY
iuSOIu4aGrjpHYP96TYrNrK7pRma+L9JpvEDIWtTxh4k4pWN9kGjccnu4Sbu3MfguHvW+b+S50Sc
IOFqPmIk4Cma6hkPur3I16miidhgnqNWb3J9p6suWHixOUFeCrSDsZKArxSTsjnv5jmytwuD8aPW
PqA0yojU5/F4XnASA2lvS3bnnRRxVZ9xrM8UyayRzSh8ej7OSolK5XnNxDu/WSeBU+Y/jTx5wBGO
9l6OAa1kpNd23IaY9ufitKmW+c+2hPc0qAtymmOBBWG+ahYSHXHzca4P++HZidgvQSVVWsJJJFwr
AE30XWKxH1/R9veg/kMl9LB5twDomprgPu5lv1SQq6z2xDmQK/BRKIdeWeVfIWN4/gxfBi04fNh8
/LkdRMDXmv8E4e6JdAz/VHDMw9P+NWHCJ9bQuBUEzCtcvzLcBmLpSX9deH6nhV49dgX0LFyePSMO
9bO9hhGbqdpbrXrAunLR9LCUvzz3xWM2GXSbR1/aKSV1/nyiNB9yFEilXfyyBkBu1yS8gIws4eDU
OnBb6VH2/+MwhTwIcM2nuJRH8UrIpnxq80kJptJWXckIFLU1bL7h3jRUqCec05MQoLe8WuA0MbHu
q815qiaNk3VkoV4p+SUkYw69Tyumx5b5/LnocjaOksLMh8LOw8yUq3h0jSHJ4u2KifBX2IF0dzPO
VLaf+Vy/WbYsCsuhXZp+nFNAy+29v7eGFJqD6K/bo10wFtZcTNH9BQpTAzs6EMyP1rDYRhstn2qw
q6XmUVm6umRJH6Bx5XSa/jLcxmKfcQkHtgQ+fiYB0OOZDTcKJs8XifZIhsBq5JwHWoqsL5/02MMy
aFvAlAH/1C/12GYcokO3EcLjNy7DSW1+gc7ms0DFnhb6G7oZusv9lsvjfwukCsonO8hX42w+mq8T
xdVgH7WgP2EkkT+vJGRQkt3nH22kTPgQJo7uaIkvgFntca0ov+anodR4WuTsRCoYn7f+j+OPAhA0
Lu9y2iBZv0Wq5ulvwpeenksydD4N1ZS0MfrHRONoWakiiVPM2RgvZRx3MNv98deMpa/Zxu2buINV
h3ihzWA1AgkDwhJHoUiym/m5Zpn6sL6h5fB4Gzyy6Hw7Ud89mSHlMufLIHhvgHTe5VjDOh4bLrID
FRTGFGCa6iv659LL5mGdLJx1H/T/MH9o5s/S2lxjv6Nma6clwDVBW71ewSxm00yYGyD498B4vqqj
c69CBhGAexqXpkZGvV+UarDYMflvgYUXuqKT3Ir4buO3xGbfAGaMuwbDk7qQpKrCoC3KIYSrxu1e
XZRX9vjYWfSPSdzk5zAIA6vAOX58L0fnRO977dOd6f12sEKt0HCCRsSqf9HhDC72V5hcTCypAF3b
31TdfgdAJmGJBv69xI87doWqZAHc2jMqgUgYZGbdPgN+Dn4MG8r0Yz+xsy/M9zr0AR5MI+yR0pyp
suazn6BGHJ1/wAI5mZHvkBIaQXURbhytzSCkigFxHVstasMG6g8oHFQxgueKZPFNKmhYh1nN2929
mQBiWTZbmBv6XhsFbk/uBGMzg6u6mAt7Iqqt/NRiGlUGN1ABzUpYP9jGf1PtqWqxfpukGIDURpvN
/ENxWKtT6MO86Drci1qXOh67HaR815o5HuL2mJkRVMwAS0MP74z3UCvGWpCQFliCJArxmXeTtrMU
ZfcmX+cvuK1tFFbeLjhOS4YWYHFIYDFRlWYk88b9/oXCjxgcP68HQZvVAYjw8dF+M5bTkDcG4gGH
7biSfUj351SYPgwKnlbFC/YMYnKzMQ5KafemAiFSiijs/7IvB99BDTTXCoTYwZXaO86hyFy7esOL
8G+bt9TmZ71bkdmfOB8XNoViiMJQOb0h3R9zPr5dGr6A7gzGM9eZ0nDbgisqai5ztOi2XrxyFe0R
Q0Vn7pdPHTlKUZAxCZQyq46/D8pYdPc+glW2OX7KqedT3J2VtKB016P8zOB7LsrCNVXOynuCdWHx
mZ52uXby5j+gxicq9mAlDRYb+HLqQ6LGwf25gxZvPb3t1uJR4WF/S70/CT5il1XEUChpteJhaHVc
zo78C9v7qqwebgHX+PxdBSCe4h5zWndBvqUpnbqsWuNWvAwk5rVVGcOrW2ien+NQKdkIxLQLPRYM
cOA6pc6suPWXdI5Her2D/dzdyS7RL5oEdd21WP0ykPBo/afDPoxK8ZoajB9RcJEglvNVG+WKOybr
bgqkcR4qZd0glHhudXtzjaUZ/8I9tZyqN85m14qIq8/wK8d3E48Ai0Bd/Q4MqQw79vk0qR8Bg5Mv
IBVWOJVe3FTsNgAEYmEd2qJW4OlvS6nzZnaIhWW7dlo7fCbXu3HPvcuKRsf9VLp5+CFnNw5UjD16
yYIR4MNgoayVu57SZDYHyFIGRvr53KK0pri39lNRp3spAvawVrnwMTgXEFwEDf1DYdeq3RzXlF80
G7ThV/3ZDUKutBIzt9vw+nJJMEyfw0nZNVvdpnIQl3a45rN96e5+5kP2cnvGgCWarJEDxo/ZI0JP
Fj3tau8VySbnX3NjUmsj20efDb0gw6togRhPQptGOlw0Wc6aWOiXKeL0ti7vddeM2i36KDopxqJl
NNTffqG/G+brLLHCRuuXcjfd5Agh1z1CFEK+CHkjWVk1Hr5Xzd6XzVieHUIKMMQ2TbjPYvtY1iev
nWGnFci5KPNqjfgaPg4WGff51WSn4oW7jCuCb3yiAHSD5A7AxmWIafTw8qteMIXa94QsarkG/xGR
y01dws4BFlYzgDi9tkisjLhOH6fVucYqKZCboFPL74/7OK4fP7741d0feVH1cdRCE2dHmhCb2+hq
H4pKiu6dRMxaZa0AAoKk+K9gUOr6dtz/MeCjOb3oGjbq/x8EHrj0L1IvpMSn3nE5DPHUCl4A7HBf
qfIsSrC/r5+mFc1mZDA9lAHA6dluMvLGFroSHavgYQRicejkJJ22YaO6ulPAV3K71psT8jcgWE4s
frZqMvFjq/daNrSXbHCOS9tnK2fk/eVYSVbWQgKlCRKIZmdBSUYCS5t20kMTQtf4+QEhipabk0ZS
793Qj4XGuAA6q5saFUGyYLjeDht/htz3LqW+sCr3JEpMMFHWSUQ1KaDZgUBZId7zhE1Hr58bf3EF
FErfioYcAhLpUJ7PKIz4TOK0XNZITOmdAgijmKrEJGHMpgLrPkHgua3z4UYU7/9XxoH+npimpQm9
bT77+f6oeWYx6iWqwKqDVWdyg8AX4ViKEA7+wpFsQ7XuleNeFGKADCli3mRW6nO8WRkbykIIVPPu
O4UWw+6tim0+/ccf+Vil1B+3af9d6REjcElgVNTuXz5DJs9k7fw3KlsxtDcC82RYpRN0QHVW6VIZ
+F4FhYoAQZN27PYG2YDJSkPIacpM44XfwpCPGxFMdorimt12ls1X0+ZWwfyt0731FjiLtgFNSI25
yZQUa1ZQjrb6d7Ffa1zKcvAaifQhuJkQDxTGS+tXox5i9W158gNxSbGa9/czSl9acHbve2INHxMN
cFkb50SCqlv6mFZmqn8wfnZGhF7nhp6qteTsnkNmtoG6iJND8wvfqkjh4+isA4LHuvKPY/9UybnT
TVw43wqUqmdv1nUsFT2TIDaeDWdWjhW2RL8uvn7EQ0mPH4CLWhvKGBufK3FGddL49l1/ECATgxws
jcUB0OS7hkwuBHp0Q31sQ4B/8vhrBTmWDFPC3qIT/H2S0n3u+Wnsgz8/+Xyc3u6+rDct7hUoqACF
eUZd2sXQ0wFPjryxVR7YrnjxHtx8N+0BW+53y8ZfE9yasMCYHvA0bKrVZrjTY/EOG7I8l5qUTWVl
5jko+Rq/zv4nhGhny7eGvnuccETHnci3tA2hvt+AJHpIpKZyIZke1HNBNOQMuwq28A5hKehJEG8g
lIIGavAC+uLLTvgMTMg2Hhopz7uvgnHORBsuDewJ2UD3LDQ82h3MyqPSiRU6uetLfsAhWrC7RXbO
Bv2+CMvDNZd4SOGDj4wF1qMOLH+1jnOTN1ynHlipkESJrfV87796L2fUM5dDicgAWvv0gtJGXdQv
XszyHG/eJymPrmEXzgjrqjamc1Y7/5fMddVSvganr3bbLDH413N9l3OTDIARqnw4Zf3PFT4TSR+U
nylcay1nCUDr7lWPe4k+y548uSSc5SAHklgQ1r2Q3yqyQa1EMHtgE6L6zSwJ4xEt7m5m23ZgbDrI
tUTpXY2weh6vZqJcrc9UdwNk3FizNze1ANhtgwDXpq4BR8kkOMa+4FxD8r6RHml54tjMJfUFdiXL
8/FZXRaxPfMk8fT05Pdsy7awBp9j83gfHDHEZGKpLGHRCjlbTV4zcajvXuw5I8xAw3TXvU+n8cfd
l7tr5a8xbWGKKVsHC4lAIoUP4E0OPRRdaZkWtLOux9l0iCUe+plHC0AjLV198wyViicHCz/XkZ61
KR0ucz5NLE6qBIWRbaSFy+ysye1l1RFkoz6jzc8nxZyhtNBrRQURWNcdDwM0UpC4HEzFgaK8Z4WB
22A45n6gRcHVNiBvP4SUPpJlea18hf6BaOZ863tm/vqNH21/Qvs0LgGH7sZR36tXwxZoYxSqJ+0B
tUwTdmUQMRdkihCc8Yv+Q3DxGEgBUaiRjCHhxyH0NgvPvQbbY3dQmyVPKAX3nJWbck8TlMEvWhd8
qj0MrUGui4ipPFwIntByx11tObNDToBHAPKyKxb57Xp9mlExblix7/j4sYxuso5Z6G4pd7fy/LIG
/YExQnsT+hbRPemFOzEHjG49We1UP3rQ7is8fOeuuYq3/RPCK03EOdCh0Lqr7T3Jxt7dMkFYbpBQ
RslfqVlmSUzlZFgpoMQTi08Vj+O2zNQvwgRHRWxhGiUhUMlaxcpn6SDdhY1mPsuChibkDL4BJddB
BMunz10Ckdyy30E2hZ8SK4ZvUA/vMN2FgOkNu/9HeSb+UDCmgVTdmwwiF4lyhbwl7D4hhuqOe+VQ
W5GpRDgKRowtzZfNHOJ8GUiGvM+GhQvJGBODtqF3QbARUTaz1hB9QHg+njdBn5SONwsp83w+AJfd
6aNcfCJNbwpuMgTxFWnWTuGr4q4Z6hochmnLxI0oDgUfOw+moZB20GSoMfxrsSJX7GXmJo7yYXmv
4TL2M6dFNY/DsFKImlUTlEpSFV3jE33uwZ/m/GAyZpTOp8T7AHLgaUFD1tf7ZlXmCjwfkAVMvSlA
AAZ43Jk6ckBxmm2NAkBI0hnfkPWsjVFwy8LfsItpB5BrIN7jJ30PssC/+u5Cp89+1iBiep4vjoRs
+GE/R6IZWdqe9J5cMZKpwCZPzQvBw5TxTEV/Tkvu9qRoW6d8JVNd8UnrLEGQxIYlIz3d0F6gHGSP
s1tftMCzGkljrO/kKPl4T/IcoZ8Ch85Un37Zxx0Tl8zcYcu5PR/d+hHHuMmvvNPEyj2gcnCbfv/M
Vkd1jwWayJr4X2htGemHf4voQUsV9V6v4Q0oIYrkv+GeIZEGbg+HSxBQJ1l1b242DS8n+PLXoWTf
yjUdjdUAaXWldNF7I21xXsTrqaA8gRGUjkJCkuozxULcdjiD0BKfjRreQAlUa51qfHEMcohsX4YF
CzkAw9k8PiIACKa8WmXKFPxtSN45l8k+E3ZqbEVuvEsMv5Nig578+orqXQfPid9RQ0nDFRItXjtj
c2U5ptTOrnFTzFZlDO8QUN/bvj/Z3zBXbH/ozn529c4Pj1v0liWxU7xe54KTKVhnqBaHXodgmrLp
eZVviMo6C1iFe6kLM9lC/Za31bqHU03aQzO1nAI3R3kq0y8N/cH/1ksN1L5STxJhCbO7HTv+8Ufa
NOlOJnzocopQINCxQueZgBrHvy7fhwqIEJf/2cj/yh9miJJQ34nmHFmZ6rXtVRQeyaLzRcc1ourG
/QzLeXgd3UHI69Al0mzhyE+BI6/BlXy9LLOu5vN5DHF2Rzfo4a++p880u4jTge6KOVvXEiHDZ58B
m1qEpxE52eMf6r32LWxa5ngTH84UUk6LKDDQAQFMuQTcSAhKYIeQkRC9hovyPSfgjXC7JEuojsTn
2bJu7B1TjY7qsENGOrUFmY/C3he+xwiASAYfbrA04EKLSNxX1tga5TpSehFmOmAYUTku7zffWalU
AVFYJDKWnzMV7G84cVAhFIdT/114XlURbtawqCt+ydDOOmMgM7YZ/okTnl0BctiiUk3gknivObiF
/cxbZ7EASsZgy3nqdZ2cqQBtW6/YxUOCZIjBL4VeNxhUtEY//EcdsJ8fLaPV6rIvQuLry2gdI9uB
AA71xTZfxr3wN9eGRE+3mGnA/T25+WY76CczjCPOG3Y4Esy2+6mqr5rGH07YQ92vB5D2gH5Q7+ew
GMI+oiAnzZl0+aF5Mut3mLnadEtpQ4szKwKAb3NJn+1BmT7aTLvdM9zDVVvTUJw/8IFP7TbeCl1m
OtwAHTpdq1Z63zhkXjlVEhZm22JC55El/FNX+90e1XHVdfiJYK4xt57f7D2fKj9k4JYgKcErgXD8
FRZn1BY/YyLcPKt9A113w9DomfAfsmcluLRW/dfJ1w2Luk7bgZ0VUfmegdZ4KX91X3FBHZs6r5KC
Zmb6e7Cz/uIXF+xg+h1hyQLi2ChzaRtKvsUQ0RgFa95Suxf79TB+2i+Z+9h7q09XYAICea+fhrYR
QXq2+mFSdyv2KLER4kNb/2Mt0CgFJLrgLZ8af1rMYQ+iqmmt4+PWdcXaQ6VZ5O52jeB3LVwwlz7T
TZVqhkhGGoE9GDopk0wRmHQo56XQBmBQ0RMSgoSMEKwlSHm/2BCt1rh0CC2mzelI5ubOBze44TJd
OW7AJLxRS7hh44n46AVovUu3hxFxqEJo4S2j1gaBHmjaol4/5sMvoew3uVsmEShclsxAs6l+hDXh
BBH/1LdeGwmiYo4i18hoFDmcXERiwfppMReUeDYKFNVcFWlsKvto7+RXUAxJu0rZk75aulmpCi0P
YU3m+11owAQEBTF/ngT8+IIJjYE6tEMrnFn00tA5rTSJ97vgrTV7bBuyge0KExkrWMnrJVLdpQCd
uq3JovNw+DA0aVeNUJCk0kg5oNGOUgBF9UFcvUsl0gH9WQzvl9mdzCUm9sv0D0055TR9OrNsbd3j
nlbjZHadh7lCmTzY2+UxCvMdrM53+hcGJprcn3FUak3sf6orwiOa90n0BR3wyo66CkNWZm4CUmU7
A6fwwL71mjniQVXzo0JvAx/k/dQKrXEQ0z6jlBMUnx432QHkq0EvOyKfwmCUgJxMhpRQgHFwwUkv
Kufz1M04RC+f4qfkOhBj5TRsbZe/Z/oJ5XYQnxUFL6pL1NP+W4QHpRDeE2Lcq8StT+Ibasc8rMlV
6TLnxQc655nCwUrljk6a6EqRFIaWhXj6p35Zfwg+vOSmsOHHubp00VlymWMuaeUW+co9kD27HVqZ
QomhuJoWIp1tho5WeWBHT5JxbzsrQMRNuvEjt1EhcBxITzz5aeZoc0VCF1Xot8DiHE0v32NjQo8l
joLGWZEtKrCu3gIA8GYstXhRxoWEQsziyujce8H5878ZeIle/Zl95JlnmwmvcefRZ6JS2WgjKeLg
nRa5JO6TgznpWT6PCJnLxk9Ii2t62iX4YYGsV4yQi0ed2Vu423K/OnDWJRIyrnRMYutBz+XxIHms
1GZb2JaEAL+B64aZSvAdPt+X7RXpSw+qLiVwr9XRYTG0u0bnixtkRJK1GX55QVl9TwWO2vQa0BiV
7iZ/uTdGFw+jYlmIGr7pvJd79WMe/ut9qQv067aekkCTE7DCXKALjfqhPZf/kSAy6pOOx1w0RS8y
i7HagUV5ZP3bRZyB7UbmQp2GhWnUdswoJyqDYzmNZisBTLYKLvDWjhK0fJTqgL7WF97U4UsVTeQx
+kRlf7KGOBFUDMbTS4nr3delcsmfawFMsUOtVmlQX0rMTF4UzJH9WHTJZeki9qElT89ouGDQxJVX
jaRFndQd3YShWUZuT6FpEzGrSr5U/TNyA6Y6znxlFEbo6FLotDQcqcoxUPPjpcHWot+Ng7TISi0b
LsxffhBtbQaQbh70cz/ajJqVJz0p6OrB8wJdsAAv9rSlwb3PUgQ+FVrH4vG1WaVhg+ti8BhWpLuM
z8G8zekRXVsPdqaPzwWVuUJPTOww0vaykr5oNlz6HLFZ4pymAvGi6DXk7xY+YEQYvahRLihoGfgx
rnqncboM4lM/apmxZC2Fz226YFBPZ83N1o5Y2oass0HmLGAlC0Ob87FAqPQGi6xqtgQ6KoN6+gaS
M8I8MKEtVi1P8OrGOyoabwZMdtzZvmVeZX/ly9JfFawJ4cjA/cgZxnGZ3W2xjdpB+dNuyCrXZiHQ
DPI28HZf6sLKuXfYI5aXOrEiK2p8DYTTXeEAfiJL7truWt5olnZxgfmoMJsEPlwYC9z2FIGcfvSu
8Lp5HIA6ZpB9gbUexg04orLh1CMBp7aC14luL00MaBKEJQ+HQdYtinBdt37wEU31HRdImGHkloe7
9/MrsPPfPw8avgzB9RlE6vRrFNtAUNpA4aQEb8RvU3N/N2lHXyl+6DjtvNHLZF0sRegepGxsNOR2
ijX641TzPeS7Pf9g3Agkqao/riIUDYVlVY6yYWI/QkRTEZSFjPoPdIWey4l8nXcg/E7CAy2rgpeb
5VjLHoRiPDKUGjstqT/plWEYg7tUG4HWR5zDgcY3DJH8Fwyfmmm3wapEWhE9Pe9rMMRWhX3jfD4d
66GaIG8RGa3tLHBsvRvTvp7jyYaDtBhWU7vRP34ji9G4RfCXBLtwHUK6cQ50vYx4rfh9cLwZthI+
n9NsxjDH6Aqjr4byOcQc4k8HIaW1xt2ilk06YPGjpenmonHAdqKs2D0l9rCVjCg1N9gbipV9+/C9
3prii+j9Fh6aqYFr3akT++N+r6d63XcHV1fNq3berTYwBLmcnk2B3CaaB5364t/RytrTJBGMr3gN
WCYuSx9GEzi1tbLx+dkdsfcgZ2u2gWSlXuiXoQPEnvy4sPGhbTlJSZDyh/9d+zeyACPtS5lJXrET
LpSINAuLTV7crvoE2KMIjJz0V0f5n3mv7zSTTFCQPoodvheY1Em2OXRVyaXgkI5hjhUpxt2YGEt+
uhuloOfakss6mPVm6g1j8ya1Z3b3qpoNBKGTyX1yVuS0YqYrdn4WIrU6r4tXp8TyudwH+NQE+wuV
c+ORXyDljdYLihwYKn8OF1X+2wSuRE5cUSumCMJ5rou43zNjUpTt7A4EMXQ9Gqw5+iykcAYIkGC8
U2SpJ3Tb8ionhIoXzSut1rQOxeb63s7OLyswuhBQIjRDs2M5FPkLcUFSx++RIFublJpk3dPh5Dms
HXDFTD8cf8/Grq6uttItZteWX+Z9urtG3goBaHj4qdIUWNL+btxNrA25mw2FomSN+PaPDMtMp8wv
5V0pdwXb4lU8+Db3SShUQYj1fu44vneE3K95ugn3JP8GTn9yRNrdaGCekqfmwwC8dXuW+SOUgmtp
LD+CwxfQR6yh8KwbHZQHi0WxC0FGRkDFzjqDORzLSVvJ1KZVronajlalMVGBpwu3kvqmJH1wpT0R
DeTFZkVLlj8rZEufDy8i5y8mdy5NapGp9qr3jzoOWW0mz/SIQgz19yMedLO1+K+YdQeFvk3My/NO
51GZN+OGyA5cY919pw9Efnsll+K5+JhJzskpw9HdwW4xp96rmXP8SCAIiEV112eW3EgKO/+beFre
KmtRPUGXVIAQ5lqCmPesajRXKAIUr+0EvtOBSK4KH9P0J3YMVZ0OtrCoE+6m89YhODTVsN1/RK+X
iGDSRVt+Mk82f6rczmjqDbtCi6sxkHwqnA4KJqd+CvdagjawXbQhvT8TVB4S+vfygiU8JgutnMs2
kn81bYswU5v456p6R9mqlnVgSzzfyjE3vbik09U7VjwvDobTaRu5mSGtBLbvz39guVVKt7ooUtbs
1LLlzBmAPxf1Y2Q4vJIDDOG5/KJox2cB/og7D9BW361vpJQHawtwqlC5XL4aIx15tL8YfsEW7Ksv
RRU4t/SAJvEBrBW8OeMGjXJqEJiETY4NvZix1SLgAxpksNY38FL4rAPG3S/MSgJ2TkfIZP6vBekB
yCInI1RZwWCuw5eC24xXs7aj5lRm3EuOLhV9E8SRFNVhmAAS4gavB5glFdoz4NbNOGCCUXUErCrx
HRukfIVjnSgbNj8kdgh0uplbC1WoyZjGntbye4X+nz0tWnKbG6RyKXJi2OVuUVU38wu8Jnon77vA
xyN/cUqGpdq/VjIuHVoIsSKvlu04OzXYtqx1kBFxb6Yu9nLh97+I6ga2iJC9bFjxg/+XzPvgZiO6
BrHLsS+QUSL9JaELJvbNEtnDNM1FYWae78TgbFfZAEr46LtPb7of7nNRO9CEvJrNijHOE2sDtcWY
fZuwkdlmebPoNnIuqIPsAhwbNMAGXOL2rrpmYdziz0t37bajwZfbD/HXrf8SHaOy+aYjCcoJTYUf
0AwFYqxIhDRezVIzwOhP2iBg+Fhl7GDgdVpvu4Qi+HFhFwPjzwv9+WKN8weHJNjaVJ2VY4f83T0v
sMGqheq3maq8JnXHVF+soztEo/wjXX+H9qfwucgPf2r6wqIijAc4PKG5/GM0V+binOuui/9g7xT4
1tsKpQVM8AvSptGRK907Hnf5hXKqttcSx2ydNB0ChTBrgMHhu5k/XRNWDZji6IWPdTWtvzqmHgaW
hesmkDBcsMgIT4v0UFAe1Wa/PPf/UXyHzGTW14NMB3LHkvJSbPQc7usPyOVtlDdYcsP2BcdbA8dX
AEvZvk2MWsoiptUx/IocPnYA2FJ6Y6a0HBrFm+KQdG5zfdGt78GKFicCKr5kJJaNTxD7L5Mg4Tja
PLCKUfZHEYwKBktdL3WD71lpFnK1jAJM/M1KISGNb7R0VL6MOVcqvfaLpFi/S7FlfpsH4ldw8j2X
cHSWvobxcaiF88I9j2Kwc1IsmSG5WS7zEH4MQpe3cC/mC9ePcUfw+9aeVig5uVwHo0KKIVTueu0a
M+BS0MPlggjbyAQcdFvEZLJGmVpeXya4NLTuWdb0BIkOZIiAgKybm/mQI29KF2ukVEvHYMv0M3kl
/OaUbWxrsng3SJFAVN0QDiI1TUMtGkiXBD1o6oqQY9jTSIWpHjg2dqweEVldf7WaYD6UfCWZdzsv
f4gPOOegBLnpXbbofYjgsLL6Q3dXWX9aeNWFAj/6m1BDV4AFeWMScfzIyzRFJHfiZ8SJwyrwK1Sg
jz4e+TWwFa3vq0mb6FwV0NecXNNzla3M+kv17eIH8hCYhoCOYjM9ROuxXp9wI8xjlJdPRWUK+LdU
pl24dZsIHR1tPujz6xtU2QRf4d6uhtTZ3JgBQd4A25vBO7Xs7MJ06wFuuV6gulMrx57kRRM6l76r
ZRq3fEOxSDuya3sazfbKQQbRHjFx+b8KyPtJF9XbjCQvX7lWrN8eGrT3uZHrCOyN9gGKFyfFqw6D
OcClLy0QwSmfLtrDJC4DQmAC491lV9boqlrqdLUjQL1KKW2RyI8gjPrLD+tbZAduqBK2DX+8LMP7
/TkMsTtSsj2h3pdie26l93dcdIq/EL7H3RLWoToKnLT9gxFnq5Yp+Xe7WcjI+d2OH6lYw8g32cUw
1hzejpm+LyxTDtqT6Pi3fB0Q224N7SfXKzl6/AJhtH+lv/IzSzzaSiphOzVWaRyF6zVuABIisRuW
ayASaBfiPPtX08mgtvJUzQQWrq7l9WoxIq4/Oduj4gpiF6LX7LE5Hu4G+8i/jyfyulrjvojlSXTe
OspiNSnxbnshfkHXB1OolcL5GcrTDI2flSNqk0SEOghxxve4UQ/0bHnRWitvb30MiGjjB5Rv4iPx
QljrBDqBL0eLdg4ccAOb9xIvJm+8E0RrIBuY47RGhVkXsfuoInhsromensJAe2ti52MYfZD/QkRj
hrZO7msmCtigLUNYxTKuWXE1BWi4/DYwUGvJ2xLtTA3TY3gmzFTf17/QXBJgCwvZGIogqFe9B8xU
v7nFzS4kEe8KKwNY9b32zWz7CQ7spPvvBOqSMz+RKbahEu5LekL2IsEutkH2Sao4g0Rj6YEK5HEa
k8s60M4ZW7vKxhlF/BHBRBwFW98fzhdXOjJtfhFqf+C3QInFtXRWKx1cMNYlXmuhmmZbO17sNChR
ve8FaLOg5g/1wF6IWHadWO+NnrUoyPVuLosO+ZJT0cwVpDJjqXFlzCJGOgi1AOCmkbdgTasiJE6q
EoXePQYKxbKngLTOCTuPjlq7o4PMHgoQMiune5ZGkz6DzfHh/VDyeFEvlPnyYf9/VMoXzeHHLiLi
ymaFqJje53IHKXWdbDuwhvixbJeCO+C7yutWPcg8JEYj4QyuSkLN4DOThvAOK0AQ2KnPd5qBNIf/
0eep1PSF01TXXyzSP4mRuiqimVUXH69tE8E+cUV6fSDB9GQs6x0wiy1dSPpFhn4NI/1B8t40HlOf
mKf00VxkZmrl8znKay5W2s7uUCCiHg/P64I+pI3etAW0C77HksgAZ5GxpVJmxu0cJEwzBEl4YVZK
o7Vejp9ammPCM7ai697brGizEfRgUX3S/Ex6MkxhI0YOyoqEgWlrlVwnt6RfOFD/8xg67nOFn9aJ
lbFObeABEsH6MGCQt98n1jyJzJvHXQX5YjiLTCEbED82CpTvX8y95urCdFAl/PPAwNyY/Hth/NMh
tWvuyI0WH9kxUjIrBv5PDHDxV6ay6Wb1ZDx4cGlK2Jf+4191nMaTpH9D+jrhM5EdSm3Dgf2cp2K3
Jp0GGcxsgtgoxlQFJNBuhjogti5oYlW8w8PZBap+m0qcl3UgYdlAJx65a1dvV3a2d0JHg6Gt6l1E
2NsI0LZI9v6w4nu4sf3KPNBu4HzjdWJEpUXO9mf+yHki5Vwp2Bzx3dw6aBhoCCijdmHRdIGWUgTc
IuKTaYqL12lTEyMKU/i0DfqgR6XDinFfZgkqYxQ5GG3ARllOASpnIq5EWVizeyWyNVWcE6rhsp8t
c2aJ6Mivyakcxw5+N5JVIcjwVARqA9n8HpHqWqzkiomNJn8hC3CFVsP7lBZw6Qkk97NtKDDPAnOy
TeZRIr/HFFYGBLGm3L3e1WFbtbwOcUlkQGwcUKSDwD2t0fDeMfoIgR6YCNEeUWZVavD8PgE3WPJK
FpopoBjX57XrGBNt2vkRoi0SPm1A3+v1k4l5scsxGZqnklk0C/veqVo1uKhhr2TdbvPaPEvsFqL5
wpgI+hGAbiha+Gste/4nH/q0vceA1K22L+J9fG71PQb0IooPsimTcXMdpQBjwv5oNZNgF8RrWOCN
sGqFH64KmrxkHXxE3s4iuadSVBOp367UEXPlJY1eJi4CQtQW1MaF68nY9RCFPhMQj1T2QkVhNBuH
7nkBGG3/TPQHkNBz9BE3w9SJikdioEBuL20/RielfzFo/2JRasUtzABzxat2AsoUhCkMfh3ZEkvc
7fmOCh/lMKADwxkLiHK/uL02AASVmhpESdTZe8VoaJi2p0Qcy7vguFc/bfOVeaSkPnzBTAdgHknC
YIxR7z5JBi/rkpaXuwzO5Xw1r5JbUNzhZKwSlTj3RzUgkbBLsYLA2jIxEI+sA6Kw/04UWRJHfNOM
pvM2ShKO9ngCrnIYgeBMOClif/KJ1zHUm762/nfpakn7F7QBbs8HVSeBG2BQU6Sa6gho9UL3cqmp
EQvGHE66UvzC/xLC8YFb4AKQx5irBBkMGYt0hsZoUikSllIF2EnMnrxeozBZH6XyZV7s7F4CMFAY
583yZqu0Q+jccxcZ2BoZfDMCE+iqLZ2N5GRiHwT4S+My5Vc9nf6KfFsoB528eLpVAbA5Ao0Hoh75
YbsRrbuPwHcA9W0RYmYXgGYd2c/RSsf0p9iMlwQ1FvjAQopUknoYyuzrkL0NExXF6Qa8nb8RzTLZ
14ynggUP6yAp31ZY9EU/d3DMENR0x8GcCEdgcmDTeDZQ62dpo8/s4+kshej9cV2KAvFClO0V05kF
D0oy6OFMHYGzBFAKtH13TL0p36zxJqZ0VGka7XXKT46gRzUeKrd3kKOZmRXM66u2ghELHwxR1dY0
1CMYjiAH0kRk2z0tpcexWjH5wODsbOU+KPUcyq4Qr0Sx/MhOpHwzPgopG/pXhvzelsDJHHJjANLc
eCQA2bPGcLs9Fz4ICiwq0B+AZR8vlrBwXnFDRc2PE3SVbFA8fvg9I0NDFnygVvpjjgEYXzZekBao
lhXvgbXIreCEffY1EZz0QiGz4K/D9PhMbqrNzLttEFssC90qHyhDJMcV/0KhDXbMRVXL1YcvvThq
zQu1OrIJifbeuYociY7XZy7cEQLu+Ia/6LMhRD25cEZETrGxDBfzBQcUkbMIRf++mp4mDcgur1ky
s0b5tU7iFtss2lzdUHT1UGe00RVQ7QsY+tgiB8XNZKEVhDhP14Vha2EsOCu9zT6ePkkZ5NAhKu7L
xtRydIp/pgAuCiOPVOJhHb6tapb7ZqU9VUFX33FebO41BCveIUyl4Ogi9CkK2LKlMC1AnfBWg97v
TAqjXcUUjYya4z6O+USjgi8h0Na+m3e8WfHSk61LD/PJKvwZoMYvPclZ/uzVIRaxTb+55M1Go2rd
RBJrPk5eHx3LQUdOl1cRHwKu2dFAvqHJxfmq9WQrbp/1zaRo6Egdwbc535cLRO+DUxmE73jsC2C2
h6aK8wEJRx4u2dhTEBtjIXeTbYdxZwu3RvanvVY2gLur5LerBviEKRzZUF5TqAhtHQ7I3QhGQVPH
g0gBddj7l86WsO0H1VewNL7IKXKqgreF0WKHxemiJJcr/3yzeEpLVDuGNP6mNauAqgCz646oPSsI
tqTsJu+W+tRdGAbO6h9ShcayXznVgx0dTAvj5tipjmB6odayqezOV9vh8OykN5HsCcBmvcZ7xugx
CHBSTwWKQi03j+EaEjz0R2jmqdIppBnPhvf80vaa8NlC2p+N2VKDmEmlHyXfqnv/KBwV4Y/kV6NW
oEhnvdBP2O+h894aDungeUUTbzwKpe0l8FhfX/x3rOeaZgYWbRyDMEMmG+F6XJQK1EyVGTV9jX6g
/RGmvUMVoROVwCU3kgAfBAokbtY5gzb63CxvI2wxw1UMYR9RHqmURNWpVIzEp5RnoPP9g7R8BvnZ
4ePPP9I9a4ZJMgWH9r0MTsI4YFZDP07EA5PMlf3j4KnKy31X+JvEunJq8osrxM5rCXyDDp6YptFT
n263+423kenaddYbjk0Bnw11yZ/FtWEdvDHhdApDJOT9Ih6UHWHEsSLnQ4oJNyZIuYTwLz2UdCIx
yajRFgILkgNhHlNC8RF4m3DBetT9YZaXX7KFZulb5yXhDSBzOe6IsaIpk4YDmoTiKzrl5zK46ZXI
MWxaFq1aOdp1VvnKBePZn86wCgA0HqjHtt7j+v0tnNRPl/DEOF/9ApZ0r+3oZeISF/CuaCEIzFon
PtcxsxpFRbhfHmd39jAYbSoMuEfOI0/7CnS3XNas7QbfCSnJAOUFF+oYccPwTC/XSQzL8sTMv6li
XuSvRPDXUXwLf0jT7l8QNcKqLFZ0+6slCemFes2jMj28Oxq1el1Wcle85DLm8v3aN+MhoSGFDZtT
A1/h+8ZffGAol+gCCAIDpOiM49VkKCYQ4siXudnK8lnLY9ag6xFXmLIUkdBQ7RIEsnevXYCBT6pi
YdPZXRIkCu4JMJBW2s7Rf6WIsOKtSB2sPnECWKyx2tCEPz9LLmiVUqRTgtVXtZmnkjSyBq1pyWu2
nWNWvIrfxEKbyxgx5YRTmJzTxcD40/S0O398FcB+5dl8sISiG4D/lPo7ANLN3s4vTnCofq7yju+D
qaVPPfeByyMgm7cT3F+IDtanXpN82JhZeHAE7uRPi74JtkIMr2jis8crzL0o5wq+lMPTO8TyhpT4
3hXkJoAhm9z+79p53T9r9RjWa9BSipvNIThp04wN2aJHbeANd04fp5e9bJbaP4dt6BP/WemwaW1W
VCJqd+WSiDYsBVofILRJBeOmvVa+Yt4jyLEJdH8fN/ijlH97jeNBolvqzzYQ5D0lx+y0jB6PLViL
LSl08mamYnnXbP5+4kGe+TEt6w8ogu2BYxKQk1vVzspfvJg/9n3kQlq7TmqJ6s5kFkb02MbOHFxg
ivu3ZWnMTwdClXLUNVnMwa2THnDakYAWJuhiz5gn8hDnOXf4ldFMuZE4xq/UXSY6/VGgSdqsurHg
4KwyZc2dWrHwjnVAQ7u4FD7RW1u+Cb32wdFE1xQFn8rnJkXvufBi1+euRhJLGwR8X765ygbSRk9/
c0Gixs+APrtjL3Z1SwXzATCc8AFQvuwPjN74OfUvWYRYBWzI8ITRV7ejWOISlIg4TE503N8f+nXc
pngirgIM7jnn8f+6qjwHDmlruVqX4PM9agxixFygW//WMjWZEWO/amM9VbFyQaW+fx3UH4FOzTj/
U+EsHe2vxXUfA4cb+pOOwPavID0749NKukaoSOB5WFJhpkbSIwofXhkYSBkCQ2GgJBGP+eSp6A3p
5cSoJH5F+wsxTd4M8SrQ9fL7fD1Y+2IKOsHWLekIXOC1G2CWEbEXQ4dFkrkcg9PlNNMvdfPFnLls
QMHFaCHI35X32H7uz72f7/wYSqXsjSM7zuOUJoSUgEzpFyVSRRBVX3pp0HPkjP9EK0ZZbRFaXcZ0
HGAm2iorYgwnN8oMgC4zxPvryLbYgyq2W1k7Kn8UMuyUE8sZNtGNuzdaVzTfZeFwfK0dqw2QPL6J
+G0Vp/dxIFq+zdRkpBtYO5bPkTn9iq8Ov6IszzXNla5H5wzXph6spgLH+W5TexM5wT8BvHZQWUuw
qgK7Nv9hjdDJFvHy7lwxegGFn+/XVtWEHLtQcBzeoyV4KuOcj9DlzIaeFjm1/UknHyq+pSxYPA1u
3JXwjkjDkh+ssdrRivjsa+WWpQYFNPxzFxr5025BNOjFHUvX1zV4ySsOjLjGorgzR0e+NAMl8aiw
I/5mVlnT/8DC6NcgWCNDkoLho7gMEc53vQmQExTGcE78HgX+ikeuiM3/PlLlqQHYkjm07Iv8yh1i
VEBaETb2kFkSX2YGpq1OuQlqEHlFFZn2QZ2t4akYnPyrMRboBghuse5XnQveA/pJv++7Hq5sUgkA
R4974hdsCJZC2VZTbkR9lrboX/Rygo57odjw/WmKQsgNwXSqqlxjsoEPytolGhYF4jWNVUKR2T4X
cbeCQOoW+b7kj3Hq915OekfflQhW1jWeCePkSD47Rs9iw+9Ymls4hPUT+o6dO82QwBEzEb3hwEQ1
+44luozyNAHmrfZUZ7cBYIk1DVkbZ8oP3c06jqMMa6H1QpTp7JsptY0Dqp8r0uMWZEBWVrNz9rWt
TmxlqcfDUXO319qNUNqiyV+53itpWaWhLLQ+bheScIDP1nUVnyTTlol7yvDDYGvceY+45QZ5d5HH
OfSzzIfiZpxYy6nA7KlLHdCB8l1FTaJ6zoPdUp1SUu9sywaAuC5VMIvlcdA0qqeAuDYGaMkNKy+j
UvNXtsVzvRjs3iATv2JY7cTFCy12NJ0rGvuFAYUUR3L9F63SrVXYP+jV/jbNf5J4fnqpIvIaRyTc
XZADRq6YxLy7+A5TF+HVf6y2RpeyBwZ8MJqF7lZeO0RD5R5hejQtGnFUIQqUAD1yYLjkg30QvLy4
ZSMvleciai/u8Mi1HYhyIoNHfhRfuBgxJSFZgxgJZu7FYAjGQJZCFQyT3eP2WqkvWczNxSofJl/O
bjy4ikIFGAVX4GOaAadsuJjcOspptMU6yEU5/kpkCbVZHCx17Dn3/i7dmO0QXzZnYR29Xt0DmuxC
r+xHIOW4OX8l+uhJsh7jCBt8R+p7lG2wITcd30HWmmrZ87121Nw7wMM50MpTflVG4rxR9Tc3T3Qi
zTb0KnFncH1Kvx1rhQxw+EE0fvNXqJngImkSMehOgyuCeVqroU5e0WdBMT47+GwXeaHTlQqZBC1t
ihqM9k/FFnWDfMbzhtsgTLVzsTVG92/o4tnEP7rfjHQaKNyRrfl3gNwJ7nQpXMu89eey2eNL0iAv
jAIqL7mPQ9tkPvcgxCnCb5jaUn2zzDpVVMK2XXPgW3d+CX2Ednn6puL9P3N2I+ALyKhSgarVZEHS
IfsZOPtp3crlhNX2uANKMVHO2eDE+MYLmRzQuVRhFGLdPHFcp45J92W0CuwH2BKKFbJZhfQ+IVoS
aUcOAHM2RUPRb2IdUXao4Oqvc0+Fyl2DUJK59Ja4FuKuMaHRSQ+LC5pA9i5vbutvXV+ZWnaBMKnr
S1pHzwr24v9wyaCrB3hI3P0ZmIAhxtlCFTlS2B24IAq9t9bXBhLL+KVRLKzffpCpTMhZPy6aZ/Nr
0tKnPGjoKHDeacwBx16KKcoBAdi99pCxRrZyknNcvwsK4aWaU5gN59RDyPXFS2HPVgS/01GpiRDm
PNPmMD6hjeT4UdEHwFE8fAI0udj5DgJ/gwCtzx6Qc/6jJ5f8CYn+Q3zWFxNYeUrg3fGx5nyDqkmZ
viOnx2ORcj0s3PM2/7U2GN+DUMYJLjhlwWe4AZCi/5okLMFLlKTs8Nei/mFMcirQyipyKVFwWUlp
SszQPXYrpa3y69MkdhPZFoGjItxSnUdSJJURcTnRG4YAnaY2W1rFfVWcpuTL6Qtuz/u7h8scFbOf
T18MrubbvMDd9OO/7qv6mqb4zzKnk9zmzjmf3JA5Qlh/wUySt29B5Pgmuh/NZRwDdjj2wexrEmQ4
RQFL50prcOiUPXPpuRHR/E5spBXxcNfMDmYsfAAwp9jv/t2H19Vh0eAmJojF3aQeGlKlHGydKaX4
1CQ7nl5Qt+4zQrVupAqfcD3+/xR6UKHWHTjg1+YmfBAPlh3A6HvoNqhQOQkcIWyVDXzMB7P5eCuP
5ronSfMys0XNeBinz3qKWhjcZqe5I+9yjoknFcmGpTleRM8xtPzLfUEnCQLVbsRdrzmOV9jqvrZ/
pBzCJWKcCcIb7C46QWw4J9rgGtRQrUn+FR2SHgXAB0wUkYAPRnYOyIlJdY74PsXasDdwYquMxwsf
Mme3VogSl6/12XTK65kFOI/6DZsX7p909MumAgmycyvcqrTBtCr3NtMZJe/o+b+kM7Qa+pgd0l8W
qSGwz9mDRfHDVM49EhBH3AijAyhdTRQZhkGj7JgHOxlICEFKWcUqecN9xlU9AOzD4qwGk5FMmPzL
n91qcpKfDmnS6TbKEPGvwaTLnQHjdEINckqLn0duueCVXFgUEKg8emxSDZxXp0IVxAF49EMDLRB4
CJxypoa9JK0OT3NXnlV8Ehtwdn/hPWTu2OIsCTJ3ALKFTIv/tTetadfjq8Y//CQLY6ITaXcWXOyo
BRQPOU918rbuE3bq3jh0qvxUQ+yzVrSvpnM78pe+3vpykMJZf/mHt+MFCzSQlJz7LsOnOIMXpPgw
PYfZyDZhtYwJuIWGPybP5wi/+bpAuFbkcYNsFJ+wOyp0fclBhqOTXskNl3QuGr6xKIRDf7kZ8m+q
bpgX/rzGtM1IU+yE0CK2jjr/ATb0BCntoQ/tegixZ2SOpVayBm0zM2FyKHa4xgBo4a4+EWZ7QhFL
6GsKzirGRp9m4u8zfvqaA7jqwgLQ5F+fJgyWnr7okuPgMWlw66B0Uc745jHeSUsjr1saWnWQcxwu
TA+byofUrDJgBS1o9Aa6WXCGOaWK7aQ3mEKbGzHgA7Kij02SuA9yg6wZI0m8x00WZEgrx96eXJLI
elwOiq1pw/4/wEMbChQ5hfW3HC9wERuH08roDKD9WErickEyG+dg0WeegFvHNQgHqwxlnbVJWYPu
5Um4W6pDaScWp0JUkJA+n8ucgqbHidvGtQwO3JPl8mcRomp4G6+6x5YeTqQHn68+sEhpRQ0AtrM9
q4iseU7grC7BQW8GDLRGqFHO0VMLubAfr3lOQjbyHZWq5rwhjk5MX8YASJr4IGQVRfCzF5oa6/Vs
lJy0TcLR9Zp4m6Oil1RzGPtitZ6A+8su2Nc6JV5JJcLlQjh0GVtgC52pz07fbNn9LdKy/SkWZesr
JX8Gt7nZxlNh7UsUczrzYPPTRzcOc6LZIUxzVx8RdsM8X17N8Z6d6apZ5/Y9Rv8QnYszUel+2Fas
sgCkWOyofyF3+NoioktPldl8p2yqjx1f5PaYwKDv5YGJ5Rl5YkwDLP4S6Uo4Ww9LSi+50jOI/i8R
uOdYNkdWZFTOKd9d9cRh15mRivciH/w4lDOHGNryYxfKwBoVrIyF98zu8lKRhMaGw1DEGeRcbuhp
7Q1Tn66HkILK7sAvXZvXP9bt4Fx3bPo6PywIuLRP6MI81H3yZodTe5hebPy74tQv7XOuE/AdFBQf
WN6pU5AuxyEKaj1BeYI+eMX74xdwYCeoezC3DK72EKkoxejsASv8bG7ov/rLuvbQkOJsSKM+ThSB
XveQTEidGRhetMohsxjDSaQWwaULMEpLjaF3poCRN95ut7FVsvF9zevucnX/X4M1mN9gWzcOC+Ut
qXG0LHYDcPeF9jEUEHmpQHRphsT1qlmOjWTqYVPHQkl6cj5J4IQ8alZ9SI+YYl3NyU4FWRqk+u55
X8opkmsfSK7M0yQyCqXDm65wevtGQaEb/3nhRhJkSFlJayp+1EGcpZ5t0vcUQseleUBjHvQLJZDZ
JwmyZ0EoSirAjnQ/2dmgFsNT16Y8uCm9IbV4QYYwN485qpbfJEYAe61lZIesmJQiyEosx/Avz81Z
jISLMgrdxxmswR9TsNMr8s6QkzHy7DjtHyALALR9UdqcB7zOd1D2p8br7aNYJAhnPx1lKcUKOnPY
C3ctwXPuIodkfj5U+vxqlqjDZPovmsEgiLxW1Ia8mKN9G2wkgnrod9hR4euR8XhGx7UoqSO6IYpf
4taLrnI9buysAs1KoSdbxpzEP5WvbQgQHThSY19rcj6CgHaAyDI7gSKGJ5PvMA86yvbUntCJfm2l
SCNN7i2Fopl7WfIm7CXmkGU98DNmDr2/+UaRwaBKLHeaW5cjX7roN7Th0+kKj/69xOLBU4zkU+7S
oxv6GZBlisMuIUeQWV90b0l4GUfjbK3tGfZdyWojaOUaR2NxkNSNcO62M4OOyKTrVORi4NAsf3Tr
DFZCuwDTPpt0udqNTM5uqORrwjPjfWz07cBssFV9gviaVm9eC0HZ23mk+eDARl40ePhTxiW436ZI
HKUE1JP25Gnx9U7h6C0zCLr5JBHrIE4ZHcE/kOwjXSnxGK4y73MdebSNPonVGYrq9x3U4GRQ9fMJ
fKPrRXhbW4VIhKpxsJwNA0MVhPbWiNgCX0kzxRK1NISWtdLDc407f+xpW3EoojPfR0/eLH668Gfj
V2mQcAruaiXevKD3gjGxyDIPPQiOGcOoJQInTMbYTE6LYe1e3zEG3tR5IOBzZ/R6ioVpPJZR1N6e
TO+gXatQNSPHBS3ZkU3Py87n4oiBqeyO9f54EEFkrG85zMbGddn2IDUuXmffUGuD6QFAJOg7cJq9
nLPXFo/8o+yJqrEw+cSoRolDV6wvzvyCL5MqAfgXpl69jKidRbI1f2UlclT3bIneP39fbo9U4FOF
AgTsFL0rKomctTl1QuCOOlqgKAyu0OKIYmXSfeJiyUin886vhTpIH3sKX3YSYHC7IMSpa+Ro5lOj
CI9yBy1ugRBz3VLFPVPq/7zMp6yaAnkrmQyycOh9/QzzWTaFqTEseZavTg90t6659YaS6cdo1rQb
uB202rkqXxFrpnPduQ2/ukze0D67ra6+cKekSottKYzHJ8Vplzfl/bhVzAUEVFUcCc/0m47iFIpT
rLU7h1PR4swRJHzapG6f9+zpBhOSBC2NDIXUHpuHjkuIS58NKwa9in5i4ipFvPwkbht4SwGgCO8+
uD75mNYTv1dQ/yipZouPK16ysuzZ9AjUUGO2UXccmN0xT/s1WmqeSOyA+/E1Dk6QIdGx17ePyPLe
NWpqJF3yc4zDzFD1isUFzdYuV7kZsU5b6+dAXt6tOCYpA0RRz1p2z5g/SIKbkp4diBhCmozjjM44
H3krbF9gvUQng7ycfXYuyOf32ne+8yUAlvZB6tJlBpbzY2SMZTkDRUeWy5hf/7oEzHEG1quKQI6W
qn1PeugWGVuGnWsbiTDuE1zMggMNOfN5DcvHmRwZYpA9fn5tPEqjt9Xk64JVj8dEE2Iyi/Aixyr7
GaUFCl+MHT3NbnlHdbZ9TOwG1V/8nI8sVSzLG0TkZ+iO3K+ayvk0REuq0KETSwNkXEaQNndLuhH/
2IKFZg1VWZK2jnzDgVcR9UdANDB/faUgx7w+su+ULzMDYGIY9iN//RbKYrK9P4rT9zay5X+7NCpI
jp551ixfwtZg5saIdV/q/0ox3zh25B8mplPXA+AhWSuIeYG/B0d18E8g7SqsaHhI2pHNGLK0Qy6N
qaVC+3GvGEuMmL+uQW004vRCHiMbUDcyw01x780X41UXI6NJCalPBSzntiIVq8Kxl49pa3vHs6AR
m2gUHEC7LRvJg0AMF10/6r/S1mV9ZFCWMqDeJGOq1tWjzoI89RxnGKs6h8x8ed6xWSYxjiDpv5Ok
9O+JPRo4IpJWlBpcMAlwcH1tQ0YqgactL90g11nTFSJOSNH+P0sXV+v9CyWsxYNUsOGWlBWruTt5
4qvhO+7qmKcr6xgX7EAIKZVafHMe42QG0djt13JNqBMYCaav8nvQX2E6w4YiUIU57e74jFAw485L
lsztoaNQgAm/XiGlUpRRV6VYJJcpYLLS9ZK8vpXGPZyB8M4cL8f6l4pWQQsAN+ny7kxa6kqPklso
MAQkppb6syLs7uG1trhlUGzYTGVepE5RuUzQh/h3mx1Orn78CInCs1sCwuqhukgnAvWK0Cx0XZ0+
VF5rQefXGXKkYZnqzHvgnb/nFJmVoQCURYv9nlVum/Kf8/nof+XstAfgsoVMwFLORACjGeK46Nqm
kSkbloyQYY6gqOuz35wUDQISGzo+AoCca41mFgBV7OnXkZV0Po2GFO7itlBtTE/e9wsly0btE4tl
TsnckH4yw38ccl+BUb2AyNXvzepFAK0jb6ogA+br/TALomnlikGV7BjgMVSvvJvY3P+m+0j7qFW/
DjpY+lFFh9cEGvxaoWdKFJfz/R0zXWoOTGbIykDvn8fIFywDrHcXDx8EZoycF4PEorK2cKq0IWTN
DGNmIaQRw92OD/qZSIPE8lo2EkYIpR7YLjgLq+FiS+ZwaZM26vnMULneb7b9brWMDR+mqZCbPmwV
ity/6Wxr5sRBTphNRkjTQMQQA/eHENAfa15lPdVnu2VPWxpKWdw41L38VdRDj2gshHSPoaNS15ym
6U8SRYjedy+Su5Xj/udj6uGGtgYjKYqFIHx47k0BP2Z4cAAuI2OsxBFHuOSsNVEeh7nCXgN5mwuI
Xizvjfyt7GCrq+XSJY6M0cFm6gjID48IE5z6bGhv81kt+NTfJipV4j5P8qlhHBdDR+CU9oauDjEf
oe5VsRbXc8/+VMUvAfSfVeuM5wlgmZOYvetp5Q8cIs0C48X2iDi1grvcfgGblI4FHtXQwhGtrIgQ
JGn6mTgaGxMRoGeaNuxgHl0Y7qtzo2imhf7t3yyNuuewPLsiaGWCJEWN3d3fzMe9SOA77UV91Cl6
mUu2O255GBKQIcYiNxJQknxNshc+03yK58Oe35A6PSslqJEZJuaYucbv/58lCCTAFaIbmd9VL7EM
GgKUO7QE4ivwkq6H9kDk47mxHT+eqRlwogUiwv0V7XX3un8pazTl/dNtV5cmkZg6vy2aX2RdxoGJ
fiM6QDV009nOCaoXmPsnOeiupFx7TUqbfDzqqqNtQIdtzO7EUYhGl9BzpM6732stVy5cIeKhSj27
Z8ldhxpATsgejZvtZJmBzbtT2Qch8jwLdCc451sh+NdL8229t8jwCc6qV97neinpFCMyxa8JsYMF
6rkTtI6WHYNfn114QxZoDM0NXuMkvmHjWGo26P9s0Gr8WrlB5Z+FogVL4qQmmosZi/JIQpn9MRBL
wGDKwQ3FiuRW1ktIL1rzcBzumA8iH5NJ6a/TH2d5+GJdEBvvm2fezfSUEecyi6qHY8GnAEvRz5Be
ta8usJMBjqLznYiJEgIopS9b2naVg+xoEwfsHQEUaMtbulYOBU4aquY8RjrcYxDv7ggDFgtGuA74
7wclBMDJkJ57sZy7Dda9NcB4sgDEASwL1sBSGJG8oCqXiAuRK1boDc75L6S7fmeVtXLqwPcNhfyF
AERZkmXKeaFI7XnZmknSgpNvSuOXYg9VIxA6Oq7Jk5UX1uaEE3tzd+xl5FD3YX4T1r1Jvwhj2QhS
FLdAwsReVsSBUJYhD3hS6lMZPvuTVxTJCD/fC5av+b+yBg3v0UOZHZJ/3UmaN/1J168l+xFigx6R
P3nY9kmmfxy/0cQf9pcGYKd3rq6mB4zqMOrMJQYhVBTQur2+z7GUMTG9PJ2M4HMOC1TJE5Ztx272
ugw9/xmTHJwiwv0+7+vIpuF2XWxs0UrM3oG1rihLUA+UqQKb+DBLAQz3BsRzvTCXqfeFzrGngjPH
TNdvmfjsbS+AdByFvaw3QUDRa6C1t71r3s4f+IpVZ6rMPsQ0mSU2HaX88AwKJnlGRxYbTbX+dehr
Tsmoeyq3BLy40fSF5b+Efa6n0eCjVgmbg2eRj5RdXC+/8URWl9lasfVxDmJbtLBBfyx42NmdkzNg
5CDYsIvk5GU6G3EEPduKyX4Qsdw8yG+Md1PFu0FDa2P67IU2A7Ut8gjE1gW9OFedAjIXMv1D5VC7
tytK5SInM0S3HiLovVvzlB2mk9nftNJ+hFJzQFTJl1dzvj2Fs7IZlkLgfqqlGTFQz05S6DWqhq3a
zei295RmB72XZin1VIvchtwQqvgukwNtAXZ1faoNP+IpOy7bfjuRhMHI2UDuzJEE257A17z5x4mL
iN4J6Dc3kF6iMpmMfvaRuXPWms5MNTBwUtf5SvPOXgAPz26on+b/NAGSRvQ38g4x9jtcYl2KkHWA
jsFA9771RgWwbxiHes/rjhw1sigrX2l6Z9k2+YKzC1vIh+oXV38WII3byMu+egIgJh0cbMNuBypH
jT2PX0OtVDrF81nPTVCAl55+0UF8yQ+00m3khYyW2dC9kOzWrAlpqpjdtDuG3Cx05SlpqsY+2TNQ
zWfly9bJtkQ6mLmuPiw4E99/7bSom5qM6pyiiM/7/AN7DsHJYA38Qpy4J9EM5u4NauxkI2f82WKW
4Sn2wj8zBc1qPveX3OljoyQ9Tt44pNa+mDPc6uR+JtU4hOjG9kdzLZVCBYqqoVncQE5sigpTo0+i
as97YWa47BdUSeDn6OhYzK/isp+vQeT2pga5R8vXF+Ua7aiPNhDRrCub3VdffVCYKJQY4lVCiO3e
s67/dGMA8vALyHedAQzpPgwFmplUhR4XdDQl60JcOwYelMvh/9q3M8mw7i2HgvFXnrbFiZu4noTX
UyswB941ssEeDNL4CMX0z7NYlIiq5d+T0x10TProbWcpUReU0ccctod22xFMJWU+z4XLHDAAs0o1
cCy8O+mAJ6St+VvvBpuynKAlVCH2m3TZnTQVFPe3vRjLUiRTkZLipItW3sTku9zOXcOcp8P3Tzri
/s8SB4TRaSxHzol991zI7AZBjrVhup/LwHN5EJO15gKLvQpeUh7qYtceKZ5kFiY55Acmb8DVESjv
K/5inifGhB88MP7S6F/86RuGvSuRd+/+GinOfCdfLta0uwM25/31j49bs0OMLcOQgvlCVFDyb3qC
lB81ZNpvBm2Pp8fgvB+XoBSW7hR8DD5wGRaTwpyChTSofxhxwBy5MgLBhTxOuIVxSNG7Rwt8IZH/
XmjOKa9f2agP6CIEgPD7Hedx14snVM7sEK+76xMjOw/AE9HHw2twZ7uNHaIGMzh/fUpDnxuckdBW
F2G3xwEZ/5IOakyCSGfApm0kC+TRq3Y2Niev1+/3nf6AC0owj5Mroq/x39MO8elfcs173n7e37Ih
vpT1aWJsbpVWR7z3/lZgjJKHRUhY6/QWdf9OimtMgk1W26txOFWzfZ45uMT7PilOpNbuCnnLD/J4
tn4lPObvNnD8g8Zoc2vNmBsB9l1qsL6f6qtySmQgjCMTPJ9qEM+ZUnFNRENylvf8K5FDwcqULjTb
hqEIT7ZJqpneu66UaKHufVholmGlkOtusaxdDAMVjrg3V7yO3cBMfEXFu8BCB8bQduOXRO8MYHHh
bib/EiZKIy8uyEJvv4RqiwvjNW9OEWv2lMzLO08KShHjJldss3DFUeChIcU7G4Hp0N8Ukn5FBkMm
Iu6dDHPpXwCjRj1dhJfhm3Wlib6JW2TSjlVOYQzkmzqQZkmHdqel7MS3Tn9N9vRzU+ho86jbGtCr
ItPh+/uMD+tvAgRdyWkGZK4sF4cu8hK7JnBFoz6jxAXxJx/9QzFxAdEDY/B+5nZX/UUns57GpI9r
93K5oepiMKGeaE4uAslaBjdrxO+Oqr9oc/XKR4ceddLVWB+dbfzE1zZ9lZy3xszSEMZRyEbEM2vp
8eL4dTzZ9i5QMAPSyutt7ogsBVMOH0xJ/jyM56DzECt6ZWDAPNJGtwZBLtNesPECNKAjIjGNSwj8
M3xovDZCULWtShAG0Om+aEe3WvPNZ9XmEVTC41B9vJge8HpoAnlV/vuPvoTXo65uzQIMJt/3Uzvi
fEMTHMS0bA3B4OdjNoZuDx+0I7Ce8I6vgisfobrYJCAKhW+7BQU88coZvSHZ7fmPETwblxyYGJzd
piWbISbyNLLQLQoG35JrJ5jDeIeGfp2XYyHWD1OgdqMIEIl8bC5q1MxYU5RZiaxeHtnKKQEfslQD
fXBs4LAJTiQZW3oItCTYqaTbAS72TBpDxZ98h67vCfYLh0EbJEDJMIk3W1fjUseGNmfWq1s0QKwq
+slP5ZFqBomZ6h+zUcNejY9hiFadyhXnN5t/JlFlcEOIiQbjeDcS4qU+p7iLDwMyXmcNxX9tDowi
W9daBJYmDICIX2YlI6ZhaUWRp6MMG7rjtB3ba3AgOWTWdbsB7rsawtxPxfndxCNiqs4A70N3gycc
jJ0R6Yke+xvRNmZznXKk61gbekUr+tHjzIjYJxobzKhVBmYk1qknjYvez09iCgyW3NWf5/sxiets
bP5ESo+4eUt0yddBPOhUPd1YPCAsKasbKCzJ8A8R91PUe7HZQ7SoiVfhAZilJHw+Delb2MKr10aF
mMKGW9XVgKr7jUmClSnDm4KTBhqSgsPzXJ8cRSQ/lfWL8yCB9ykm/6hvamBHSW1R98bJtESQznTP
8pZRatQ6n24ik7qIK98ujMcD5l7r849cLs3tJ85b/v+iUkFGDqnooZPm0tkNF6ery7pQ/6+eyMrC
DsPlaoe2IuuFsQDANFgrtpNSUUkiS0Ns40EQMBAyHG/J+Zh3RD9/8NSbLisFRxOdzoXZEF80E7qg
WoEWM1qzvkKZUktmRH85MEZ7KXJzC9HkFzOm6dbzwXIRel0OhHoiv9q7Gdfu/lLPfP+ytS0AjJrt
XuDTUsHVE11GVNnfILaOYGS6wbcaxDlQ7tVfaSffvrV2ELgRf3FijDHd8/b+jAALLH2gqqcH7MIO
nXFHMvqBZpUjGmMKZUr1rrLksRt/h4doHdqnbn+01YQw+6tiR9DqACp1wAkyoyBdsDEH2x/iEoBB
GGU3QWmipEXcYxQVxyGdByc8GSiTyB73jhC8qFYKcWEc/S+h5iwRDAPGKjWTa6Z7POr3B4lLDL4R
KJvYa3vpEBomlflA2VUK0UMbhnkRwFIfInxrcDXVP1Dm8Ba6AnAPp1ZKsbyLFX4DMVRJfibyK5LI
m6xtnHSXEopATbSrH5Q9Nj/JA/2BXxOwIiaAjCq166+C/6+VPMoZrSrACAUq/gKriCMXfSvxD6NJ
zcZC9F8Pvablakg0QSioR957vPFUXnMh8l625MebNBrBfM3I181kRfQFjo+5CBEkr0RkLOM3RDJB
l+UiT7b/BoK1kf20x3woJ+4vJu2+Jj9BNsDdT2thDwNsPqh1jp/goqq/03b4GnVM5ITyQwapVhCF
V8YHQULCqL3tP0jKH0/9AXMzvjsAu6qZSeFXFFjEQjSoysUNp1p/12U/v/hN23owZgs+0vc/0y26
PIHADb0SIKgRiMn3bSHiMXek0EP7AZ5N09T97wWExbtNy/RhDCfrkIk8hXilhbodK0CyJ2K18ygA
COeHiAl+9RUubtjpOOcfN1hVe0f8GdmfMmjYVN8+RguZ+GpA6AG46X9coEqZ06c5lXCV4LfI/Bx9
YtCi5nKrX6KSwlaHZkYjUqbUTThj9/RqeLPcEoVpew8a8SUbwKR/6YiePxfeqaKtPD4kJ9KHbh2n
teD8NOlR/lRsD4fKEbdhGW+udDaO43Zhpz38jn+Q1B+DPj57IRzKhWzJ/Jkvl6ROfQskDPJRaoIS
jsXOQhljrKZ30MiuBjsXNXiQlrI/L6S1Jw06K66J0FfEIFCWiyKt1/gqELmicTnXZwyRYwYtnQOl
IEODVUCJBDhoHlHibN8N6B/CfIA/DlMuXUhn7FzgMTdaS7qX82OgxPOFLy0sme4wBxuT9grNDDqx
dCmawHGws/v9DDFJEMKqhFtBI/KUkmNl/sCINihVh1FqJtLdwALPRX1SdVTtE+bcOHlDII2L23Fx
tZphqeuvgNxshtSrw7kEn1maZLQQJz0dyGYDM0vFmbPbKhlwfxHYqkhLcTIhzkdgwIEmxt8ORgxE
EJ1g1Y5EmvAPnuzbzAgZnCxlytbkeYWF4qq+54y//MxJuNyDOdNvEodCOZEwLNhoImMmu2nPkyoR
Knl1UcLaHee7WkH92oENS9iFwTbbLnnq9SWnBAcNy4rMZCc1J37ct/5h2dtV4bOOL3cCsP0OuvcF
v/fKs4aMlftch0EH5lOQL/FW15paJZNjzdieyikv9Dr2+GPDES5g9Zy30fzt+ULPgtBCcMRE1wUT
cmjPAKGqnuLeQu1qvhQunky1UlZCfS9/JcbJqujMbVCCJxt0+Rfa3i7V1EL2jg7d22B6Fqj4gULe
+MhD9S+EmY6D5GiIC5tH4Isx48iOQDLBdPMaXVk8X16JTD02vffmh83YbJj+mavHDtmg4pNKETY/
Z28mryv5AdAif6jvqrZLIDpwFCdgo64u0KV1aLqvg2+RiXDIxg5L4ZnAyyu3ULziM12/k7xGREtI
7EHff/EAE7EMVbSZqGXWdG3sbEcVemlS/3pXZm8lvukidm0L16IPQMR6GsUO5eSss8G+7KEL34So
G9oklY7SbKoUxaXyi6he3crz/Hc3k8eiT3XKbB89fyx93m/XjQxL538/x1GB+X6vZKslAKfM236w
yW5Uk97dP10fPyTabp8H+eL0jNiG9RCrR0dO9lJnDYewDGi19LG0icbWop/Tgypz3Cf79YUoglPh
cfSGEHIIjTzs4ext/mGSbDZHwUo8Ff/xyBZZt6+Gtm4QuxvG7rhJFKPqOglIVi+zgR/2+b8ccIBO
KdZchB+ai+p2SLFrJKTZRiBtix+N2yoDDHQf+mNrd/WQbKnW1SSR/OD6x/z/v/XsfO64WqmIDm1D
7vPA5kAejQUtYiezeb9z199rp0hD2lAAi6gRc5hyQB45aDZnMjMmn5tHdAk2eZpQflPNQwApRwCZ
0WU1IzOtvVWp03t6Ai+uGa+wtWxcQqmnEp2GEorPaqlKsU7dPFvfSsOlbXcPnR8Ec0lz6dub0dyg
9fzJaGeycQhuK+/T1ACDoTY/K31f/HoAJFhdCPbrW90KkzcWeeYsTE8L56AR82/4dfHTABE5W9Xj
soOj/M5XTiS0KpXMHPL4BDtjGp/oq3V4y+xzTx4Uzjxz7C/TKNTw+ZGEf40h8N3uqv4Cajwcqg6h
HL1eznHskov+gyTAlkWImAV2Xuz3e3IfYaw/DoY78Gx4krwWoJdNUKul8lqqxCEuT9Iyd3XhZeMu
CjmaWmb8llPobUViFd4rBQ/9Np1VA2NrPMpSu9O8qK8x0kwfJb1RYhmCicCHQBB/VM7dmcsmIkSG
TMAso+PJvJNR2tuk9AmqKzTdPoQYJgnMbqL491i6YEnXwAXm94THDYsfz8nPmHbW+467iSwbsvmL
2d9sjtTNMCdA/j5ty7EePT20LbdbXD5JIHAAhDiD7c078t1arL3mb8/pROlLT2uWXOucmHQXRR2B
V91+z2IY3bT5C5lXZpKHBjZ+2uVlTvS7XMNC21XcIvX6PwayNNfBAnCCSpVbMad3CamuwjHJbmSa
cL05nczOwcprchFck3gEXnp6K9ZhyMurrQTWUpCIyChxk6IC5H0A4RPSzgftaHkYlNKKmLGIavtX
K4F84xDQvLdV+rzh88YdMUihEakgOUWRmJtAeoeISDj+8Ca7C1WBpzXe8Y3Dg6IyySK2JIBZxV9L
N+RHrXTibmMRbtaswGnuX5dR7iS2CV9v8+TYL9mIawZvsZRgOiBbsOKxYcWKQMEI6u+gDje9pCsP
mxKvovT1ZMlY9xI6UQnW2Q90r/a0xQE2fNAhzZgTDqMrz58FxUAJmY8N/23ncFyoylpPKS37hXP/
cLW1fVsO4/I1A7eaa906ivIwycN9YSPORnWO2E39tqu4psRodne1k01D6CVdUBsShsKXrQbat4Av
J8SKRHnaAGoPKc1W9rMz8PJovl4gcA8Bq8V0xsb8HN07NQrXzTOPnuSgOYxp8r+Wfh/0RVpgD04p
CzluujltPnb8CNM90VNT9tO1FgxWkeMTWON4xWBgocGMIQfgp2uwc14iiEfdramByYyiJPbMfjTL
kxHLz4XgYpcspZRRbPNWsW5rsg+NV0/NHW+30HhG7DPOHfOccDakCbYxhh6sIM5EosvpmJD8lNJH
76SgXRGz0idTvUDxZFrKeBMdt0a1vxzHQyFfREsntNor04Ue/rcBnShffugT7vXoF0+p6EQr3lQW
439XXg9+EEQNQNi0LgK0JzmwYFJQwRQPZUAUSPKDIiFH7eaBZoI+eP07AvDsWxCVS7Pwr80/wWyZ
IKwTcr+TxgB70gkAduZk7CIFdYBQrZCyB8A1MyTPsmerTqdl0UXv+/pAZAIjye8FovfQV09T3nR7
8vpwUjqpRoL97DaKgSmpLGZxjl4E5Lb/Z7vHUpVzOTeNcqtHICAfD8HzVse26nCDkU+VpwMfTPlv
S6eIDqo1E8W+s1pZHgAPi+jvs6jm5u5/9EMx0md43Jma5YH7NwB7fmYFPPR4e79I62btzGHUgVtt
rpHqMf8jQWtrUwOpvM93fPMmS+kRIw2cZjvBCO/wEm+HeM4in8njqNgOdZW/033duagu4XmkmnRi
AmUwd6y7N5qrqFA/73Z/0T77w5YuliSFKNpUqybAxC3lpu68UD5tzhf6RNYMyxRJFHz92rJP7KCJ
7eTtccm6VS/d5DaDPqK18f0JA+87/8Ijf68/REhojwhMYCib3f6BmqFTWBHO+gNkmoIn7UopkYYl
h+e82ok/JyO52sdbghZTy+nOUSusd4N6MoicAfE70tayTdJqXTWp4Ajt7ghVPlFvqg+q+mqdE2xJ
TRKTY3uzmucLOlD/9WBh62ZbT5dPXLbntL1EID5/s6uPQvrk2mflbxo3J9jsg6VXc/Ozs4A8cc4+
56X6ME3cj36rIiBwqfK1dY+jo6oeDRUfdM43bs6Ev3rwlbonjMohPCWMblBBQBnwMDbxFqvLcCYQ
28lC96Tcvlnjfp2Oo5fqXgHWHAXfjNnF4Q3VPqpBpNqiedUbiROcrKSrVQJ8xgrNM2hLaX69DPr1
SyC+BRBvwxNjfWQgXOVlyeMphRbwFG1n7KJ0Mu+3lpxL5A9iNgwzeF5nULmxVM5pyL+JZYplbq5d
+ezhUNYjV1krA7APO3XhKedS5GzwDcEfk/2bBP1v/8MO5YQs+NJ0eGFadGRuCKhDYe98CcuCdM2o
uWSuU/tkZucS9SgXf+7ZVKtTSB7zp2a46bZJjR0+9SSHW9t3F0XuP3RbAKRF9pPFAAGX/rrQB5lp
oBzKqoBobOqHEZx4cxyc+miamkeUdzOjrwQcN0cSDjAAmAro7Nb0A/Vw9UFYGk363NOs4L0BH3rI
qMbMw1anUSUsTs/C+h5J1abWw97NrmmSHvrgPWAI01AVyAlnT/sp2KnTUyJ36Ix0txumye4H+3IF
POI/HSxmD1Dbrpz1kuXc0+0jc/t6iJ6DQ9YnipaxWFucgS49LjdTJA8wEr/5AaoGZehcgma49pwT
46VL3F2xt4PMweiEAXt7IJIGg/7jFmsNrp2QHYf89FZfZsh3SXNla+L+GS6j14nl+N9nuy3I82PI
Mn0Zgqfw5GnAs17tntKi5pXAQJN0Fm0YYb6DimlGld0Xp6CnjRuYoMJGePW8oqYsIkFC9okNLaoY
QKMs9JOvyUpvcmtlb1EpUuzjzBTQYCZAnfySZqbPwHK77kNcgBZgRlarSbjWvZ+pifeQpzVyNol3
CbCu/s7hKeB/q93lXja7p2q3tDt2acAj4y8yza689Ko/ZAxpQZSVFsHllzPjDNyuPo+0V9x3wWrL
J9rZxZIItvP9QEGY/J8RSN7njeoPrwNaOY1M2wN2d4PaCOv+IPH+iiWRx2lccwOih+ex4vkhKNEK
+zDFkL1DCumTFet5JaRjK415k9mv9NBLBaQakZL/oXR8BPSoZf52M4X57y11wbTxWG+1/tZhkpph
PQzKQm/lxsgwLCtweusVIPZFyo8K9ep1mMKFTheZ8SB/lugTPkqSixTSU++r+v/4rsQaPH9bH0Jw
sffE3/xThLPOVkLBvWwQoArZuAzYHPqKCVKcz4Ih5IG9DeF13YOM2DD4XZSdahbIHwUQfYhTeirx
ZPnApnDAHuktzRtwDQ+x/944RwVEJpGhmnAtno+S3uNUi7fm5oObhoK6A/pEIlgrsJ1JUJR1OrDq
gxC6YBjhb/hHQyiJL8KoMBivciIlAu4cFxZwWbM4TVUR7wGDb2XAddd/fhOvNfRa8B+v38IpVwPC
b53LwfFZkANO4Jvtn3/M5skWS8t5GGyeRcrS8OxldMQEkZMBEv2nuyP6nID5He8youQVrQ6gTbLB
wmYSjDAy/5fe3UkLF+pqIBmOA0vONG5FeCPnLu4TUFuAszW14oNDgiq6qDavB9yaoucOcZFIdXNe
3xjflrqmfWKt2B1UEbXy23bdxw5dw23h2eKrfffQMGXylDVVQwBxkqGCDasn9Vl3KpyD7mXvve9Z
3jc5lC9OMux+mJ1IOF1iQA2egdqSbz285dxMNIk0YrmMS9e6GKAkId4cquSTY8EVqVMWfk0PXBoe
Nkyz5oXtG33MlwQPLxNmsWWFpRX4asgpxpiFgWk2dU3/7OMfZeSbAa4ludMw0sKw8M1vraDNP0hA
X0BWXMZesVRbcmLLGy2EbwLRMQO0PsZvHZyWd/Kyr4Nz+CcDb5MdTdsbiclvKwNqRkD4OvAISrEb
1ApxBaX27HL78HeBAeDCS9PIue5Tz9PLMfy+2B9ebPkYV0jClv5314xoeXoMaF+gjLKNn3i0ickq
DXc3kXQy1T3ZECtnPw+LB7WLUXWL7qc4LpmGcNIkmsnGgHlDS/qErnaOOU8BlZjthTH4SkCwDm98
ykSN2TcaUXrJmY2ckUSvUkw+7jQF4SjB7pnE0Ou94Y+0de8+MDsyOx0cHO8oREyCVaWG0VcS2oHx
lvY2xiq4WfEfIDUxfHlD2xr8K0YCrkjgRfFaIeji5CUtmcd4G8foeEPxFqLZWtTLfqnUFX8IiE0u
w5zpSAbMGvUkVhr4rw+xquGpavCj6RnRNOiFWwDzZD7UD4K9XoeU9RY22yPJnVpbNiN9GSKFLAPd
+3o5kQG6g5chr3cNo4xreOiTZU2MQg5NtskFYWsf5IvUkDCkRdWjZGVJlDkb8fmjfma/HvLiNKwM
DFViM+foAASHk8Qo6HZ0xCEDSlem6P7iK+vUAU5pGlvtQ203g816X+f63fYDXJOozhiuopJNUHky
ZydQLvxp/bb33Tl1Bh5R8CLq7IjEn6kkY6fbe2tGwYHj4R1WHX/Ok/pNgfdbwSNF4ea4FWRrdVP0
fBE9Rhq7JDDC8ufJz4aa+C87xOoCvEYpv6ZRiKlHM4MtkuUriDhUatY+3iPNvct8VqJftz3kBXw3
iy2OFM0lvzDMxjlzWEfIeTQoYnUDKHGE+hugrJtqTWykC1SPi6E/+1IW2oRijvHD+LnuRHNvcUfV
84QacEJe8VMEk9v8nBv9IgT+cu5NgFuFxdK4PjGw4/MxIFxulwQc6/5rJEHYhwF7u0LHQDFa01RW
rJWwpH4BYQzc1B8/WbDdM/tLEhYCPCHIpFr5fYmkJSspeazxakDL7pu2BEm45mqXB3dwxn1mfk4s
p/NGkpT3I1jnq6gN2LHeVZ/JQiiTWi+6D3TquQGabyl/U1QHMxKmGoGf+M3zMUpMUiPeZyVDI0U7
nJrVOzUNVr9FNhY0LMmimT3ibYuBR32yk1eUG4rhrSSG1oEJf51j7amrQhb1fV55GmXd6/2hn3ZW
JeaLz1FOuoBXN/SwsavB2wxZHynPRe+8ME8+UnaFwtQ0q1Ej2bfhkwQSqqmMMOa63zbvOqUG5P+W
9OejIujOekodZ9JEzdi0iYOmb/lWwrmZKbLx9bEULV2c/M1hxJUCeywr158wdiHcswaplg/+5c5Y
wA0KphNNtQNxIy6Xq31pjGSTnIdMJ3KNQQ8HBo4uRLxPZVcJCI5GsHqLzsDMh7Xx17NW+nX0PaS4
CmskRUrjH3aLFzZhjCJkcA1NGbkKKL5AbqV0oUUGHmt9YO5anCmvA3XvWrSqezjd6crbf/0xkKN9
Bb+4fRN1bNhZQws3Fe9Dw2nqyh8HCNmKKEXdbEWKXkMsKaLUXw11KhR4wjAD1aNmjYtNgXb7KmDl
EG+C/DagNmjjzjqKGXQKi1F8YuBnpPNLSQPmjaj++wW+39u/X12/PXnB3adDj10UuG8wrbz7DNCQ
JTRSMuGenzGpXnPFVGbraRYC375QSbVQUrt7F9HiuuS5Rwgu5DQqY4TYgtZvkMs9/PTJ2DnjKEG4
b41WnLg3d5LW4/Ug+T6b6V8HCITUb0P/C1Pd61Enaft0YHUu9r+MDmw6jV1MbV4J9cc3YwP0mA+r
xpe3/iEAItgWgfbbchzfgzmWvzYcpANNL4JHeerUBNF1qpcs19lzYVqAie9Y8lnXePvaJCqZSXyV
9QryTUwH0LTxLjOguM8hKpzxFG2PdsTBLbX3iMWJ50Wy1jVeFKlyb+AxFyxyCNcvbuhBH9yqVqy6
t0rOzuOfCuRqQCaw7JjAq8ySdQpfUojx2bK4XORqxDeUjLABz8kCTWR0nTn3lLD/gdO4tjZMgEn3
w0EQud+fwpBVjbHy4+gbkF2769Lrp5IOrwvmj+9K+rFTZHX0FWC8+LWeeBLkc2e5obgkxSURIDE9
daGeI+hnIViyH9tUTD7XW9yoQVH2GblLkmrhMVCgTMaBMCxMkNc9Ftzbqd+nw21cmbc3Sv01HeMd
GIK+bAZuWT4nNWVEond1Nc1gVBYfAE/GSchLnNHFdQDZdlj9CZvUzN3idKZ6uJOBhwpgGb/VCYy+
QiTpqBzBGpCdbPiAQjRLftxjlhFYGL9tLIwohoFAwVsRLhDP9PFL75kD2RJWi0jfn1gxSu3ZD+Jo
aBOHghaJDZ9BlqBHeWxU29NGgJSFXZ6uWeJSiwBYbRy8SQpuheKyS/713/szpwHhxspbP/oPqPVD
kO8YvLyIBz3IOaKMZxQxVeCXW4bbQnTtUCnfq1U3KewW6Uo7W09c86vL7P4dUROaF3E7R5uDhd6Q
cFZpt3N06DC3zSSVhnap0ozL54tr+qc29PJh+MXwmeZv+ui5u/xe/sCoRefQv57VIFY1/jDZlZSB
e7CEAV3UV1eSulN+voXeO42dfI1igU7YmRwHSxwLIYh61H7k5TifsQcYTIyfYlKuwqs6sxqhsow3
NzUGcctP/lfx4m8pljG8RvZcW6JnvsKrywfxIQ66ZcbU3DjghziZZeA/8K4Koc3pS9x31da28guE
T2jtUBOR0eyNz4HXj+LvmyZ1CnybxsX1MNF3Izif4jYJH8zoypuEVIt1edEgEzCv3qaAZtJ/eMbK
VNs2uAdNrsNVG8hqg8SIowQ3zbi8UMMtLlgumOZdqceuzxET2ZZzg16QrxttZYwdmfMcqnd3fFc1
eVPd0cvUwY+6ngLCfeDtCqyIrcj51xGLfE98/e3eGejdpoGe03/3R0xrsuzFxzaYkdQusRPHCX9/
metxGHPLjuSaPirKbtBuowHZCL5aPffPLdsDjh4fWaT4jXXZe5QJAPWJf8KKQvFKTplKgdlEdN2y
sNMaDGFPXkM5pnm+mAE/WDE+TN0DRxmqy2azxfTUy53Uws2MJKZuwsGYY2Cmr/yx59Cev9fhE+B5
oNF5HNE2TPgL1InKxZDnwvwemnpFAnolUmbj+PZ3gGc4qV71176ggkSgYMA70zqfGxla9aEgyVSj
cS6VLsZoBNozvBNyK6LKOCwjVeC0PW222XDtElYIRtkHr4eGqspDrSbIA11mPHpstiIA3D5iJB5g
d5BuhHILRTJSOVtLOeH9cDt/+OgUTTcXrfBjYCHDYrwta5DewRGmV2/RVUi6Aa4hUNIzoP4vygkG
tahMpLdarUeohRCNl5c3Sa7EcefRme5+wKf3If4qcNsMuYS8qoJkqQ4y3AHRomfozKB/qE56+J32
LvrjI0JQHDgN8sgaCy8YsXaoQGdvq3FNUH/fwhk0j+gAUaov6/240taDoe6Am7qSjsfgiAbBBAHI
LKcioG/wyfQujRexISPg5jKB1xowS3xLEKBij64hSWzz978dzMK4yLwbJCdIQI63Skedbu2ogj5D
if/3vUsd/yCCkKfGRaCM61tH7ggZ0mrKGhVi1gvwPdNgZ3Xu6ne0LCppmx/PYhuYta887p4hsViM
2Tydn88s5eofAsV2g3OVSciEUB2vUH7pj+pX/BPdc24lUX6H+OZPmGW13BMhflzYcrurNCyvgTzN
0CdnrrMxBEpDlkKOvlRbzqYnOTWf123gdV5mR/qYPUsrUpCwBtC2eOl5H9dxQElm4QHNjKGB+Tnc
G4GqufvjZsXQYf6tsg2x8h1vUANtQbnn/oA8lHh8i07LByCuW97ZUYZ5wdEXwT8o0Vcsb1rd6paA
ujgd6bT13KIJQ2TXVFBwbh2Dj0ceIlFiqOUJCKLoFQSkmlDh7mmKM46PdKtavHpq0E1IIL/MFrtc
mbnpLtRgK9Bz0QxwO85CNIQf16jMi8IiXtgMIl0NqW+2V/Jn4SXaddYInBxjjKAM1O2F5wvHYBef
+mPJLqmDKscUizuY6j3C1aytGmFOddiIosAkaue9gIwYxljAgb5HVBf+bgF9M9JDdh/I+k2vcphz
98ZuYXGZq2TjKEmiJ9rGGqT2PIsxfH1mjvRhSZeMwBqrLKoYw5ByMraVZ7lbhaCt5A2EzisFUnVb
gtUooEwx7jF9aEZK3Y0862Q8VSKQNcFzh/YrHlwwo1FbosYIpbdDUtSC+neyTDmi0qyF4mCA4DsW
7k4MBU9W7Lp4whgSL+aavxl1x4PX6STD+rn5x4jGp6UuOH/4vDBhaiHZwhjVW/SHQa/ZYW9QqAct
ndE1lTA/NGogCrsBuirBXrBxnaAdhqyDCEON46mdHn7HmJDjtQ0VZsNZSYD7tpMk13+2yOTsW9KN
Q53e5uug3eaR9kzvdc2HOVzMAY1eAeRmBetWhXVHk+GGVicVMwUhzNKyd9fhXSBgGCGzJFhDJkx9
yaZxmVog7MpElqjlM8iXPhzr/COncC4GdWjP5+kIjGH1ZpghfZ++toBNrpzNyx4drQHgNkVN5DpW
Wlcy7omGmpDj0IttY8DoMRPj6Dg/d0jvIsm7oPGlHDxgJF+/t8YPWH8BlXbyyp8DqMq+QvwkUI/x
p0wq7+HJq0k7wMXXWBVNnvcyoQOZryKFo8BS1FDN0DUADw6KD4Qn/PRD5g4Z3yd5Eg38z+mBknhq
pVt8xgGH9snP7jqctkJYdIfhudTOJJggIB2yqEKsGA4JA9OUopt7L+KIcRlecTrXbe83XSpyd6Bz
gMDB+umoFYLdEuTIvsnOp6RQLWX6J/coux1XFdtbVi8mvJ9cpPCgOE0MYKU1PwEK7F4H6KIbyj1k
xB3YaMMLeo+pcsakFkq+DeuGZsRolXnd+YdnbfRC7aHLdeBFsrIr/Pqgg++1pmIsU/13yZ0gNQxU
dgrb2QYrgRo2yAZ8kg4FTLrp3nbk4G7D/RT9d9DefYfy/CMhj7QfRbSJxTjCM0K64fh8lILgtd/+
P6oCNOm0Rry/lGdHQ0lzYVIVpfB3ir9lPPuAooUx22Du7iOExC+Gt/k1Z8LhMrk8OCe/6M9FtvjU
pfNxvZ9E22WSBpxQ2XrsU7bpspSNsJr0UJyscDbDrmi6DXCU8cYM5CEz56a1XaIAvhPRxSIJE3XQ
h+6k/PZqYrR4oHKfHNCkrHsn7iGKzm/hnfUr4SGPx+/+lMHWSrvDvPZVAPLXhcJdclMPzFGoHFQG
vQ332gWPSqwA5BJdp4EGRIOf7gWN2L1Ob9cEhUyTwbsDZ0xjW+pX+CsLHC+xadk0CR5btmbM1R9a
QFQrDSnDf2sBiwh8A/Nib7BkDLUJwmVyguX7Ok2NQiB5834IS1VrtR6czYydB1ZWzI8XAufE1+Fq
lvpT5JYo33TpR/9Y//8aa7qa1lA3X1mRqdMGUansIe5TEgFiBanMtFmGBWMUr0jtEFd8gInrZpaL
xNLwPgFn0aNeU1NVp7S8gjHjJXlZR/iaX7f1g/vC6K/YaolodmEsEU0UVS+vixOHnpy/dT9FVdwK
pRE2ZrsBmC4CZJvwb5U5IzNYn92X+P41oE/fXfE4kW7ZEGgme7ZdShZg9Gfk3vTnSrCu7X031HIg
mPbxv3utPLqIOxaTGOWehltlY4NsVfTBNvB2KN/cBf6Oo/z/Yr73j7jJcz64SYdAv182Kc7FH8ag
P78eHYnC1l+oUBzMWVY1qOVPXORCyWHftmfPKEmVr90KYGdPhn02vdGBjDOZ4CO0g37mPCF74Vdm
YHQ+9MUgkbGDrNsJnpVM2u0/b1C2VF0am6zNDZDTp0xUXhDBBPZr5Q8IppUmNVqW4R3jqTy7p0h/
LO8FtxvV+B8q49AeNzujE8TtchxtLC7M7VOqAxm2LvulFzzvQczhJA7YrqBaK4tF/zIlYBvecLPv
R6qI1yZWLRIRtNNfoHV8R9Fmyh8McATvsQ1d2ZU8e7Ej0Z0OEgx8ACwPFu2T0/jNR9jlskEt6u0B
H6n4ZyiNWGUMWgyo7JiTHk1ykOcRLv24pUKBu5TctpEjHGaCg8K5eYkVJAzmWcRI6rGkNwRN+51D
tcTKExedyhMXxEUuU6hb+l96xuwTW8eeOmkiIAViSrKEaHBLqqz0a/GzRd7Dg2076/diZEFgUAiS
kgxLHdnyfWgxkL6zoU03E1wFCk22el/AVsCj1jBo6jbMGgtdcvgGEboSCFYnMoO/rM9bWi/E10b2
A7Ml8BbDAAY2LlnIOdEbbWq0IK0a3JHhsK6d24z5uQOVCA+W0nWeuIO0QEZzv77IhryIaIQf9c8P
4KqMkGtY/NT9Y209+ewviA2/EBXEs8zpAMM3PhTut+30Raok2DvyxH527JIDkBs6Q5nnvLUuRiiS
naLoLsQDktXhSJi4ZoqbRr2fdkUBGS7aQBKwi/p+KnwQKQhEjXOZ41ja67+cmlbfOfbhO9vlVcNF
c0mshdFDLLgIc92A7XfyGoPZJYOXjqy+xAbmEFr26BJMCszCcoFvIjRU8mwZ8jNC+17hEBdzYZZA
1EbkhS2DAAVnO54Df19MrR/aBOPxIjhAk/nYMoX2FqVjt7fNwcUTwRYVDhbmMlf9Lh6FLojqYoOG
mRqbDsEUEeZhmZvk3viLUPQryzPoqfzuz+FzrbyzqvaZ//DPWlt8UqzXCa3BjTG4+H3Un/c7Wu8K
3GZeevhua0I40+CoArAJfZFu57pOirfMCx06Kxtbc+CBv+pYetfMIcwRNVnjjvwTdgpzQ31FAH22
Oheaza4b0dKOlpBw5r74byhsIBt6eJ4w9E8TReUKNv862Q33JXt66dz+d3QgwE9J7Ls+RMGUkBsH
WmCoDtcx7RLQStHWAR+yU2toueoX+hJMeeWfTZB5qkaGGj4XS1AsoDASoehtBTYFTaHnIu8p6QcL
DVnFXcx8QNbb6JtghmDT0foteu1OsV581NSEIqiDXeH+U5HiMBsrl2poPsnYFVdedvsvEETtgCtw
7Vp0HLrWBfcr3XVYmw9SbhGBciJv7UPC4GqFkTQjZuYhGP2+a9/rTmXUP4rIMHT7A56HvZP3iSOs
cPzROP6iL9UGuHfphnG0/ZN3uGXDpDHYxzzqBhko+o/85zhpj8KvtTPfi/jsQD/ailNVZYBcjXXj
A9GBvZSX1uuB4HiJqBU+FlJ4fdFPjmsyWJz+VAEG3/b+tzIv6lzoB/eZ2v89EhC+SMKZPpZ29g1J
Qwe8lYaQG6WbK64AudOy0sZtNOCb0gQ7KYbS3p8RkLJ0iBUdIw9ja5wMcLu1A8rpYHYbFoZb+tfS
wpF4YxNoqKeTAXzxhfoMruXUa+hUkyeILdU2w4rxXh3ox/N20oAEODXzEx/+NdRJAhPEmVQBknSk
YliDK2Hm4fjWufGoSLdYYcbqLxq06bNNyfIrtEcID353rUaEtURH9tBDgEoNPtPhg4fRfvcd9NJ9
XGE73iAql0HarFyUiWkWlovKzaTONeB3Eh/NLE1XckYA6fg46bDcm11TOP/EIVy5z5ko2FUg1Grt
vwHMkxjDZaBapZcY1xTFKkuo5iYIHeQtSeodq/GrAljuRV2mfHnfTaX0gOpSq6Nvk6x1J9VraXoi
x5NnRHOt9+q0rdon+O6NAL2V9bKEtt+0akj7P5DYThfTB4QphksOR7gg3LRU94ap1JbKLr6TZj+Z
kRMrct5oB81BUIotyGVZCDxWRJ3NetfEwuXK0ccu8yxx7hrsxtiBfk0GEp0IJEWV580WSfBJ5Mhy
zd/K6FJDvubyqbam5pSuK/XcAhCmn3zMldwpEn5K6mxhfCLo8dj6kvP6mmk9Ay0PqNAprSebD3pA
HNWYSGZxa2GP83cFFRaZThcEMxFMSdHRrin3pNaMXx9aabN50wru1OF2Zti/04flCAvT1Z0GLDLS
Crqu85xHQG8SBSMWoFA1qAHUNXNLrZRx4zbnpG38RvD3rIMynGUb74XEZXUP5+GINAxG3FYgNaT2
/ZkTR8zHyWy0ZhIh1kOFpnXGD44Mo+NvNNWYceqSiQkjcQ5NMpxVDfwNTx4kN4IvJPSP3+Q3CldU
CbA3GGHTLj9MQgzoqIhOaaAEnoNor6WrmuFDnlz/YmCA28qVovYek9OZF6JKbb764HifeVuCK0q5
5EWUB2/Dbj44hHmi+nW9DoWVrmTgUFdkOsj4h3V5n1DFAWe+l1vuwpdAwdxn6yeY6oq/0rB+goDR
jMK6IFli6my4Fw+cpFRHcJ8splnTSFiqMgWvsRC/NlJ8sz9MRJQv/ljD0vR+2m/hbb/e77AaxSLN
UpGV+q9cmrgV4QmaYQ9qPQJr/GQNKxzTQn6hRDH+RmD5MHYkjPMNGn95bDxoJSL+sZw3MQbQSzWn
qffhNDGzrTWFydP/YUO8Se92+doiR9QJbNSwbsDvjYd9Bek2I+nqJ2x2kT8eXM+mID2HJev0bfq7
Nuul4i/PIhIzovL+2WMnUqbZzn/J808fKNxqrAR1Sc8ScThEzm6Py32nsBCsrKwhb1d2j/CdD7Al
/8Dp5v3esY2jrN+wFCqeVRnNXF9pXSqX01c0H0bra9mFPUI+IQas7lJ3ltcK9I7rMjtUKplGW/Ju
wyVaijfBaa7gcTAO4w3F7TSnpfl12Kgsx8wZRY0V2aka6ra71kzhoL/z6gCsuBxX55nIZzgHIx/M
USeQHcOzfK3AGv93jOxrzirqH4Qk3H2sXOc9spfrDNN2p4UIZQUU/XKR6ElFhDHwHF/c4tMgbCpJ
DIne7+T8D9cntOJyRqjkpALQMTU3tiPdHPapofbOvzTc0xTmJfOag3WXTzhqGIPqDuyng3Ai8Xvz
RyBIdZS2e8t+X2ykKhORN4qRrL5odJhyBVrNNZBYvPKFJ+v4QxSfj7iSESbSwqsP/aoXP2eQqXzh
FolR01bZNuPLv7qkrPl9J1Va4Ku5NDU0IUIxQdNCCbMXcM1l3fg1EZ+njOV+OvsgV+4vREbRqthQ
/LiyTyEsOnS0sMvQ0cMS+Vgj7fl9L6Z17HQ/ULUxAw5AvyxU52X7tJmAXUeqhEVmDcc1p8lCciLl
Wc0M/kxHp6OuvtQziTtc9q4MANBJh62LYw5f52Y0JRt96jr4HZVxVVN3Rd6YXB/K7D+2JwaU+31m
Snc9eUcCN+J+HHS/Ufz+kXJdwOJ61vq5xyIjYFJMEMcJqMwN2maAQ+xgJhNjangMjxYtm1q9im/8
bUmjRgVC66q0nydg17+yZE46z6UNhcL1zlDXoM98NOp9gQG17OJI32wzSPC5xxI4+nwOMJooDcWh
2HFYksv0zgdnykpUZMUkXKs92js1envR3/OdCsyvwgkQgfncrBhZYTds3i9Wz2cxb/TPrg3TOrQi
9cCcysBOfa/agWcg+j6UV/mXgw5ZnOhiPAyjHg5jQkX3R9/P6h4E4WqonqxxtAncmZn21g59Odjj
+1KdA3uG+Ia9m9JDmwd4HKoDIiVVy5cLpTzT7BFp4W6KYVUxlLuUl4A3aovpkU74U57Jij2+RwSe
Op/otUu/NujV0WSbHQLkxavXzyQ3XTtJCy+OJdbTsRFU2c859HrpajP3l87TcAqSoU4sCz1F5FC6
wq3wnuC7jTPAldxBzldlMg6UNzHreCwbUpleFXXRJQ6B1+hZWoEWOJZiDFqUwV3f/gV1UH6EWStr
OCbQexbj9W7F7+sY21quNHWjlRlD2jewGmr0HH4QGOmARjOW6LsMmax2N+E7g37DmU+DtARWDwHl
uJ8k9bVVqW8UN811/0sBRaRENaNBqvhwxxVTCF1dLxDdj9EYcLYcfRCIIhuZmv3bz3A0YRVozw3m
UdbjF1gK4RnIyq6el5SMpnmFrWNIl6WMW+lKKLBcoQJLCc6YsxouMjwimFRMap9TAUNPPySwBVd9
4biWE6e6FU5D5e4BxFmsFrlnzfRmHqqMq2l4NK9pkoYVsFb37Z4GwpcCTUyRQySxdI6tB0gqdqw+
VRL7LaYNjovGNQlY8wkBube4Jck6hCeRc7gUpTN/InHvOdLoeAd4OoYr3rGeRmIADuyhxaMexvzo
1BEMtdhTMs7Pc4yFOe2Gft2ytF2Os9M0buh9uRtz3fM7ZG2hFg9yy6JJM6qlrEwfuJ85h+5rW6T8
tqBZkWkbtVwWaM43fL7vb6HvY8aRtbiBLvtZItnv9R0K13LAjdmrZCjkceSRbzcF7zUI9CAXQBJO
ySc1DprZscDeSGG0/SOgfKRTOo8/ah4iI0F/+5VBc7jt2FQCsXwpvNJF8ve5fNXD6FbcxGhsLHn7
FNpop6dLU7727tM6G2haApcK5flX7PPcKTGe3v34HkHGHy+Rhoq3dINpDV6Szrzuxg16Jq/y+NZM
4FyUNjsf7v8HzT/dfewjD+0B8Hu+voGrTorDxTAeZaOAsgjlPG2qtdIZyS9PkonAXI3eXBiepT2x
UuKx9HEhGj6SfN/1ydei6+LuEH5iRJcQLLCNNcrGVEV7dInNhoncdsqMxZIV1V1yiPb7WvTv+xb6
NwCU1TJSZ1kkMAfuWTz++M9grY2UQKbzqwmB2+yzL3BcLWUqAUO6F9nfivPLHgVROJls2BC0PX0b
kuUZL1guAEQiCAIr72Lj/drGc2ng0UBBBijv6XQWDyG7vx3EEVrFXNvPbtc4QR44rIqxqLHcjw7x
mhM5hlgNAPFFSkOvvIgeEuGAFtyJrqK9iO6zCrEkozbdRvRfZ8ehtlkjZip7WqLWBOnUaixa9rAb
Dc9jkhM6XCzaHXqcTV31j4N1gcRlycB9RQnDDPMlJFdY8VRXid7TmrXrpS5+BDyIGb63uR8swr0k
tJOd705nz21YnJYxJOu4HCpBTUay+0jom55tUEmSWYquoOT/tkXnbK5zD/UrTpjKznp0idyl8FW5
7kb4hByLV0hKjGzz5AuaC5iEuI3vXRzYU2x4xCHuLBAaCpBD+VvyEvEZd40/TPZ+RBu0FC1OFsqs
ic0x82tQjqfK1G1gDT4TQd0d5r33NasMGDhjTrLuO0MoJwQa9RLInhnfzw+CzooDMF+cvc0C9lDi
fnYxVeS+M/RqJ2bsEXLdcYuwpgaXIeREn3BANVwvj205nWlNZ7LFrDmZkncRooaPL+wqlamnkKOD
1mYZaAAKn0tb5oglDI6zGPkWN0CGFrjzRvp8sjBcEMLXMVr9GBN+e86Gbzi9Het7NIaBSc5R38K5
xyOZvh6hp5Hh/KmlmsU+OGTCXRskhgi5sG3GVTVlkMBd777RkWd0vAD+frN+W0LeXUHBklI6BTGh
4s+bAxf2mYrT2z7vnsCbli0uN9mDlbpD/QRc4Gj7DiMeMfO87fwSi0y5s+CzJjy76t8EhCzbE69J
T5sqAzf2iYUY/mPfSFCoGsS6OEGKTn4P/s1tzpWjkDeKbSNR5nWW33idDtTfefYdWR1any4PnWjl
JBSJUtj6FbVV0k8+bZsCXPWoj3VK3XS0QuRtb6zuzug9spzSxrC+WaLyvTRvuSC8d0jW6PQIcEOo
m7hTsVFq/lH6oywEmsYBXj+d7iRjHqVd32+87wW60PwXwbUxOFePwPEB+oSBUuOpSz6NXMXuXb/0
qJ+oJxHH43H6JBhzp57RL9R09erSW81/qndReJYufYCMm5EbcDymxZ+cmpTxHT3wnvHFrXa9Fr8X
jmqTJ2msXK1oQNFPYF55mcGPFkMLeroew0awvQAXKVHRwOwqMKl05+r9qh0mRKF7LX3juOl/l8bE
/xOhP2cGmRHAo9RJjrkQlHSBATGjqEFFpTuummkCknsVAKXHnDBO7MQUkn0FTpWwtTWeI0CGhGdR
1y9q7nbibXbakHpXWkDR6KmGXUOtJ3+E2ZlnRTMueW+JR+Uu9P6w92ekWs046YHxwEWV90HbJsSz
ZatvPIOeMq4MZjw9h1aGrD0JA+j/icok9ar8y95BMvSzE05O5e3ZVdeL2vF3Cl79Qx8hmusZJl37
Bi5RGBp4rncxDUazlpCjXAPPeQbR7Sda1f48TjNKw2gWGdh9b2TlmB36ojvMI4P0lKl+VXGyeqC5
dNvrqHS1AE+IpefRL97BdeC5idUmsJbhnwlPK+QiJz1zSqohPE/AzWCB8vmj+yaXjeg8jefnSqdS
gUzwmQwzhYLvAdkW0UsQG9eroqRR9sK9LiBHrld9cBseXyScpU1TH+QPY/2MmNkIYm6V07ELhNxt
PwpRddeVqcIsdqobACbMkZpLsAIRpA3Jur4sPfiwzbByLQ5aqcm/X1XxzCnYi5CnRhIFaB0y3uYG
c9Kr0Z6lQnjYNNhy1MIQYwBfR2RAna7Bz4S/AB1wd7Gj5wbA2Yd75ER2CKBYblQxWNIJzS2oK2tw
CjdZ2FKdi5lG0fQYZyWlSdRT7XLL3vqEEGwf1mgkQnIpPMOmpDKjgIwQiAPfAUM1k0DBbFCiuaaQ
KU02SRFM91ZQGNSj12HCq3KC29fB2cNDZ6qHQTLbl/Xivc/QWgjuA1B+awYwF3ivNXBMay8Phfn5
HwokJuwPhh8tf444TvKjbhVm+S60D6BMd933HU7NCX2RhnwwJ4WlSLXo91lvGkqq39E5zP/wuSA2
kQC+7HFhhwWnc/OgkAiwr54/vXYqdJ2d5WtFHIfj/oOlaNHg/MMZcS/ELsnWDJjG1VJOuVksisQU
TCmkxxVlINP3B3kmQNpkO2eoV659wUWZnXwfuVGHjKcO+hDEs5DVnfd81h6I0ePcRedvHs6Ya3d6
bcl3kLzBmtEwhQfThYSx53JNWR3R1pAJpgBzOepgQ2HsfUsqdfNtusF7G+xcw89fgXw/DvJKRk4G
tE30grw2U7Smser81fvD/XOHTD80FVCG+2v3qkPVOwGMk/4YG5ooSKuJtjNlTivhqGdWQaBvTYV9
heXS9o6LcHzvczLbUg4qyDlOY5+QaQIyugCjFuWl0ZXLgoTSqAkWG/+Eo2CY7FzTzuNFmq/06f+R
wTCyrpzT5o3oOQguh8EdL5QZNYGb0WtgKxl5JCKU1dZUJN2448/6ANTEmdRXYKEFSiAvXC4pB7pe
DbFj7VEo2h4IcnN+MWSMbpfZdNcZnrzjdTUney/4QdsLoHySH/pRhpX4mkZ+Q83aX9rgr4HD8/BM
uEdWOo80n7KEX2tu+xHZC4xNsPX2BudAUzqHGXa4ChaGZSAA+oWHI1oRSw2FPG5pWBYpS0CWqgvE
fl3KXw8vEIwBYG2VlM17N3yhZicx9N9XDgsFyi4vI4PxwwGct3riO51Y8TP6MFasolYCvI6K0Y+t
/jF9p8AX2Q3sJJisWjDWLCkfr+Q1sByRRjseABQXNpeTV6ds3OWuBhXJb8WyHoj40uCT4sD5aVMl
I3EBjYBxT4QaeKRP6AkFJWYkkieQ3+PTdZVwzsJMu69Cmg18Ok75qn1Y58MedEUIHFW1rjOyB0yf
sJXOd3SGJ9WBqK/HHqvA6IcbHS9kdnkGJyDrgDO1X8TgEDJikjA6jVwuSSn4MkH8ZG/6kiDrN3bu
RDH45pEx+Wd/iWXk4Le+rgobHBNjgB3HDVaPVAUSKr/IZU32k1+5hB2ON+1CCMAx3g5zhEYR655b
F6637QevGTQoQM8fyBb6kdEQGJKu9zNyA9/hwUuQVIG/IPVDKVEV4LxLXKOZ0KmKyo2y4vWo+3b+
zgBbBvTAMBaqt/9ueg+Ic6TOyGfiPM9lHdbY+FhteZI2YbhltjcceNULsuSiNCjOhqwCc/9z3bJu
JRbXuTOs5LsRfDLeyVZGGdRHhdT+vRiPJyMq6J28tohUDkl9CUMlTjYXY++9SGOCiQZH5NGcLStK
61hiMNAKiZQhALz6SGkLtTgiLtcvLfz2J25aTuZtF7Go/c9O8WbOgurOpvUB0JpWKS9/Kcul9sZy
Q8eUSjr7OJJ9Vq624iwMCWLwc97tx9mroXPfj0ThrNCi9F09MZu5Dulg5Lhq/MDLV6FOwTOlNaGO
TnhiBpaASd0RUkHy0N/vJ7Sv/+Fx13LeVZIOlZ3rmLLKVKmqjMKVrAi7UzH4cd3fW3R0QOLVPtOk
F0hMSnQPjIuiCJ2uB/ziyyo3VgN01Fgc+BtA8tRrLylkdwDh3qGEbFvqh345kOByjT9IM9P4yxD1
sERKJyYobJnnTilLS3bbcY8C/G3pmwKbSBLR5IwxdHUBl6sFGnzZWuTJSekiyhrNI5qoojrJATiJ
z7vA+zqoahUkF087s71KeojWev/1bvKzY+AceZqqSe0WPX+ljz+uvIvuG/gk/Q87icg/Eq+bwLqA
2b9o/XDC6y4iniufZ7GaIBfHiRvDVg3BpfdfwCIdJgirmAVwtpmWQwRV0fUBzMcKWs28RhdGSxdD
jqUc55PSJaNDT9L5dJNrpsqdFw5NTaTMpXDJWLHgdwen2tZqte2g1yrfnEoB+Pd41voz9O09YQsD
YEJPq3i9i2wolUVzWcPWW/i0XoaT0Yo1Uh8/zEse/1iX2sKjD5b1cqrEVLiQXZDhA/oDryulUSBq
gRl2UsryZR1OEUreSt0ofMXYiTOV91NucBvOuWqTk1FG0RAGvtcodSAc4+wtuYWnkL52GVKZ8WE8
Q93zp3OgntdbyWAa/16qdtDkgV9AltaMoT5HQje88Tvqu894Pxu0tnJkTv6RpqFGp7QHuuR9NQBE
qSDkC/ZzOIGSzqiS6oVsq33uQEB/c/vc+Uzf3RU5dGofFokzj+yqS31QxPt3EjzppnMoKHn6raBY
kleaeUlJPlNquIAwv03ZV3PH4tTibFtRKrNn8mHqPQaOfa5vxNTeWFpXIgmYbpJABY0nr0E5gdHB
XzBECEVHWJ4m3i0NDt6eJk3BC6eXAqwf3ek4CFBP+PHvf48C3VP1T8u2EYNU2lUmTLBgOKt5C88w
4kc38gRrGriB9dVBCOFqsxC9yDHIpkrqQFqtshTI1DzNBa/CDdchlmOXouCn3hSmNSDt0mjfUMIO
MvXx7VcFhlGlp1uj8/fY/qIVfPrq9gkgoESCtyknJW6kl2csiZADbs94oDQsQF7d5J52XX60uVba
Q8QyQrpWRseUsECSYhN4AtOGvIn4Xa1p/HUJasD0Lu1ElMJclXWlsMmN/wY8TrbX2wf7X0Cmd+5w
4ilze30DBvfNZqqVCAhdBQhWorLZj2xjM9D1BMzCfB08Hys2gNt1MzCsmDigqStKQK8wQkxVBcBH
TXLPqGAX6f9KzW52Tly5MeZtYzne4DOG4so1LWQ+M+nhnOP9QtKvGLIGORSf8o1K/S2Pcc8/BW2n
XDFG2k7ywKqciR7pIVI7Xn5F0lC3YaGzvAlwHiXBS8J+Ks+I/YhImJRip3Nnw/hlPkqPmcwNfR+4
EZ+LaFxoBl5A+fli9UMjH0cY8rGgq5jvh1JA0TLnOh1m3ceLIeVgLH64Fm96nYDdKv8wFtk3sJT7
sptlAL7vrqOLYckzmz39go+sQg4u4ObgYfiVIYstKm5IdB/O7SWGHkpGfSxbT5gndRJ20i+3c7WY
2XMr0ohn5J6kDAkh10QDdK+7JVNHzvpc3qfHZ+BgSbXPcm7wQK5CIVWa9kYZmA6TWwsl28zvdUu/
yJpk5w2LjNUwg/Zd3cQKaFcdr/TQFLc9dsAxvRgc3CdTq6xVj5gtbF7P+1AO1w00jTvc1/ahXJKg
dB1snmgAQE8rTuG4x3Egw2IGzuS97DNWG57vFQ10t1EMxUNnFyMUzaz4UnL6avDb6yjeVk98J40s
TZ3GmHk+9tAf3on25eknmOFKYXcHsTr2A+FcfCLzfNMiyi0ggJEDrsaz+du+bnRrsh2rAyZDvEdD
scf7K9e3WxWbyt0Qla2qh301rFS5fhrx2hlvKqDE2JBU1A7UkBEK5r+k5FnJMNinTKXIvbWuGyYN
vpjWdarcq1joaoYGqJaoXLtVYBc+z4Ovf/sXzLu08pSBaWVdoHdLvSLVyejNiycXB8G5SOPb0EwJ
UsbyvxU9JwVfotq4QEE6cZRolCrN8zj/jYsOF2wHOgf0AcWxzmLqSJy53+ljMbI7BWSk9YFbgaDc
DtS9kWr5hlj/nNCTF4RILohblqNBCWgR8w8Ps1MhTTFea1vBLRHYFnKkcFB54lduYUstT0j2c2qe
7Plz2OCesABmHs1evYEqp405ZDtmMrnZ1vt98wpOcK1zbCCBI0Dch17DTeF/8rs4yqTnJA1v3QkQ
9qCBaipT1LSBw51CKYrh/8mSRGcIAB5wHvoNMxiugskkxhu9SkmqnnLJDKZrKvca3o4zN8JnNCo/
pvJHihaFB5uEsNzhe/djWAzGT2eglKqmcr8MXnpClNrUxYNB5Tuf8GkHAmDcK5voxp25lwmyaIbN
1Hc15MlwHWSOEj/42KqU0Q69gcPOeC3B5ID7JelA2g7L/rW9RR0pks2zRdTiIjfQmlNQOMch3mu9
Sz42YEbc6irDOFMJa0ZwuJvMtjGgPK2+KPzBCDlSiFDIAio5zaVDElR/ToGq+UWrNRjRarW2fM4z
Ao5uLyPt2rK2+hElj1jubyTEnwrB/xgClSzvYdxzNG5M02V04GSHRRlVQWxCa8lM9Ju3X3mYwBBJ
Q8/2Uzvcz8YlgiLrI01qH1N5vDeLlYBC4pcc6DpAh40W+Ag2Mr9D8leY/ZyR/NrGWl/LZ2o2MAvB
5LXL+7lJ37+BmUSCX4eYqeKQiYN49l8l8solMmWqpVEJIbV/tUgIeW5MzrjSX35Ri5DUkybLX1Y2
smSOSklZ7Ung11hhuVZ5JxDRxZThukK1b9m2r1jgBtO/5nDGYlNkR04CZy23PMwo6qIQMHOAKbTH
46JWshllB+SFB8X3MmcG6Smk7HguIpYtNvfVv+rDlJvBALOVzKvGvrBWRM8IzDd8qau1+p5zrOwW
AlqMi0n0xbX7YDUUNH3RMPeSlZApK4zsAX6eZFhcEu420lGNgC8Fr+ewJ4KFiFLlpkMDOrOkBIpN
igc8BMzoj7FUnszPlXEZfhEcHs0lgB8cORXsL94yLL1tbq7GmRyrrPfxeN4rVWMitcDKtfLQthzr
M+ijM7aDF9KqzPxmaWnUpxfV4hzS50O7PGMMB7V6yR57qIHNok0iWO6NB86wI3+5ZLD22rEYPZMF
tkMHkM+fLjQhYfp3/Q6vtSNcLAvYFW8ZRmbnZJrM4TRYIulP+0rxMYnSsXVaejEz9uRPdLvQT3KC
jeR0hDeDecF5XypsCVmPdqVGBJ3J2OOgnO/9ZDuR/D/4h8rHXN9GD3J9YUS2dqBRF4t6FNC4mIha
fAnvvxVwTXvuSK6oTqHOgC1Ri6l47gSV4YHQi5MHxOUJEVYEVHkESLBpQKGoONu6PWtBIjzEe6x+
4JJhr/Vad5v7YmV5Cl1SRe16ZFvabBY7YHvEUkC2Xxm5R5QmR/RlEfD1sHI3x6G1TkHzDfEcFijF
N+PuTnVpTEJfupF/aKLATOT5S+WP8PG+jd/tYl+LD9zmP44Q0Fsdy/g/LVXW2FS+qju1rQ2JBdtL
yvuePIejtcnhGsztmCB2RNuTiQj0lve/06MTF+TtDSMTkF5NGKdPioWY/KJ31KOOwCIutE+oJTBw
OlnVrnLJM+MalJN6utQBaOUfX/QB3pHtnCBvAkstrn19InoIgCevL4LqnZwF5+Yzitz9eaYvrwOc
yhUJiO4+2ZOd8fM+97NuANES8463DP3YXPQVETmMvS8QzNuuCfOQqrpFF9H7H33G4oe/kjkT8/a2
YXlHKQYbkXQehm+kaOQQ9bD6WIBEWV6GQC5ndn6tgdzJc4nbRK3fK4N+KP/Id/vV3RqTvWEnNf9v
/60AFzphas7O4L8VwJStPG63VAVPL7c2RHwGzP72wdTIqpRC+G5M0IbSE95IwCdkeGVRH1I5WVOk
jPt36PgkPke2iwpEBuG5arYwHgQZyPYOBZO69LaTUCA2FV+DX+k6bbDDbdrCBiXKUPZeGf50dq81
lA58Cuv209VJioUcqLgHmIm1WMvsWJZ3FCd36yDR90UX2SZMGcSpVu2rqEQVJvbj2Nog8ThpLX6P
jv7qZSffdnv0bI7Zvj8P6AgqNiLXr0FDcpwigvkOelUALbFAPYLZjVYFeCZE5i5XVA9oQViFvZ4X
5QwAe4Np/4tG75uwKnU6uDgwd6qgzzTW6ioY+C3lhv1w2r4u43WMCvCviMk08R2sDN2FJT/8VD3T
ZAnNU9cl0aHNVB2V7Tm3a5PUzbFpfqacjCJll2M7Hig7scHjb/VR8ERqZ7zUtMtBxI3jwEmXd4Pv
X9Ql7LVK2G4h4g+IDuYeP9cgB6DhiwPBpSXjkr9C1bMl6IOzDl0exUToracPiH56/OypCulx5rgH
skrs3/ahnIKo4E5BlY32G1Td9Afz/9Iz5isR0FzVdl8qPqtp2Kc7ZcQ2DlrICtSSFaZlVpRKrv+P
hwaSj713MmRcxrl+Il1P5FBnvmbpQKX3uoz1omUHwABWCYR/+snOoX98IapapFLL9fttB2hqARdP
fI30BMepIxZ6Tc5zRvM4RljFDX+C0tB8JOoPE2NbiIRWK4/PRDWQdPrWeFzPJ8SfPlJ8XHTF3Mwr
4r23kNlAV5uNkR4H8sngBPP3O7VPHvhqOO6SHZz6yVSZrK/uO5Q3x0HE7LapwE37LcjkvziceHaR
Kds8Brv1SZzMj5mt7w2HtQFLG0rWFX5Ej9U7vuNlrzneXXt7BXM6VZQ3ef3rVVtnr69YrUA05ft+
QC4BMDx8d6NVe//cA36X7gsMv6RaI025blt6mAdLNuv4ZpahF8Q72u+bpMfEl9zrF9k6ptM+TkMk
doPdY4eay6PrQVqIHDUT7HvnxUy/WIxUr9+0VpPbO3YA6iOzQtJhL0g4FjSdGSOlEsRS8viyQEPy
2kWUUhQ38F5LfjkoxfsWi/xiTVYOMaDn3k3I1EZ5OTm1q6Lud+2Vm8FiQolKtGGoivoOQ+vURo+m
iMUreSqGHzPfXQBAvM0K1QJp80kKl4MEG+qnTfkgWE8XnTQhJZN84+TpICWlaasW2x5FWIOB37qS
3KgYcFiOTkEZfG+pNX3vcb3QdPegYytLuGJexMtbiDqiiPHxfIGS9rOsgiTHH8vpd+S7IM9XyZAq
hgt9+9ICm8qF9TUs4pY+50fSpa3QCQGugYXI4fdy/B92bHwgswCqQRKsKuTM7aed8tFQew+Z7bz0
HFQteJh9i0K5rSGMrNLXfpau6gBJTtKXuym8RKGaUFpxo1j3QgJDXUCAVry8loKj91/6AQtS/GQt
R5IhErYgvslGEj23x7Ft7KoIXdFFxKT9pwvGXWccmncD0Wmm/do3rKjNq+lxwpcNt94/b93w8zWf
547dwstB+T9GwGSdBpLz3Po9GN1HTaFbZyAiJERGmDkdIUnjrGipjd50Y670Aaf9dmXxflB7aVNc
hJLY+7BmzPwtOH7Y0E46kQjEhwtYV80LhlUs3UB/Tru35t8Don0P/3pWQTvHry93Fg9e02DoMOsD
gqLwpjMsIgUSI3q/RMkQstDjBrnQCB/eAOIdHmdaAebCrHiWUQMnrFTxf6M+pWJ7u7/Xd6IrEeEk
g4j3idbd8bc/xxfcE9XVE55Sxij4OkIySEPpLL/Ch4dXsuGCBjG8h5Jdzc0Ex9VpsPA097UVvKDi
jE4a/vghV6nkITiDqEmEubmfqQd4mr8n0AifwDLNMZJepcxPfd4NQWBmEQrVmGzp3cPkIx3fTAPN
LuvXv3xmvvlRRpdEZcFQ+Ih23MJt6L360q7tNnUKwgioCSVwKnUBEZg3/JPF+Qpmeg85gl2ToG5W
69eYCG/lkHP0tciXGEzZ7lpjVUiXrJUpmC6JDsRoygkeGI4oKBxBa5ptuxoFoaBnryBMaVKHbFeP
crVidtLnMkWPyPkIQ1wVm/zUNhxnQzlbK2NxdVlWIAw5SmCAttwTMfbbwOCAAEyrxRop9W+fjbsB
rofLipQZVWcxaY0L1CpJ76JgiJtZR5skQitfZjJpOT7gTugarT86HuJ1lmc77hVIGhdnL8wuKi9N
YblVxmujK4L6sW2Pxq9H8ZIvaMerNi0poC9E3ujbu3b9/WKwRH6qR20Ji4JtQdux1RIOE/NPGcYy
wx+MVCQhg/zC0xSHjT+967klhbNE//6/U9jeaF47wYPnoPa/7Q6VDw5lCDvtzX86RDCCPD7Ss7x9
L23GAL0YM7AfUHTKxjdb5zswhUlEJoZEeiqogXsZXdXguGMy6Qi512pFlllz1ryiCxYiNJYY9Ewg
HuYA4gs317L9B4DoL2KLTXL5bfDzXSfkFkTG/VsHzRRs0/JkUhQ4Gvt6BaQkXoTX+RVbvwOOemk5
vCBhJpli0J1uaXOM+GG8iahEBltf8rg9WAo5YesVxZh++u8aaPzi58E8gqEY3DeWTCcSJGYaMr5x
Ia/jVjI0pi7/zvwdq6kVQm/1j2BgDa0WaYgRzmOXjPFaILhkctRlvxXXHciNip0v22T1GjiGcWrG
H5mzJqPQR8eTdJ+BpeYZYNJYRRNFSkGelQbo2j/OFt5qB12ARcRlxwcApSvnk0Dvk+AUyE8qBiXN
mimuunwcM1ZFKnukaBzbkoN7WRE65qo3Q/nOUeF3Q6bwoc5gIq7J7msJKisxiasL4yS6M0tCtohu
GMhaTY7RrHHMmtG/L2th3ttA+8NCQCA202gLk1omTXfMxEautdGMwodGTQlvMCQILJej4/eF8iD+
mLcfyXUllmgHXktKJ4RUni3xV1e8JNJyHZTN+b4QQ0KxqMy9oH8B0msAsDFVGbYx8mPReBuP7/V0
8hUoVIfbVaHuuAMqEYE29l0QN1AKcBXEp7Qfvm7NfzXVI4rMpw7G0KPVuad1ye8rSjluCmFmoV3f
/w9BoIr1nNBk1TS24PIRaZDpuzuh98VnnCMqeahusdLpJzqwIe7CdLqtaUTKQCwjg+GTFsRxnaSU
ssAd7kAwrMkKtfz94ujYKUbnx8gRSU2i2RJSQpUc4ahsgUrcu4y57FeeTnVr0aB/UkFb84A+bd7p
bf1tq3k46I7waAYmmHzFgodj0GcQDvNEfphlzYUI0ftzq9RDyAFfhQpvzyyZ68B2AYkKBDSJ1GCe
Ywor3vTkrzmz5ekHVsUQwIsxcV6fzbG/+QAo5lm/RCmKkEdVC9ApjVolRidPjmldOPyEr6q2ijkw
0+0k9duyWTxP7fUAWZzs1eYUtLEjUon8mbobKkP2Kd0r0n7J+RMvnaOy1VWa2mZ+X60eJHHdGUFg
R1yvf2s1Y95lIdXG4mksRSxsSkYYM1WmQ8Tusru+cZI25r3JqOkyEz3kZM7BMRMFUiaxdpiimbAH
d+8gYTFj/PkNKLBu2TpeV4KwY7BgtGNMc1lUhcjQO066XFO8i+Tr3RSaY3QdobENUf7e6iVUvIPc
S8ozxPym/xzaRrDLHqeOZUG06wPu1FcoWZ9le0JsiI7pAXxTOtc/14Ph8MIZ3KEIEnpY9lTH6bs2
uk+sD4e3OsThuCdPr3NPDkXKYW+1msNpNvOmDsaHdYfbIJrXj90WgL7qHDZKd+GXylaRf+lp+IH0
BvRKbowB8BaHUCuHbMwMM7VpKNoBOQ/0LidwjUYFr2FsRjrEkTRk2TBc3AQOgA/vTfnydf5VkdSH
j4Pzz+8gpT6Vm0aZFCK6jfmo/4goCHur1FaUTg0P5MlIzKO6qXS+sOyHWhu7DemKN57SurqZ3vah
gJT6ERRrGTYktnWLNVuliQW4qHNES3ViJL2DUFiCVrn6xNzPYEZeBhvVM7GmYpb2yDS32GhNy4nz
RFz1yZrKf7VmsetLCP9/5iIDi3F/P5wvg0hbmxQlItp5QcM/68Wa/G9ViEfTxZwW4pSjTIaHsZ6I
CHy+V0Lr7r+bQ3qKKxSntjtJKn632/Yk0SxjwqI6AQ+1tlhIDwWbifTNGCNuz/ldgUfCj2l4iwDa
gxvRe51DparMKL2Xc2T2dLd2rjOKIJREGx5iXhwbjMxsYH8aHDTmLNdsMMutTT4ya2h5z4BrkdlS
fQjL6RdmwPjUd3S9vmMFMuSumUF+EtNmLiyM55BY860cyUiFNu9ku76ddFjQIQEYIN/TyNderjC+
1P6k/zm9vLOD6352ExPJ/SQEC1ERoHKOu+ZeQprT1/8ByG4S1JoH/mbdwlPs3wli3HJ+bSstEYeM
+OjOWUVQOTXuc8OKq2VOKBvnE/YDsZCqsajWcgT45yIt8jyxJDAXUCcfJBdKw8qWe8ov1J2zbrv9
kNBvj/cNj4l4ATUUSaH3hKmaHrmsZ99XLNlzaDQKngndqaSKgUJ8WI80wgFofZ9kUw30v9kQiMh1
XAxqB0ipoifeo0bcPvZ/33ZE4a94nHbgtpWMcdmlbeFA8TgyooEqXl/YPOHhm/OCKuVP/HAfNQcg
yASYYc0AZeOohzHX+eOpkIh76NKZ8wAJIZjKLoHLp/cAzH61fpf5WyDOHDUN4ivsLmhnmgNegOhx
f/tZWKmW9qhIEKa5qm42lZCK4VNklrOLBRHCA+0lkygHYeo6aFEihQK7FdhkHhSQGGX8tk3XjxHU
Qxfm4s/p4sYAFAF+cAuc+DYEAc968WjXh2Pp8sJ9ClhHPeh3wZLOVSwF3+FOcJ9099+AurRMXByj
PicMTCA1tjy9a617WsOKg07+3zlAQxH4Fs3f07J1i9L07PqF1RNsqJR7mrLhgy4Q6sdcAbPUlKFc
cdL1arcQ8TE7RjJAPOT4Ob4DnQlwkTJrO0vYRk7ppagm4203l/z5oR5j6nfc1xXAUdRievGhV/Gr
gb2yAClBbXAEIN98IUA9iIzy+AoFy+dJSUQmdhgf+Ku107l9gLZTcn3ayKtLnhBfuaVmYUp+iiGa
EGI9sPLMnGtgQGlQZcXPjkTC9jWGeysq7yEH6ykqeWqozVqNFnXmYxYztciAoJ31L992boFBEed1
o7q1UEAEeZVLT3Fpo0UVvdC+6WNyjT77QuviCsRgrMy+Yo2a6zs4esqOp+NeFnu0O5UiVH5xvZie
X1szizPtpQJx0yhTdPA99no4rmig7OULPqPN/JuYKYRIY15/154erQSck3tqvLMlACQGuASpDeK6
g5sGPMF3jzrzW/3WVyJiTm2JIZwpMGyautTDBEn/cTTHrDM5TQcBd8Dpc3bkx4vdPw+CcXsgQuhs
r44rPP6G7fOo7kpoPrnnHMJWk1+kJHHlqS/M7UHDaqL00/FObitmFZUIZ96rllG4EbOWDoozLOCt
X0BGdyAVC1r30CS6gqjor8hY5iZbKr+xoJlC57fmG3eM3/7nZOYLlscvFjun6OD+Z3oHpo/DxtFq
rqtnnrvFuUVXNZ9yJuGNCz2QJLGrzy3CSAN1+CSuOIo+LIdjfqzq0GEGF2cX4MpxNmq08y2L8HH8
NE0+H8HtdnOxmuBduTZoEbHIsm1fyBJc8SJYDlD8apTM6spvJO35JnUN7rCwH/psQ4dnkar/MFqv
fdziHKV8srj0Pz3GxBIPw773YAycPtl5aFa60MCXagGNjPpdWMul7BXP2XPA+51eFJeLfiFznijy
2qJ5kxTalm3O43MPPwXFidyAEQ30V6oG0Ob0WYVcgJLe4oE1XIeTUXSIXC/nAIJXchZuci0O9vnm
VV6t8u4LdWxWkP3xj4EvFCgDTE3i/vYYMxvg5xi61jvo9yoV0FP6FosyPuR6iN9nEVdEf+hSiggm
4JS+k3cRLfiuL3r+9VvdbRdTwvCze6luU2LJlcLQq5lF9CzJVw8Ub2r2bA+hu/r8BQDcAXL+tUxp
zNcGHuuS4Miz6R2pnMXW2BlsGvotTuhV0ujDGINgS3Y5r8W8nWZheeIE+UqVcN38HOezabGBCr/5
kftdenBORY2ya+tBZE0TkxkuHCBu7atgCnqoHTdUquiFXzQcUgxqB88ueQuTkS78Benn4iYKhKmd
6eVqJgE2hP2Ex1xVhwhUCHicVDmnxrrXL7kNmUiN3Cw3DWEwzc7u9txjvW6wyaUMQFp5hX3Uc/ZJ
rj1PFUcfCisYS+c9Wesgj7p20ohXKezVzLRY0EguUGSAvv8u5Ue0dIf56dDWIu61tleRuFM/WiaH
FcDALaaf4ZGwNdaKhBr54mn3DUPQ89YIOfXw8YhD2aA6qOGri6AhPM4YF+cJfzrIzRrRg5xe5YOg
ZmId8KhRySUchMKMzAYAPUn2b+9h3DDEmhlE3RAvRG92PbjdZm5s+28b0Z5UXZsegdcF9ZlVekjb
JPS662DZ1yIu57wlBFl0ilyIxkV0B9cDMou+ZLV0NsCfXvvvYF+DPO9SzxqScV11ry2kNIKvQXtZ
hzn4DZ6mBjKsTtCjBCDnElA+kOrMIIcxz2vLeYeNk1nYLcUkNHrSlrG6K9gx2zlFB3KJ1aTrSq9a
JwFRmhiNe363qaZDgq2qJTLiwtpiW4SmJtWji8UWEspI+AyFPtKlCIvWxfIcX4H8k0+pPN/cYmWx
/hZ4DUk1DSf+RklYy1tQR3LI5Ru/DVTKA5Bjs6FdshUVMkRMIlMS3bpj7tdcczdgl3TW4i8BHUKO
Oab6C3Ry3FS/7+ebVObdqzx6T5gUmxM0PcQZ9Y6T1ucR6phkhjcxaPh31Q24m44Dswq2n5P0kJoL
9+x9/cLN+aKV8wiXAM75ldb18VaQvPWJ/IbGUO5BNBGf+cUP4AY5BUEYphoqhTGkCDpIR//HIjb6
tI+KH/jcvtZqdtP9UrN/1U3CJR+uJeGGpB7F1J2PGS0SozvX1L+Z59/rTZduj8lxTDnR+OnqZAWv
FMd3YpX5ll56dUsziFyzdkKBgHQkf6DqFfc/F3iPT9MxgAx2Sv5Uxkw6MHvvE/3xf+HeCQCkueiQ
KhM05Z93n2eh4u54Y8up1dy3N7oOxi9TuibdCRFDp0uSFLha/Gg5GPfcKR5A2SLJIhAnbakg5uuo
ARp9czVbfg/hKg18LknKp7CKKhhLvxYOex4uFsbzIFUq/BAfuSTDcd6NvtTUDVZzT5EKuNyYxw7j
8L4ptqlBj1kRIZGH0Y6x9slqp4nawEh4OACWB8KBq+Pw9MALea8goQyVqE65QUYVhbVtWiHSx1zj
Ppz2xsGli5dd4pJqsPobvShH+fDynNJk0SaO0uHJD2jZQ5gT1+arqN1uT/EtZEfv2eg4Z/dNKGgu
r2dv6T3AY2X7qrqlRarx9s3xN9NBBppM3GZNsgAtHemQbvlccYTQPzPGtkBpTUWL9wmEUDr5Ovav
0LDPpdvWeBDXShcyOwGkyGWlXSFN5srTlyjlUNiO4VjNL8/R1s/QkmW2lRUkGdE29GJWwSZgg4tQ
b+jWJXBQsIAGR/Y1Y7kiINpdYF8q2UjV0SG2y+8YpG2+gfpNrSShyufOLPXKtTI2cnD1DdTSd6Um
NQopWZ5q5QklhW0mtLFGTpvEYF/Ao30YUh5TIatyvBP/WZ1dl1H9d2gCMAi09xQ0h5pSlPADABSX
LNgFvdhvzmuHIUt6xbEH9rmv8YWNXsyw4/4gyr9Aef7Sj1jv+whTcEDWlp75lv87SEsIPwXWABPt
HJjLxmT09W+Ttw28Lc9RA3W/5Ju0uKWdnfj4R1clJELb52c6/WBDD02EmM2wEbxM02h0ABySM6k+
Z6IcIM69VQOHx3fSYt/a+vzty7aWWBaGdBZZk2iUFxdP+6+Q2EFaty0y7yXwumzDMrAjzkzkGF7W
FDtUpNMenh8ZdmSc2fCeSj3o4aibjJuRvKc0dNiOzZ9LAWPSNWWN9/M8/2sKZNyByoNlcU5eDUT2
3KXaYL7+4LfIjNlVwsCMobBxmACkdPWJAneusW28uVMurO+ykhDJYBFsOZsgnWW728SSZzhSS7MF
jr3vCz7bJ+F7qROrkaP/yaI4aByj+0sLpA0x3epP5KXdM4Dr1DK8x7y9S9xxZ339L0mnBbJswD0g
1FPptBA+3qii101FwBFQ/e38SGwSB1xvqR9PNn/j8XHmJIZqzY+H4Z0ZtlIMJNnAWUpSWOC/K8n6
SBlvf/LGkydo6mmMJxZcAm8J2xiEjtWnhfLvn1WdoNi+XWNSokVfzvhKOoasYhaNC0s9dEPAyC9A
9u1J0RrAhySR+Yl5FqwV/F5OWKY8m9bKa3uPAhXvKsRC+UfEZ0dSnXE3kss/GRKhFsJU2JbG7eRc
swoD8CPCRxTJCMGaMRYviAJox62L6xKRVXw3lWPnt1Az4l8sZY9BeeGXpW7KzFJRaEP8hpJpb+t1
VyFSv23xM0rH6Y9H5CsJXnX3DMTzWzt1doOVg47HqyAjX71WzqKgjnZH/ci3jVjtL+BdpRUL9tiS
qOFj2g6bzpBxM35Q1et4t70a7PzKz9Ylrod8M+mefmu9w9HUBEVB/pGQPqK4HK+FSAa1bNoxY0wa
PciSmpFka0XV6uIxNfB48axdqIRTDFhqH8WFNhG3k5E9OJNY7fl3HiZInVFQ8Oif9V0crPhHVGK5
CzxNfHmDFeGkcBGFpD+Vl0JY+WErrCOQyZZs1i1QC0837h0I4gr9dX8kJb0KnDs6lQ4qT26qHvSD
3tVvw1Jv3VLCxXP/CLcOjJkSajJEyB0obCr8oi9d9uZ0rlci7bhaaMYeb1HgrEIIYTlEQWnvC2Hb
qalCLh27DZUjQXA7U98UcG/5F5TUjR67HoABNRauiifep5mAa/yHmj6ztbj/ph+l4AOhLiwkEJJB
y8nRR3yFtGoo+vcYojWHiLz4mTPqCShrxRqC/455YA86gJdbgaI6aLoYzocI2rTxed2elnJMlLf9
70c6fdRHseNqlv/JYDyDijMRhiodU1aAXQfU7aZplNqsOHsw4LqK+7j//gHsJ2+BhT8v+6DqUDBJ
rMFkaOWohhwOP6BGL2ujXgz+QFwvua8Ldvb37fER+fNXnSTeQQjYFpKEqdIQAF7z7inzfjqq4zzj
CwVr9Zf0jdBE9kTLzgRGMoQyaSfRcyDZp03eJ/qTSk8++HqKYVm7SBzD1bYiTFDcTlp3pnETWTrF
7YtZyo0jJGOOsQI5b3k9mEModw+CrQNakig+TScr57+iagCxyvCo7+T6LwnsTK0579+gPF3Wa5EF
PW3L1HHRrjGCLqzX35O9D8wWNlW2Lh25E5yIwze00pjVJyWVmFibHcuq+I0Vg4yzxDFbdYXu8W0x
D3tnrEg2FgM59UVo0fzElnCnaY8QGipEA+qGZ4h+WpuYuVSI25nER9qlBaDA8HbO/wPXbWXDZ1Mf
CuGftyUDgBl37cuhOIEDddjzhGkZ0FSI0SEb59HSRy0HQ+DfdnbHbHE7TtAPhS9nfQslSn55b6jn
gNm7Wlqun0CuFDMgpNGRYw1oBZos7svrSnUaP70A8WzwvqdiZMu1ft2zOoM/2Gv08YM0aoSYbN7E
KSm7+q6rw+pzEc6GDBMdKGe8kqL8WpdS2YftyAro8kSsCtIGoTggGWzxF8MRAMyMhOILTBPFzoPE
r2IF+Hz0xVYWlcpRt05ZXl9n/81axfeRT000jp/6j8vl0RgPBfOxf7khMWzOjLDoiOuLQ5IEXHo8
rHUHdzaKYpYutYSddGLH4F0bQ6c4J9XGhuov3T1NHe/QMqAua245TeuhzsO80ywLCNsWTQd2Ohum
kzncq/oJjSOjqqfEt4d+hIxHYmQeXBs4f9EJoEt9pXVBaTG/kzs05uEiWaLdrkXsMv+6mhZCPWfS
AJ8AdOZ1EHxG5oEU65llU+B+P5binTbVNGMzS6TTuMgrltnPhSSRriyrWynfNT8e1TRozSRAa3Jp
FEwBHp7Rc47HX/6hXVTt+1wGySjfrbzMq34teZyAk0jEMskfbcWnqtV6ivo4R9vphcxNA0A339qO
v6Gd8jRCjPtiTYOc3/fDewZy4ux2wjA4mSZmsmr/H6pjCB/29ag1SQw+JetRdm1vG/CjHfhTCJZ+
VGJ9DT5YrfxRc2JL7AE/wg0sPh/sdvLjYcmkck4ZVhV/5AT8xHXdhUOTUcWj0MKUSPvIBhkZeGNS
WMFob/4JG5IcWZTsowA/yxU5LIN/2HzZPd7mbrqJvtc21cZCYkpRqbFdaH8XsUphXgl53Ak6nDM/
6jfpgLcEjBJs3Viv5jdL7jck2NqBw0dMlGaFzPPTUad5AbZ9z+H4r43NEJp4tRq+BL1PxNqqYJFH
i/fqJTIzHvTYzQQVay4zHcmiiDwbdteYDaJTWMz1BE1h+86GSv3514YXDwqbBusnYswRokDxfRuT
kPw3VSe1QKQjjELk/EdRgUTZawLMV5JX3q8CDpvhPT+ns5iTBCp1RiMmHuw2xepBtPg49pV+JRyM
B1b3ZwPmEVGql2WsEqG5o1IXtfpMApjH2bWNR76ab7OuDN6Trb6nONNpSAv54Ad60EfeUhFPhVeg
kLNXYgG7iUNkCtb8Pm1C904tnGAL0qLLasIl88QFfqscd4lVtAag3Y9u6eRVGkcpAbnPK7OWFMzW
Kcn+xeEGvhqALRz0SowdTmYKjugZ50Ma5C53eacVIqYOyn1EGTtFbU0XqPZ2MvsLv31hUAynq8Wm
YhoRrRLYFqZNvvdCDnNzDacRi5Lltgv+6XA3LdLxyDBAtZC5u33CuG6QPljZ9C6brGddjMhhqgPq
i4saKQko37gC4QO6jP+o4oNAqtxzF8ds1cF64arsqwk5HmDsA/ARYGB0HVVz0tEUBue6mbSnS/O1
4a1JaPJJnT/y3Odsx4PrPTsxpk/0b90j6JJv+3lomrch1W1wWBKT4kzCRdJALw7RI2hNnKFhlwLd
nUc19akn7WM7AsybOrNcs/j9NrSxomiaiopyLb3C9zd7JH/Xicbl590C+vzIFANhr0FAXaIClE3Z
w9QgmmMMeyAVfL1/K2w8UPf2kcfN6deGSxuiQUpDRQyszRYjTULeQjIOdmpY2grT73nImrBnc1aZ
m9YAks+Y5e43gaDoMHlKsJCwpv9iO1KaktS9N4WUq4kv7uuMBVGQNG2hYAue8jYIMonZ3fG5U9wU
+DdiK5DA3kqDDapb+Y2+EveSbY/v0J0kk7SwbMFa7BvIU48RqNoLAqR0Mh9BBNY0RSiqJ8fpBJkW
cfJRz1HiOAu8Ho2LlZmLXnMWcQJ/Shl6JZAF1Y5cSOz5GC5bOZhIgXsFlSZzSOjGrNMUECflPhIs
02IQmfDeo+ba7M+kAbVXmVHotYDnFcWlXvnIO1RDr4d5Apyt9R2RhVi2xgZuwUtggb8XeHGxqPF6
Hynz48OyCbfSUDiUhxiV/Yl8Q7oE0GeEZc4Pwj2bqh+17hSKm288VEfB2UfFIniIA3vih13iXM8I
whVpknBlxn2j5GVM8GnNxCfT8E/wQPSVSAB6rlifJ6km37S2s+dKYthNHThcguVoqvFq40CW0E2I
jSXNLwEszEpWYgxAWuAQY5B0v8Jl+sALZ5FEt69rwJHIZ91QXOP/JsXhLBb5julk/CjlrMji7uxk
WAcACaRaP65sJYEuX5vWut38Z8kg3Iv8xtAy825QafxZbOOGPJt4geG8UCTyKCn7mxJNpLRSRZpr
wDTpT2JjiOazfUosRGNaJOnnYHKH0yNU4IlLrJbPvhU1VCbwA9SDt0A5zD8m/pD23kImGKrmEfd0
Vsg7c0HLVWJ5Lcf7pAgqRNrO4l092DikekromSbfaSb9YrNo9nY4FHi/YMLp3rCNp0Mw2eRS0zsF
0xMUlgN72I/+lbthhxrqYk/fDknVb7ij1evNhFpyLxddeWwvO1mbw9zxFRmi83OU7ts1BRKkNSb5
9ZQpKUOEVJ/HZfjBRlYqqAKkzy+RoVjLcgZ5QvDTwKZbbR0E11gilNG/Jr9+C+jVYSHZINO0AHm1
4Q+zeEEdMtJeMcwkJPepg1MjN4b+fw7SZUIAGlzKHdlArx4+2+iFRfEEaN5y2q5tOhmV5IwK/cnH
gL/R0IGZFcm/xp6HAsRozFENDC2MB79bAgaSMoP3PbwLk5I6Ldc+Uz+qYHFSeJuORholH3U7bdoy
efRTerWgDaLChBl8KvbmOxkOu5TZyBXPu4pmqJB4bX50DX09filJsg25byAItJzQGkEzBTs4ctYI
p9h10olFkGL++GoQUJCex42GudcYbRr/lTWsgeln4U07Oc7YnHzxpeaCIEU0i5rSdes5mZW3asof
cD6CaEKYO7M+Lefh3fkkMhV55shTjIZCEKZyfmQeG+o3XshnJSlLsioNZ3ASVFCVbxv700ker3UZ
FAYIOLUPuDmrZwcWVD4d89emilguaWHjZxNRlJVsioSS46lF+NFFBkLS6XmbFNpFpkC6TKycUXtg
GfrNEb0rbBIUKKqXPJn3aOFGU78o052fVbu59EONvw8g+h7/iaskslUhnYRB9TRO14KaBsqkS1IL
UiUtxx5ay0ImLVSuy4B+4kZS5LXwzTfKzhA1MyEOvdBfayBOHQ/N4IkNZkTNCcfd0yANfGMonyCw
YeWfeb1jlikQ1BbWZxtH0+GxLGvYgScBR35KrsvgsScyIfyGKVO3cRt7rMr0//iZhxQLJWM1Rh/w
gxXxou43wmNAo8NXAWgXZSBbGeiSKAgUNY/Aek/g/Q5ssuK5bkJtuukmS+qDelUab1eM0GTxZMYn
bbQufOQG/4dMYhAYmYwJW0ht3Ukr2VhEDCyH/cuPKkSnqcYr24VAco4ylJABPr4lON27OjaOCEcr
zeDs6SId12rIrG3PMzoeMlc1UCUB/Gxj+mnFa81CTYdw1mJQzL6C5SbWXMpfR/m3BSFS75XcTEiL
IesuMxtm/l9zZq8katD7nyj05zdISMPVcR/oZteWheGnVvohXoaLSeNtBXk1d9ox8Qmbw7Vacur1
DN2EXTQQpF4xrKYGyBzGT7Vtj9WDBOT8zeeh1VzifEOYmQQfLFdxNTj8I2vH7n2VtZZZyh4s/m5T
4BKj2oFuoBeySzIk/okcQePWKpqDj0UkvzKscor1mUGUa48nXWSeh5pxYQR1u/Ta59cmb+/fzVvv
b0DnHzwhWcxjx5cdjmVn5RNLcduqdz4qx0i6RM9Sn0cvTpy2mfXuPscHOt73x4EU+3F8iyI8q653
/30piTkoGFqqUHtiJn0CfC2GGsvn0GuU32xfzJCKKCH02a62PCvSwQQsB5uWnLi0mtYgZrEdaecX
UVxmeSo7c7OghF1S0M0FhZ/OdlOetTf8jlOrv6ApmpdXGI4AbYuauFZg0FORw9X9OzWKqLc+XDh5
HSMeda/5bx0WUhOPPBz9yvxJ3IkC0tuDh9xFnwejmWD4U85WUdLOupzdfeF5fe2I9TD2IBxq4mpk
ChMBDGMeniQzm6KxXCr7l5TiibCYCELgmiMaMLs/wCRXloaa8umds/oAfben4HD51Vxra/fu7/kH
QeTO9UGezMpHMiq4DZ0YU+hmAArRU1uSRYVLQeYnBeBpqS+q/qe7FFavkdMUyIu2CCf2098PZYvj
oMFKXxSE+FGjn11JQuYUcFLxtCTs1m8+lP4Ru3RMKNvU/OIoLhcXFQdZT5yVn91iMLOdfnMI4WDY
8npdDJl6FKu3vU/NU4G9GSRlRfiX4paGWDbbbmuIT3Da7HFl2UebQ+koeKBWM4oK29MQJbrsT3hl
sNs6ljMUM86HamU1KbwAdTgWeOcM3ZFnHwERYE/zOUo9SmRqToBQZpt357wNuEDQzCjmEOFsnLA9
HbdS745SEf3m8+Rbrm+5J1mU9toqxE1v/acwEhRwf5swKn/896Z8sHMIs6/pLd5ppsh6OMSXynwI
h/MjIFdhfExicLQDO/ND/2X9OToKOk6oO0tln1llhFdfHZwB62reCqGvjb1t1LIqqoyMNm0OPMv6
wpFjurqk8IoFqrkX6dwSnKPVaC4hS2E+g4RcXvVRdT3q1EyPpNX46nPvJbBWw5BlTLgpSUlqKv0R
963xVAgdqyQ9wLQyfUkZzJ8hGZfq2qg24CUt7LqM+1AK60PBj30W0SWeNw5iMpIwK66J1a0yzjI5
zLi0U5fzj+Xr8i4ulRvjTjfECeCm4/n6zsCjQJAuF74fHULarYQ0YpYmVSxXNEcUt4OR1AUulQQz
TpJu3ACdsnfpt+t5KX0MgaFBBgecCv6Ead9nhuyHp7ZGMzWCLYUdy0UJ2/ZhhICdoipUtT4HoeaI
aYgBb1cJB5LRRmra52cJPo0SblEzzkfxcO2WjqQqUs+mcPglYT4eLZ/N+q7TxXsNns9o9YnwvY0x
7qRAm0uBdbvpIdeFiX3OaMPEAg/AGl7UoYwRQoUhynPms89B5bt+y6flZCDM6AH8bBy36o4XSZbS
LAM3e3mvbV20YifpHXRZGuDnD9nvMTAXBd8BAr9z4C9jnI5W6wopQdj9lnD7ClmzO4AxC2ILyAL6
Hy6havXdTQ58DKeRmFMwY+os8gfqef5cA89CR1FmTPo3YgYtp7RqpH2+5W7950noUgX5ucZqerGl
GkJnMrnG3Yq8t2k1QhhaPZgotjnDW1WhTekN+HbJPSExPo4iHCdQcBuy4XF/JD4nMuqvRKefu31a
QcYea3FarMw1dnHSpJdp6cZc7dw7XABnWXlBHYYS40FrHm9FjMVtMW2J9RTV/fKS3qeylFElQlSC
/elIhLLKAbtAPePVXZkqVal7OGNbKobeSBNEov6v3Mz2qvypzTOkQWIaPmoyZ3lAsjTeDebtgbVu
Ou4dnP6EF8pW2ck+2rk09ynbymJyon8/8siHRzCCR9WMY4poXAECkWLLyfTsTvm1fYll1HbZ0GS/
+mG6YvUSEEZ/+26PuZZ6FmsYhZBc9/ph7WK90jo7OCeCX/vbXPmbFBJ2NClZvxXdpjT8TOY5ApdI
7bqtzy2CyOyBwPwpc5WKowgEzXewukDQ2TPQfkN1oPxh5LyXNnidOmp3E4cQub9eVOyr9lCiRMSt
ghCzjXFWHL3r7amNStnAexBry7yGr7Q9hNW6Iz1uJ1iCnltmEjBRr4BTuOOmB+DgaozjkH5RiRi6
paRRHngTTvHnSHj3Y8CPceVWnX5yJzqmetItE+S8JtMnxhv+Ge2xmjMa68kDNxK4DZSkSnFseeZW
gbkrUI123ioUFwgJiNClJ+4HaSNoz/mnb52tBbVT040e3iX2F+Tu85RQEorgk2ioiDYlPLzOmdyO
6j7tbrip0AIv5vX2eivtqoHKtwvhTEPEO436FLhAgh+HBKpYc9FiA0uNP5XO1LKkCi5GM9oNDhje
U9G3lF0XYLfzG3w9pA3RS+4NVelK7I4kr8S3TVUYh82mGkIRTzEozcDwIZUyeKeVzrzulO3I31PS
xcS9C2fQFN4JLrUbflreVJS6uCwvCf5uTG4Ce1s3xndsVfKprAV5MvIM1FFNkopdb1zzjqE0ZPuj
Y1PnNtyb2JNWCHRbE53DFfrnYuTGJc4SpM43NWWiOXSgivg6BieM7igV0IcwSCXHUjfohgNRGDaG
d3SzeQ4aeTe4UgW+Oks+p2mS3bfbYu/x/K4UwVPaPUdvbDg8Rnil1/qbkJolmsiJ3gVxZG/N4Emv
qfNooceYaL5rnFbDtTzWj401ZUFynTkUMgiqamQQyZ8fMIGx47Sw5PssbVRjAHQCsebAo03BMSuF
0nRAzmNcbpX5cIki2Whasuv985A8lZ3Zb4hn7AGIxllI8ouA4tXzt06YVwDMDxNnph9oOqmt8Oa5
7JlayyJNKSltnioZFftxAmClLB2U9W/R9DgVio7Rj52ZAW8JlCPRg+tQ1bY1TA0RQeyQylsphGOk
scCnzsCjJZhaGdeUPKQLV9D8i0+z0vv9BrYROL39Qy7TbtsLrsPkPmhk0MBWtSiWQp5pzSBPbWMo
wWlGd0wvS2RzlIBunnsKv0Fs+JLyDIPTbND9fWpmnILWGR9bxz8h/WR31WPxNa8HddoAozGfyOXB
LfmvoJg9LSscs4yXCoBUCx2uO1qG+2eFKLq9OKkWudHxnfMHBi653v5J7xhoUrqRw73FgDRm1PXb
SoxIw1P2O9yEDszqAc3B/wMz9PhioOsoRLu4X5waN5VWKVzKKjP9FJ2w8MlhzDPbLSUEJW5X4FqA
1klU3punGKNg32JQsObBizMTVmPYcLxhi+jpEMnpa/mqCcGGDSnK3/wWdmuMvgPhsHVHiVnJsPC7
+xIIXsCzjDcc2EloQOzFFDthUDsv+OUs7FRZNUXQhjpzwR4YOjrOWJm883HcFccULreMzunASXao
YFQ2zgtQ41F7bgboRu/3Cht8flil0iNCIcKN5In4IDG3rL0qfp4agjWbPHC3mDk8dHOT9je8/n/2
oH1IpRTKbrpaIaX+AR1T+qxa3quJUJePHjhNN33GalvdFyG4JIzA56lj3B158PS6lbWjhJv/ETR5
QGXG4D/Fu0plBRC3at24QCEXQ4HB9w947HMqnoO/Uatu34EvvW/tHDLAKjZPZKdXhNVKXNvYZigS
ykRX5C1lN0ZAMYcAqGJ3ztfPJCdD2WM5KmI1yNJbUpnwzQfY7E+pphP/exea/ejXuWxVSzxFf4Kz
l294FJsN/A/PhOJKP+tQCQMuPVCDLBRjlQLe6uSyi0AXmIBlN2JPqgbf4XknLQJXlo0spqBdeWGw
9tGK8X4Kb4PMIRDk470+4T69NN2QWCqp8IT8dRQcPqvhu4TBnLgu7LuxOuCs7PW1BDNzA0RvzCZ5
wvZ5zpzCwmQ9HeyiKifx8HmgDQdeQlmQuhx62OcjWDpu5+ddMN3fd/Gmr9BdUmEMixiiE37aUdBq
Lo03btzAUZlZH1wEY942J6Pmreses1HQtjGbddwO71zg32BIVNzFtfxoQb2z4u7VBKbzfG1w6OYZ
z3ahalpmModETl4XsLVxU/30JCOWND3xzPK/DjGiUo3/T01MJcXjycVNKlS0ounlNhpKP+wNczWY
uEcGYxdnBQFntqfWpzXf58EIUJi2mkkWEhJe7N5R3fgXO2d9aQUEAcrXngsOEQSZNerXHskfaDF1
AnlgMVn2MUPqkGqtDfvuk0JV65iU9K6YNFOOoE1QAcvlu84rguN7q/LBAgiS3hhQAwdPtRTUA+Rt
4s6o+sk8zIaxONnu0nhMG3qV0xDIpKDgpJbEQ2DsvbxS+5OIZTkKr3QLQknVb0F2Bsgw/yKNAf4N
7/RmnIpQKtC26FCtCcHzQDK44j9uNeSQ5uaZhjN9M8Q9pbTa0TjUY1+D4zN0M5r99XeUA0Harp7H
og9+jIyaPA/cK2lKH4j/6StWzSb2/6E0SiMWx4KqqDVNwfdG5fEa9/P5Ncsl9czx4BlINDqm9pQ4
0LVx7KEh2d2UzIOov6h155T2049HLxFogE28sM3K6jN3AuLZXzRoPYe+sAQ27YqzGxEdDhNYDHhS
qoNy12taHgZdUHqFx21EOoDI8Okr6zxCrJoXgkNdaYRz/WpqLckgXnhoNsf4NVNuZgeaPXbPxmdm
VmAPdWsYo/hjDQW/3lJqv2+1Lh0XBHMGxXG7vB6WFOEJnWdpv12OjPr8Hvigis/yNDybQopz+zDe
14vaqejfj0pjT1G8mqPtB4YKAIW9Vhb83w+I2vq/Q36uW4hXJlw4leNnWzGlWUn86qvHIn4YgFzI
s0kjO96CKT6O1uupLxyIwYPfbJf8Dt1LVcmJz4OeMXLvKn+XevaWf1XQcQbQMIDsXHenKfDQeACD
DBGFQyWyT4ISvtAFXYMTnVSH+uUD4gSck1T97dGixxDsjxvcGiSDXn/plFc9UWFc35IDwwDy/wFN
7we5EuuODSiILA3L+7SIZfA9iUM2CVzyMGakHXXHF83Os9Bdt+b8wSsCi3vOgUXPYXu8MLOex6jy
RxrdP8WmF03fEm+KnPlS6CLP0xLLyi1p5fcpkSX/JS9KHal4RPkD8pU3ZADkDdIurwSLp5dQFmv0
5YN4jFSiBY/m3T+1cetacNcFpsaagC3MpKrowdNXBK9rgXRQnE1RxCyCzIBbMAMiFisFRLF3ipBv
M4dNkY449oJjzH2oPONHBVYL+BYDkFhKaG2tzp/rTQPu8zlKweeYAvegxd/xGlYxNy6fcOvnZ3Fb
ScPNWyuOG48LnaD54h68ri9p6jGdTVbim7PRQ5Xg2T5OtS+wfCEH4+A3mqaxJYDGkIgFzFuNQ3W7
0HlrtztKPPcWvtEwdQOWchqVcSGSLZmBQkKj+w8wXT980vR7/SIZzZPNYKBCTwTG961FKqGC4IUG
V1+a0haww4h0VTLnSTWwgkZtq9Y7etiOpFOqVRKiKQm49XGWGb+jbwwn882CBXd5HS4EWxCYNbAg
G9Wkg7ZsKSIQBulzaQCapeM6dXA4Yh20o90bjtSgVDKEo8B4ULPCJjXWA38zq2q9p716XaGMTPS4
1T0RwIr6Ay6GDc/60JC7WDJBizUEfq1MrHxQIp8mhawekuicuw4SrYnJoWtHU1TzmHJHHkNPJ4GI
wCAHntHGXtRAxTENW6TVOJJxRGTsGtOLw7vyYeS1dm3IrZ3FwEHVITCY1cOLLr7Pl4xZmDNucp7a
XFO75/k3L01wP2C5GE4YVitTgQIpAvIUYPIEWck6mhGtPRj39nmsb8mbf7BJHvNsAhd+jSS58xzu
oWR03UfZC+nYKBRx8mZvbCe36pNVEnUBcCU/3oFh+snxy6CfywavM4jg56Xk8rbVQy9AEQC/2Elq
ecpD7XbwTCcBJhdGvXTfaax4TK3iKOjUG2crJpPSHiPtGFb4whqiUebSbABMtso6teMpKyf0uxMQ
D5vUy6lbO6XpvqPh0IWyJtULN94WlIiJbeihBHInlEg28bw9APgTH86Ot1R9HqmZmLC8eqTV6yEu
0xHydb4aSzMLqwhsN1kxtRLOCSonTrdetubF7CuG73eJizXDNqljcX8jWLNHk4URpCB/YAapVZ26
dbHr7R0MnbJIN9pmeATW9cBWoXMJ8b3DdJydPU2sClJ9DaOny9nA5Wg1NZDcj1DTquYHZNNCvUE+
bjqt5wSM6z7YyKfu3bCIYTJEeozFvfcpp2h0S/yAk9GBdeUTB2ncAnwcxHrqbo9tMktlQ72LeWti
JslnjBZFPWTs9resTFr02E5lQq0/YI+SuIC/wB8GDcum8T8MfTb5m3ntjh6vOOBGXK1CXDXMEf3O
O8n6MER84V67jAW2eJCaSS3JTyywyTth6zkhG38T0N8adpSwt85v/DS8ixEWklDeIsyfjCeJ4/fw
KEkh7WefJPRvUJ20J5PMNpmh4rWXcxFoh45urnJXNoKCjZ2mo8eBbu8yWYTtm2+aWRcQvAJCB5Xw
XdurRAIkwzaZPFa9KLClKnI+72uLYsBPQZHUY5RXEXvkaFyZlIYrXqplaT8DK8G7z46xVPc9AF4u
Vy9PlA+M2SNPChqtpq1YFx+pSb7S7tuwnkYtc/sJ7FA40B7Qi5lyzsid3EMoWC6GQ0P7XUfVaMJA
wutzNLpf8x9H4exZ3++W76swg3n0qLzjkawegfncjpxoFewPZFto/k5vBI02qECLcTO50ECb96/y
HI/BLLGCf5GmbUlPL0Ih6efJyNMA0a4t2+gsOp9koVbbXn0Ba6UpocWrEJRtCSp+qZMmH1UWhiJq
yOciDINaxX9IonRIJpbaChCojaHYAEVNXGR3G0152x+hkSsmMdVoVxkVRzBwPsFNU2xPKK8eoCfV
xmfm4F5ici1e//gWus26XH8g3onhOclak4MT53BUPi9KhmlG6SKO7mFrpXjT2Nvn/jxAxtl4iWoj
XqR77ZILkQHfXFmSiV2hNc0DXvIYrMX89J78flObhVPDaU/1vHpk4/LM8NY1qlHShWzJ9+ZeUa57
pRfjR9ylTzLAcTDFwHh0hszU83IaFV4Z1LzhJ2VvyvSHkR6DbwVS7BeY5YJwfjOr22ciQWaRB/fv
9M1RmN/qIEbZA2+eO38iJ7nLT9c/rLPCfG6noi1zUjn63gx7hOBDQra+mKT+vX6251qekwOcUl7s
rozaOThUVjhgrgswByfBM60G1qeYqZZTyc6VH7Fydj1dgI80wyAxxlxHX3WAmo8yGKDlKoGO4H30
kv4U12zoIwYE4Mf68rO4B1soaFO63HxgDeoQB5aJGDRLZ1pLGDNVzf7D/asj1aGXcR3dd9ygMRQD
P+T3bz2YFlZTFmRLxk1rFkDuBW47MaV91chDzPWpGdERcXQbT8R7fd3l8vMqGSfF4uQqX3fkUrAF
B1Uzx0wIvuiyDV6wSKe+VLDScWBd6SSVBtSsonJnY9PtZNoBkWQ2QfbJLZFvVHz8FfodDjmAGDej
YhTIoORHZl9lEVQCkMTurZ/M3FEKDe0DpPJJkycAx3zsQl1Kwl9esuW+m8u6jdfZJ9RFXdWiO0tA
D+aggUg56OOdsToLI7Im9QMgF423MRAlFD1T8vaVwxUY0NWeYtFFokkLYzWnrIHc//7aJMEQ6e0+
B1SFnFuRengDk/e9XGxTwcZRGc3bnjVGz4PHQqnJZBb53KfD0fVI0Q6j2FjU+y1VnBvIbpyZUuzj
rTU6bTSvv5n5/FI5yZL7y0A69KwFUivauo3tJ3OvBOwsHT30zrZw2IZS9Ppy3sYIXvPrSu2zXjBb
Jk8G3xQ0LjjKdyFRLS7akuOGeCD80oZmC4bjw0gy1DFpn6Nl8V8vTMjdmyPOlaRbiu1m9OKFXu5p
0AE+d+XUauycmYLoYZ32r39VOxwF20EMbSb4U+SKHFA5zWniip1AtKQDj4zOOn+NZYAHkvvjrWP9
ksdywnCaey5Qi7Zfb6prGGoQAW81q4pI7AEP7AXYAjL/uuDisQbtSCe9S+29dyB6xImvJvDqu7vD
Wx1iF+/07GA+RihSWXQkFhatNKAHJzwoo9vEOPq3ysfmckH8y0UaPwtZAReoDTelBZrn38fviltS
TSnE8hycq8Q22vu6ElzlFcq8jd4TYrWWtnEg8sRm8Uu3bNNOyrH/pD2gm7SO170omyf1GbMMOslX
YeOXiNv95X6Vd6sDPfbpymbxdlMjFLKh0vYI/mAKOLdrv6OXY3PHirFacO/mUkx2f1pX8Da9CX7d
Lr8+CT3NClY+gHx2LpXxm/dmRQLd+04K1K/ZjnVVwbwaZchn/A6A9C0EzV7MPTM3eyX+9oRKVFCw
p06jGXe4AloyyW/nBFiBb1I5MKpEdTbBzVoTHpIWgxMbJZq/0jNCrcK62gpwKQGfDn01r93yvda9
4hyKtECyWKoRSYeG+dvTt9Shc9+5A5e4Zs/c8N92p9aZ3ou4Rr+M9eL/hu6hDB7slfrZFSjvP2U/
poeISCClKb8Z1VRMjbz7NGsXgbD0NNcQcVOFyzfz9aEW1jAWsiu9pUugnfX/rJrwVAEHpOsaXf86
U8qus2hlRfdOBKFhv11w/WkoQaoIAlZ3qG+WV+ColDYBs6f90Ku4EYxeghqQtmC42Fj0z2uC2ZK/
Nkfbo9OdbakAU2xSYRBy7i6D9g17Tco2lI1ZFN7Xn4YetKmfZYBdoak0rycpifMkne/FGGseA1uW
h/asXJppahAzHM9OiAIeTxbRPO/sxDN85wNfPL3T7TDwWMeWkcU/vcLMjBaSpL3emtOoODL8+p9T
zQ134sqsC68nMdjbCR5bAZWjNTKWphlkNcG65ZzE7WAVmpb90NNbBV2zdRClhxeA8gszK8utLEeR
BP9jNszUBRPuGmlSRPP0Ti2hp5G0JjX4/brY2q7OAAZPxFjbk2JxWDvRmESPg6WD6eUAckzB0Wct
NqprATgNkfth5mSyykvUHmSwkFeaeG0llvSFZxSrW9oDu19OYg3Lx7U7I0ThP+5Owr3SW2Oc4eiw
2yjbInjF4o/zePEhf4tzpino9ceq7quCtHw2yMpdY8tVUW/vMVKwJdb/ZNsOCEI4EbQzyR31iThN
mACD03E1SOde3I319Lov5VWh4eL48dhiElHPK0Wx4LQT4VYEkW4IC6gLNZLNGTIaFSGTXV80J8XL
z4TOpt1eXQjRmGj23RQsWUvyxijiFgW9OFggAKokKmMzUUu+/MS/V0knoSEVc/cN2ata0qpZK3/f
QxjuLyMGtJmipWvXXOm6jL+zgPF2J75TG2aqY/MSJgKu4H2g8blqWhTgFI5GZbH+eYIz/tQDro4w
VnDrWKlT4IiL4GDHIfmMlYmLTG2QI8V+xafEsO7MDbegPgA8OD3/U6r0dq1xoY1zPf/HwJmS4YMe
+ZRUE4UAwNrqBSaSTUXA29Jq/uBMp0pZea0/IGz0qslb9eLHnlvGopsZPv6ONZYDiqXWAAj8mBIf
MBS+f2Fq+aXCwSXZOrvHr+4TNc/pbGHCzsTld5cJmOFs/vYKOPA/iHIV7r4HhBodb55nlov8z8+M
To0LqOYZKoNjFY5G61W5hB44EpPSSt6r2BTW7d6ZSHywKCmbVfPsSYmOQAz+LDPNXlFbOyAXFyNi
30mFoBtGPBL8LVUQnF3495S96lKTN3BwmXYhK90EH2Jouf5rHXXvNj4UU7IonnyYMSiS6tMPFE/B
fCEn8u0nhWK3Lc8/k5rkbD4IZyC102H5zsBBlb8VjSnma2EtXsw7P/TFInHYntUaLCFGrBW5lqFx
AIvnSQ4cXtzqjCCcRfWmw+BrHmYEEHLXuZTfANX222EWWrSEx7Jh/oQnFXyi6dNdoruEuoMQdlo8
QhCQO24rr524pdJ46RNJTWp876/B3Q9vfy9/sgXaSMNmG5JCzahQRxKVUydc9oglEbjii1Sx8VR0
gX1Xp8BFCc70hYmebyTU6DVMcVcl/kMjk5fPWN8WbDvP7ceW1QSbW7548W6rcSDfglVu+WXIfoqb
qv+4roA4Cmre+GRqaOw0qHm8Xbc85sU237Jddvvgc8Aa5scopEf2McFFriHidagP0+ZkxJoAvvVv
okL/YN09/7kxaq/7mRpkbFNJtdCyJYimmBsgQ+DMLEvTs/6L+VbZXnz7uebUWpbkeql9Yi2kjYyi
KSn8s9fakkDbn9se40uWToy/bdQ7V6gW2Wykz+WZpISGp2PGdGxxfE51kCWA8Y0PPtA8PmeUbsrU
cYAvJGKp/ixCY7rzEu7vw+ON9vVPrJ2EZVhHJkSGDlPkwAstmgxS0r9zVrT7w3Z85rTBe1pa5Ldp
lrSG6pEAHBF2JukpQC/iE+ZbRfO06pk9vnSsC7jyHFDS8SyRmp1ebtMwYXrISahO+zkzpp2DT1Wy
rN+OUWZNoyqq7SyB/QfqkG125Q+L9/x8zQVz5zK/R9UADAlWA9RNQ55Z0T/IXyGG4HmtXbozoFng
mw1bnDzpR5c5fUvsLiZ+nr52t4/mT+vGD4ly4/dfV8kiZAOx7Zoz7xK8Rjy1pfh1lClQHrm2k8QQ
2JTS/tGPPK5QvtHdRQrpPIX7juCXj20pCyL256qVzltRiBCf11smG8HEBVhg4rndQASJ8T4TkcTS
9b+KoKi5S+Q6QgklHi2ITnukgAmSyF+9kfJC2u04CRkE4G8UAr248HOmLN7je7bjt9crBzmgdGuK
yM9z24Q0GBgB51ehfn2mFYib13smUdXW4+ml36roOLnCKroh1r8LtVCCMSB/ljVcX/G38cISOPIV
+yVm30LFVXAtqEdHKhW5YMcMoJvwPYk7pI1Li4I/XLisDCUvS+INbJi1ntqTZsZb+bZqp5tWHQTM
d4MBsX5kFUefJ/jKo6Mu+xEPdnRoKZteUBjDhWBnCAC83un1aP8XcGmZXYHS09He/GKz4zIOBMmS
bu4v7YRTVq77CvA4OjP/TAwTTLLD9NFb14DdZ5lbRnESoEErRJlkK196Qu0cL5kPBBMClDTAPD73
aBcjGAeOLvjvwD/wJkO1wy0XZ5HRDLNd9Ts9kAHCIrP9yG4CsvCrWdnLwzGQn44mqiAhBDmJh+q+
I8N6Kk9owuMkCkzUuHW1548tmFpiBx+QNwAFykg2n5vvs3nlTw+XFvOa1HniV3QTtlSIHXKcEOZk
venzWBaa1hm3l07dYisRS+d8ktA9toZlAq7CdBGGj6bwI+VMllrI3lv0Sb4VkwuxI3c+ZZJlVVbE
KNLIO9+iPepV6GFw2ZwjjH1QKwS7JwfPcAGVhKP4dkVkGMSYseBJ6AX5BmD9yGxUxezMw5JZqSw6
WD8ceu27Mn7d2ii2PvJ0hOc4VE0trBLWRicGSgr3Dq4325VdGjR62UMKy4y03brMmw0iiYaX9v8S
jDdJWjKUe22CxAS123Q0prlMV3N0O+htw7jogzC3IBEcaRzlph/i+L6ZOFmLkbP6ksRaO65TEyMD
J2/u73wf4bGtrrQU/wcWY/W+rd6EF/2En+aD/zRTvOJittdWVS546jMPQW4/3F2o5s1IpxYS2fk1
1j96mYUgW2GmOUFNgcSCGJfwMcZyRjxZNgZwx+BOYhZcyo8jhCNl7gNmJKa3p7/RXuYlcvEBBe2B
sGfXmqPdlLx1k0YqNhRbpJ6T2L98v3aSNImeJ7hJ4Da8uhL2hCpMo4XaZUfAAwrgWxqe+Oribt70
AVnQ3SZk69WN9mYb3cmdXFfVEKLY2C/MWxBu0zLvAhnwyA2RO/gumiNmZhnakDS67gIrx7FsTbWn
pRBM+9vRjSV3zA0CjaPHwTl42bqWBblKDa4vlilRWeO6YHzpUObtcZxSb7jM67+9K8WTouJI0uFA
Nmqn8NLbMbvPk3aDrosSrlENltP9ABUbJqo+E4Q/CnBFvRlzUvKmJuhnk3uq6oRmvcyIMoFbIWoX
U1UDK2CQhFmXAhZZNaiEnwveVE3WhwHiF2IjU4trmDwWh77zLpiIZGKR1C8El77X6twSsW/GVqcm
ZyRCC5uEnepj8KwjlD79rAyis5a+E4NsqiQN14dIogHuGJQAX9/9lddIX0qO4agvzg+34j/Jy7Oz
tAVllHTpzG2Z3Dk3WBRf4+pTF/8Jphuqta0yLESCksIRRkb6VQPZmt3uM16N54zXUbSXXf4nq5Ld
jYjUvq4RWivvrJ+DouAt0kfh3EMNnTxFcf40mSSuIVpnWyr+dAw2CdurNmKQLnXWaq/RHeW5Fs84
zB0OvztH1CWUEY9QRXopQUCF6xoSL/nbdCk7ARNcN/PgwpnSfXAH7BTF1MzFAyR/BsA2EtD9G4Jm
IM7i2m6I02JWi4VzV140bYtxmT90z5pF2mz1mR45ZjTw8BxJQkK56xYklTrWobjkfkPOzRqE7dYQ
Bhqii+GB4ndhgnyN5ja1FkCmSm8+DDhZyCgRgnMvZVt6FDMA5I0WYLMP2EWIDxAIzrixlMYWcHMP
ttE7+nn7CTbZjFuVBmygMRX30mQacbMtxKK5IS3sgoVdbRwojJFULCdh7JNQn5BmAfHexC60qaaT
SPwZKSIXIqO/Va47FtigoWeKcOA1QHAkdWKwW+pUURMCpiATTmdSOxpe2unbbqeR1pqW1QuCiju4
7yJm1t9kUitqpIfq+ZLVj7a2m9UXnI7Rl19wbwJGmD6qRHWJUsJNelZqeUWDkVoqeFAjUreQkVMJ
2M3503riBnZOdiz2MgGoioLPw8fnUts6L82TECtJc9Sq4AjZHWTefMHh7j6xlYPzFLx4KwFSqYTd
O4fdOyI1tYy3tcmO3B3UmJiSAPTZSNvHqlIuIRsAxrPUhv5XYHSuWcA1p6ITPDS0zZqU3Ifrnc0h
fNgajN5sp8cxdNWL+5X+5qnN0goYpsTZuNbaNXPCD4VFlaIOWkjivb0XHHuRURwNmNM4m4BFPSRo
TLZjTGm+o8NdJFBPf6kIFbRukn/mnMhqM4MMjGG66HHEMZjpvRePtaASXtZ0rKxxpisp71hUTu3b
6EhxnYskqOloaiGq4H1NuvQ4zUUXFHSVH0K1rI+w1Mht8qR8kYvsDepvbvz1x2CGT37fmW6oDOmt
dn/fRU5g4CiV8bhRTHYVP2gSnrlWuTkKKDKe7i1UgJP+kWINx/JqhKIS274v8cVRXd79ZCW77MVa
z9yXVSVQXNPG82FOn0QgXcAoMhULpnKOVktlarYqehPmxYV9+kk3q1GxNHPKPR9eCgWPRJHGSBB0
Ijt5zubZx3MKiZxxPtWPNWKAoTzlIOGwQGrfFDKPvWiQMFw42FITRLj28DZ8WPhBHzzA6kmfUmxY
GYLMb1sGxXWrhI0OBBITvQlVlHYGvDKK4YreC8qoLUXTRulGLAeZhAwKUyRjjMPqaJUMwxTwYZNo
3mKr1iiF/Ad/mbAXpl9FAQmFcQI6gnZhm7ouEBbKLNxFw/fIWGqYciYo0fTPP07enLK+hZUY2LhR
u8CUNWRNWjYKK1Z1YyNLa/dJtKf8d69u2jbVZtJ4mF96BRZL1tjhbyyG7kSmtby+EUuR7EJAdyk6
E6exqMsdu2G6d7kFIYWJReHD7hgcH0ny1IIU0dZaV91FsbTO5qlesqcmTvapq87DkhUfVGJG64ln
DvMr6jTOXkWVJp7/8MCnO/IKZt/eHPcbLmLNIfgYAlIG3NKfv0BReFTfFaql39wb7q1z038LVO2w
VaEjLw2D0HrPjgdevVj8C0ycG7CGIjHl3SktcKlD80QYiOYwqMfiayj2i9Tmf6onWnxsvNxVELoS
x30zmIlT/QrZLXS3RFpBHOH+IbTj++dhZcT9a28T4EVHBFtzrkxgjCrGQkgsYlP6+o192S+luzSF
IZCdoXlwM6OMRforKTWUZ/C5RcWIU0i37fDk/KHweftmCHZLDbukFQOEZPjSDKdoAamsH2mvkncc
u8J3G+I2cJc9gGAauyVDSO2i8iUpi0xrXQPI9Eq8ag8Cc4R7Ra8rP6LUBCiiYKTl/D4a/OxU9F0u
IGZqh/49fxCoy3/9SBknH8szK4yB/QpXdbU/bKu0uC21llniEV0PBmlsPg/7vJxcvilBh4oMyQwC
rsOUU7vb9d6JrznPePun4buMz8iX6OBBXOLCjYLKUqEZZfVjzORWJy8U3fMLU1ndej8oIYo6j/5b
3C8qX/rJFpicGgZzRymjFVA8AgIeW8AzhuMWql9oJiIgNW9dJUzQ7OdLLKr5Netyay0vJ80qR95w
H5R/axmEM4VHkSFA9V2SMZtLFhfi/ox8NmOMNG14gGO1+5HtfHaHfeAgbLA+h6Yk4u9jYmcSeDkc
+fIh09AHRITIIgIva2/D5cYx4xGLyOaKMP++w74PQv7v+bEvOxMkvSgQdhtuw0uLuEgpgelbFjiv
hehzKEQefS+5PxF7w0qRcb44pN+ebwZOHz5tTUtmaTcEzz06Rg/u62qqrLEL8VGcYezsDRJKUjwm
qREbCfu1NBq9nMVZOhZ6Qc6/TISVYjdpO/YQXfO2fHeh+0z+nPhDmn5NJMhBGOT6DqrR+aeammOU
QpBm77nmvOaNPWrsl3+A8VvUrMd4dINavp7QlPIITyORP5INWPqL3/EdcX05AJydEZW5SjPQl/lb
bnQ2ETHvomJI9Y+SrZOb5uhQB7SZNX63ZtkKjgqlPlCDjgHY0YzK10FVPdPc3N6z6JHEE4iUZZp9
TjgUcvA8Y0ox2SeaxSOLE28kxg4JqxS0tX1Q8H1Ty6DFNBza7Hut5YR3Sf1kFFLfllwFFpBqXYBs
jqzbutdctV/x3N6ehkRK41YGM2fTViGm9T0XvAv41HHgQKsN8lQUPgyHpNLcpj6u0YTJEhdib9y3
F6nx/JKg1gR5YCOA01AcvO/dxqOLhYlFtslDtXTX2VVKxNav+I+m4+XU8Dc/2FFFoW1YZZ/5CQgI
w+zzZF6YhESpdFDfeRVvNL2wvPULPi4gGU2Ve39FOF5BqftXA/25LqY9UjP/Gt/Sm7U9j1OYIR/4
R8QgjE1mltJMlwKhh3BFTXce44r74uaOiHaotSWkF0ZMAZgHA17JTsHgZPknQ6H4lJSnvaa/OOxe
EXMJH0qXFG9lBR7Ph0FvlK0OpkcZ/Qu1ivI3isTV3lJwCQmejGQR64c2cjqMrLw3uDxk3X+4Irr1
/Qt5yqHR4Fe8gZu7/5pzmOksjwWWAlCTmwqqFiWHzsgg/O2JJxXxiQCsm46Ze6+q6ierC5iz2M3E
ft6iUqGmNAIvf7MFSVelr12B1216v1z2M7wrLK0xi6A2KyZ52rV/yllsA+VEIFxlk/bMrPiruQ4w
Ptcj9oZFQ/DPqq7dF+7H2YHJFGY4sim+wa6FoOrXMnJr/+8PhXzqh1wjJkT3iKQrGhup/mBTvFxQ
glaCYKYQF+4Ep81VUjaeDursJA3OHoPtEtBcGCCeouaNoqTy3vE69/FIwcGXLrY1XKjwJHax0xXb
7oYKfCiNmYsd0/jzG5CqmlJtmm4NEpUfeRFIFKA56HrBg8zLp40k8ev5qeUoML29tyehEnmj7PpL
ydbX1fux5pbP7UUTQj0quA2MQRvWYABgCmCqcUEbjj0Ei1UHEvAY120Ce3Sd792wl7WMK5sY69SC
d3ItIA2nNIFvbuovEFXXWJk3bC1y7bZ7P8k30on7ZTFNpSjY/UfOWP56RMYbgTRJJchxLtrxZigs
4EdbhIt1BmC7jBWCKMCcC+K2IdBaZ3Z29T5+lglD+w/4wkRzU3iPvmLugKr7WJ2Z6UJvejCv0BqQ
YsRpnzbbMvsBTyo+FufR6Wux+TYKLSxnRDi/lWxlEkJsEZRWiD84agYlidVSnvvLE/PF6JiHJoUQ
TjEsKWsLsD5XobEwBBdaZfYDRp/gSJbp7R1qm4choMMiDmza588OuphrhgzMBRAoYG7xwCBlJb9H
kQnLHkIJriJHpLxNcLqtRnaltovQ1pI56rjsS7ilEDwo52Isu1vUeZGXcmmogGZWD5lH8m8pB49T
5OJhaOyDgBEOeRKextScdH4a67GeC01kjs9SZptfvrSsWvgGlr3IsyT34z44B+SbkB2DmxQ65u7/
xFy0udNZu1RO+plR/N+LKUWoqXY0qM3Gs3kcsxtPymWGKOURbD/hLka0pI69ZZxbLIlr1M5YcV/K
sjoD4qThx9NXXHEWvJnOIr5IJvICIFkMt8gW++/HTa+yT++KWhFR0mt+6lwdXDLeuNdAjcAmhQKY
IlHbCPidX+wW6Aer73OAKZGsGayIwWZxoThAh7UZNUEbiHtCEWeLIGKZlMrLLy13U3P9Llfw2O0h
MqyIkfkp4YcM3N7QPN7azf/5QTSO8rEgvrc7U881BvSdO/5htdtIwns9yRuGCl036UG3+PkhaNEk
RijIEkNgErMggCSPfAD3sy9KTNNHVSiMkwfViq6IORCvy6ViK1eRpYL7Au2gA7Uptd+7ykklTr6G
jvrZYqhPz2cvTi+uqKspUcxDtRTuiOlxaIkfKRDXcQbTqfS0JEUSCyw1P2iO3VsaNOax6i4d9hKn
LAfxPhAYtyke28Y01gL1XvKaw9h+5VrnaBO+pzezF2ehgckQolZtXPPs0dyAmygnDg7CUVIb9y2j
ouNqPu0xkUKB6DoKuFSYt1B9NfUWKkmrn3R8RAZpiZJenyjhyq5DzuTZTo16sXzRFDJFG/Zjepxr
E0OOFJI5ZJrILTuFBkCComfemcxdMxEt/OPtSMWzhYx+9fM2My5pK4tp/c62YLfNlINP75cwo/s4
D9DJn5m9ea3XBLGXjdNQ6lWEjEY9nglrBjenD5JwsxomsoFLroAu919nSBYNOEfdbsKhCxBuinz7
HDvS7wrVZb5qLjGagHgbr7oD5buapu93fXSHgHG1YAFmdnYGM7rBqWCKUEqwtC/4YzRZ4KwswwVZ
irSx4NDR0G14VwREEYFg3QPd/oHm8VIxMxwsb6Ks/QdaOZmmdtv5gclagHGIN8MYLB98NFVqkQbJ
YWER8H/fX5ASS6yFuw8zBSekpsddi8k+LhaTwQ8lVi/XYMFXigJgRbt4TlIsnOmmmE89DaMwpZak
LA4NjL4i9NbBTyx6Ylvo6CVi8hejL+vwuEjw/AL+1Qo16qSUYZsMQajSfXkRfr/m0oJHAhO6RN73
l860UCUB0nS77d/EGn2WN7YrQIUZ+24dP4yot0qWRwOtb+Kl2UDksaQVouaEt9HKsx+2pcp+SOTz
fcpifSHQhqrCt0WBAdDMUB86Xunw9OjkNbaVlQUnNx5nn3MV5Ybus97FVj9pe2UwUHx2pYqO5YRK
GKSEi8JJdCjR8thNzHX6EyDSATU8UygmGV2RPid1MFj+0fllP5SVJ7cUbOsoTpVz+LO/R54WscF9
4qbzd0Zijng3em0YDDwrODwTTmunFy+BK5P4OdDGSdYDPXKoHonNcGpS35ef73ILbmuQOE3Q61HL
02BBYzcopZH3UUP9WLayeGm42QQLsBoLeBjeZ3dJ9NVssvF8rWAwVRI0k33Roh/QfrjXPuGVmf6C
oOgtoFnAOHdUtkMvPxGlKyQlPenBPV3xLafNksA/pXxqa9eqjg8c4DDYZSAUW5DatkDLEDWIbs/7
MgjDqbLtsnf1/GeAIbeClRGRKPL9Gnx6aWfn04/i4EjHZey6oDNNJX6+SewfZYyD+RKbshr6KnSr
XK+AAYJYkvOMsnUgLz3rd8Y+zZDORIIwLRYune4lQGZ2m7TxA9ZAAkE/81viXlCp5sNk8Ix3J9Sj
+jmkKryKzQzYw7+f0qd0qId+1E/IUjHDCuY+3eAMgXM/CAYvMBxxV4TxurNdOD+BMSR0lVwMUicf
V/9zSVRGUT5wN14Daj23ulwSKwKkPRBg/Esw3KPlJYkQBIPCjl9pqqLb2MO4/KLdvQyqcwTdo+9m
UKrht+IZbtLrVqdsJ0wNDbLTGEpeHDjvRWbG0mmMpRwq6IljAp8mUxxYPZtHBVkmwk4yn2gZoaMZ
DYWsUpPEr7mzSgECweinmPgEgWmZUFqslMd3DQSOEkScP4fCZV/1pWOtQSrUjy21kVEKd1pyV3Mh
mZ2drOxe0f20D1efmTaRCSDbQtNxlAXhNMOQOmBKmjoHZEmDFdZ52FzlzJhTU2l9Oo6M3qqWd8xP
RkKCTwFu8/xavqgHIVlZg6vSZQ3YIzEvsDXZbJSsFrmLJ+ja+jibcHN+8hTmFLAtdajePY4DEdeK
ZER+W5qyoCTdOD+uvWPdpuZ6GxJ2jTtKEufJI6ryTec4oRECez5/cboXPLbBFbcxnDKITc1z6FRj
bj2dtlEiK21YCFn0eic+w+6nXmkr3PC8JKC3Twt7dpgip4XbJIojIQ07F7Wkz9hM5RLmCX/ggHGB
ktv7izem4lYdH8WMXiQ8y8eRnG8FrRophWyII3VwZDwEIfy9xvYv6wKx0aZGQyCTN50NVPPgVAnV
Asxr/gKr1JR0kfmHX5csuNdV5v4DBDsI0U9/aGVllwc/006N09gTW6ZUoiICrt8FwvrbSCMfVxwv
OCitRO4JVnNSdwuW+iqTJJ8uyvGovqjOkFcakQP6YpZzUTWyTiprQ+/MHC5p27aMZ6msBlfYcExi
vAglPCCyeO2atquvI4svN02vL3DYfuEX5nHB7PxwirJdqIKyC30WnYkt/r6OThF3F2C9fc6SMFnT
WwI/JG0L0HEu5knlPpYG19otefUMOsRpUp/4KrcjqoeqGAxEWS8VJljANzpA+4+qeay10HxMWziI
MjH9sgKM4YlBap4xdgmbfRdVs6l7NwWaupjJ87kc1ZpxF9Gfph2QgKu/vdohH74Y+FgDazC3xSgl
QZa7uWdZKKBD6Z+ZbajCOuihzDH3sUlhKCNFVz1rl/sFnCAMaLWmm+eCOxesSIwuPRl0VzWl1n0H
H3i53frNX0ISwt6/GujkVIAshSL7YccjRqUKDAdwQcQ+yi6W1LwguQB0cQU9a98KJlR6xuNuM0Vc
ITCxDk6SjodWGT9iJsMhWzYzY5snbig5ThiLLTpGKZdn2VRcOKKYCC3DjU6puVV7nB7Z0BIAQgRF
VlPpoB/EKubBu80Y8nAPv5X8AHM3L4hUrE1ljkIPM/s7pc0P4d+s0xC23dRDaY9SC1OcC5/f7gtX
kEruwYY5yc8ec/6c2aPi/duF/eQ8tQqgs9fQvnCDJ/Zxm5vsoaUyAPQd6ekWx+U33HFmWC5BEdPt
23YRyCzW0kmJEBWgesupVTRwDIQlwbAxP2s/jDIVuIDA2fhVFIgGiHq5OByaDi2lUDtQnHeY1/mp
YRXGBOKTnukAO66NP9kZ/K4s7ynOKi6iqO1PnU9XnJxXU7hLuNlX9eHA9lF8hlOYK/rLK/4fn5nQ
hTGmUM3h5V0YEX9Glqf5zZ8slj7wIiswDe0oWfOg3qRl2nozTZAl4aOer1+RAg/XhF2LFPMBpJQA
0bN27QVT3WlAamXweKq75ixUcmhMzAI6wRBClGOkrnVpQwhNd7f3aDOTpOyCcaPCOeBbumVjllRB
KnlxQgMK2ruPNGhJg3R/i2gkm5HTYC8ybQPIgh7yboWTf5epR7BarNhlYkJeh+RWSzfCjMOC3FHD
nHAVhrwTbrA2Xq5t/pG4zVlekP1nkImxEtTeGp4uKBj98UfYgxIO/xW46ppBy43Qli62ptN7Pqiz
dUZHVZrEFrRB0XIjvRUo4GQBbqpwofNaO2Vt8kGr1RI3rkprfSd0kgUMRroagjDwq8c4G5tcxv1X
gDYuL9acTV03U03jj9SggdcNoBAg4OVYnee246KfJkIJ4bl/EUuiGnGPswAjO8dp77U+fbHha+xE
UoUCh5iI7XfH7vmskarDoC0LRmjJetlojUIoG7T05AWC4L2x3oN/RYmgN7iAg9Av/Ym0Z0Gh6IEq
8S81gFqUl10a7TvyX5Y1AAL7kqoRTj5I3gRv/oqozWLuZ6NdUw4Q9wdvrmP5Oqzh+SRc8tw2Ry/n
lIPm88FFSuZN1IGDwMSL1b+4/IaNAnvCqnF+XZ50IUeoXnXWsd24SwA3aqwjUkQIe/Ena7JyvMVu
Ik1S3R5cN3VNcQnN0TkSh9v2nDAlllL7Fj5ziT837dxqKfNo8SIcmXrf+jxLAaumz4Vxza8UOhvj
XPhiv1hqSukg+ys9mxa2vPb2bVpoBqkk+kh6gwQCZNZbn7ILgf6WvviezWq90a31cCaCS8PIxuJ0
K0bdCnE9XNh221iBe7hgxQUY+yVH7RHhs8D4GwD5pINX00ngkl9bVp4fxpxLWun0m83FXYuBb+yg
5wo91DBCaFlQAoL2/ptfpj3/sKw24qJKjFR5QEhkkvPhXZ2gFPK+oo50t12Mt42RaBOMHf7UbbFp
yAXTxUBNmwBFzMyNRRkrQWN07bSg4Cc0/ihSUJc7DZn3Wd3wq+kxeGsFW60xsSph/5JNLHzL8Y86
zf4wt8ncH5RrssuwIWZ/WOhHFz4GS0AYj1rq5IGPQoB4yfsx7NrOPcfFcMkC5ZlCj3yzQ4747qx4
8Xs7BgNrKOB2AeKQZokcVcFvzRkRt39IAhuBJaOECC2jGgExBmcnpyvakvjmtqmRXqwnWvT9tGY/
7Bi0hRwXyxoruxiGNcMI6JiNQkk+YIr7+apviXk3asmbTpMrpzb9Q9AWby/IUcNBdoLoWV7CtkRE
4Fx2LumUNnvw1WmH6vPGZTTxAdX4ZyiuQ8KQRSO0Me9r8a9gxCX29aOGAIUY5rg+crGeIS4BU761
YC//fopN4fT6i7Z9qSlgvfyIb6kapSJ8dIVoEpYbwj9IRIlCFDpQBAMd4toCDGwABQsnrA2FLKUQ
wE0TRTPsjkSSuWeQrjh3y32we3of0sHXsmFW88AhSwyRBRPmCjnKD+rgwbvcRbRWsy0pewqgm0wG
WPU830qWu9jbBJigUEnfbEQpXdoP/OY+cbyOmM9ZwGvMhZMVnyPzflaeiABpJiEK5oMgyyZRTElb
xDKFNeVzl4wrqD3lMA76tJMzSIt/CM3nqxnDURXKeXrCcX+3PguAMjpXomr3j8Dq3jZTFfdgypYx
BddjUojdwhNpds91YixWGbcYRU3xiYx+XLbiPtlVlfmwHKEh9crqciAgqc8ue7pk1/JOiW5HKejy
AwQr870zkaXKY8jlBI/+P3lnUYMGcvZu+hvnnhURgbD5Sb6ys+lm97ugPOoAEMrrNNQzpyDLEouP
W93Mkes+evWIspIyK2Zl18UVT1yRRvgLEyz7IbznRrysuvz9kiJY1LshVW8J1dHoaP9u+LqBxQzy
+Uw6PBOHYigPFT7GzLYZ+5M97sg7HsvmHylQL0lXUxTmiv0VUga1us0AVJ2DbPDBdLzs85eyp4pX
GiSNg/sGklrSc5B85ew/l0CZ83dt245pe4ZBIAbY7lRMurem6F/SHxMsn1p3UtPCJSTFetDeoJN6
cN/ZlrayfX9jRCB6ZoWP72PBattw9N+aAdfEz8fNr2OPg2SLfilN2yOrbgOOFc8teUMDja2U2TTq
AsLU3r0vQ2azA9UsuuzXbywukoV7mCegIbVxMgBAbcauF5L3NFzy57ld+xVmFswhosDOGWQJYAId
Msdh5GtE7sIFJNyOYGBugV0AhdMySLFGrx7A2x7GCF97Q22DNl8wUfOZCmttNICFImebjwuPLa/U
BoroQXkCbihgd2juR8l74Iz1/0XyL5xzDErW+QXM/DHXgHQ7xljgBpYOHDfBM/LzLGTwsaxEE+TK
FE550hDl7TBHKpSeGjPzokDo0LxwGLUoSGsxLevQ0B2DKdefGvc1wkFttSV2QUa/7gUAzbGByUdi
C1YAYotqfcIxub+hfhdj2eyAv5xEF78sUnkaElV9F+kTejqA0RmIg1O6pCoygEGteAAKj8k18iq2
qQ40Eykv5HjtLcDMVVLsMCdAUdhdjza7oRHfqMvjRnat84yOK+fzeT910IiDLelP58TtvlSNlHqB
2V65ak95goTQ0RIVuYnpzu1HsNfCfZzeXeGj5mL217bDdHWIVrH2AbPHw3AD/H+PaAFd3KlGANs6
ca8qFNYfMkNb9sjUIhK9uHSOXSYvxi3qUM6pCE//QPhbTxNQu5liUwp4y4+xXDeUTriZqaoUJhKl
1ex1OL27W9RRZGCt5sh5VnJPcdgGD9MiF/lgbR2IpRB3FK3tOalX2Xak9tU5hHGhxqNTkTnyPh8Q
zGXMzzJilG/GaxDFLqtKdaBXFCzehILp/d321pdgDBcKd+uhm4kDsxscCZ0uqKyUleYbN2twIW+p
Tb4Uo20LPZ08pqnXSxCMlmLdcmrvY5S5rq+ITuv4+3pKhlE0obSiR/x8GfnsVQG4MCx8rdK/WCMu
HXJIODWziBKPt/X0cgIqKqWZbaXyp+kV4l/hunI9lbxD2mSs6iZvFI3ONtN1I3Z4TeuSmCean65b
QbMZXFXenllWQLKOiidFH4PGJ8be4S1+E/CgnwfvXqbnAN3rBqhk0SXIcRo0FY6obVVIa3wDfEop
N/0N1a6w992w0AcobxyA5CIDHHqCtTsydJGfjV85+lbFsAcOqR+DAPfnetUtKGrJZ4Us7aszPOYi
SGPDJHrrBbvcNviTGzy19TPM01MDt02kESrxm7Jt0Q0OkO4MP9QBFkqqSC3deK6JCWKWvKu3NcK4
Qr+Wy7BlsYUgm/lpnzBzg6QNyAs5cgoUxHNz1ZF1F7kBBFMUs3pPzriWEHPnBmaCPij/he//CqvC
TJxnCJomYJfurL4WXtKdBakROtiQ5+BDgff9gUCzwbeMubkpeonj4SlYzDlQQsGKEhxQVeqWo5wZ
mgV7s6aYZOgVhz8MxxFtbBscti/Zhq/cdzH+9V+/PakjkWsGkM83l842wy9Vtg0affaNT2waU+on
edjFWebNkS3e4Vq1kCa9xfhFeiNzpJWnoGmJEPN9Z9rMilMC8/kQxz47scaYPLPylPTxUuhxL25B
MLMWc4M4UI87/q7OV+HEbFOs91gV4DKaT8Ov60Mvdc0PGrn/BC1aU+yO+aefWe5kYva27w0xRxjw
2UcCAHd7DvkIG5J+1IIcRvPJn/ti9sC2xd6fLaUHjIb4zJqgcpVczOCPpNnBhw1GAHxF8JZSSNnA
PXftZK+gPOkA1ZifcjADTfrlrmeN4/wecq2HFXYIHCeXRyWXtTzWfkIkkqXciT5QjJOI1stwzDvt
3XGTXhtCi6wZZ4lGqqxiRWprJg+oaKfGf2PZVmoz60zSyRZU0s4HUbjWm48In9bERySXY8DxAZZM
WhdtN6TQZbyLe6Q3xNexXwFXyNa8n78Rm/Dzw/USfEcfdjQxwr40ldH9RvXXnlANUH2VRBjUMZdT
fEKv5GV4A3s523MER9D4hpNyJK3gMwSu4Rv+xyhyBHbWlGrX0OhHe0XccY27tXNsgXIMnG8DE7d9
dduknMbG+MA2GIHD5rRPbb8jyQ3yShbMYjr7isekcq0SQEsOJ/02KIzrWSTRJRP8ypaRMe31Magj
8j8ahhRhcq4w4q2hcCN2IBIVdLTXM8sOuR7EP6U7kzMh9pcRooXuYhMLLUbjMGqA5ug6U1zRkbMp
MzDnhnHEktiDy3jC7VeZNwkl/vg4fa1aNxMAxgBm6yFUU4R1YlafE1hm5IzmiWzUtIA1Oz/Fl+Ju
PpeyOHWgaIYoFiuVNRZIe9g46hmNc4AlSQ4E0CqAudJiow5cUvjv9Xk416jUyG3sJsf6w19Th4tk
4Jsy2fsfPDByP9kufvh9Xj9tOoql/l2RffZn3uAd6swFtb7ORHJ/eq4Vn/ZuIw61LZy3KVrT0YHl
Ey2Xtzk2lNmyLxn4dAbvnSX+hRbVIRyqShiogVqOM9WicJxn8gn5n94P0Mtk0A93hJBQNmfdN8v0
rQAK6FFQ8ZLC4+qMWGsjFcarugs7KydA9GU++27PLO1wGlwMtVF3Eh7xn9+bpMgL3uqt2O7vcF15
62+fZZ29NEhCkxdZnftcG63S8gyUDNo65IlD4ep02ECB8MXrTlR+21K/1TRsYkWTRRcpsEpHjv6L
o7XVOG+lsOu9C6I9tyGJ/8jumL3Lsw6fGAqn7Av0gIEaEbl46gcHjqNWxhToxqGBwCB13NhbixCi
7NlegDZX8kBlQrE6ViJ0hCvDaoul+b1PuExpKPJO7FhBzFNgkSi7HTgs/+GsWTd2ZKeplkLomKMo
hSH1/FtIRdzIGylQFeXF/Wn+7/SSg5Pj6SUSdWTGebjNXVoOW/MGIyC+C29+vmagYiAPDASzxsj3
Ho3lOOAMJFQUf69XOldg5p1O6AtObv8xUpgErM1nkReb/CVzzge8BlaB+99bXD7qNOd1Wn4Zgt3C
K2cVPv8z8fXn2IjzckQqZ+me2pW17jSjYEkjgexV6c4ofdYY1vJ+DOBx9NBxp8SJ8K9qwrQtFGU8
wdAzujfMQk7Vd4i6CJ19BWK+4swKkA2CCaXeIUYN+bazSYOiEyvz13bKwcvuyzx3keDWr2aTnOU4
givtM7cZefNkSB2R+jF5qoQeyqa0UWKGzCCUxF7QKdLdI8H4XJv2LGZN2x0y8FjgWL4tAfXC7tfh
BA5SDPKkfW8AM9E0DcLuJuGrRGLwzc9HanleQ6Zpx4EhrwStj8I5DCG9r6D4vCmvN9HirufBJ5ci
RH6MrNt5iDodV9fM1EZRWNAHPw+eilcO997wrM00LucKi/pfscIWxWouLlcr1F6WqVmjTLJ/9l41
sdPWqUDl4tsAaGdOPr/sM6jP/F2+udAlbvgf3VFLCRrt2H3WIsHzjNKg1wEAnBeHPjsFgI6UcFub
DX5lBNzEJjdBYCACpAitS6RTOpw3twOTj0H5e8XYA1m0fV6BU9KkimYJpg9ObPxBXNQOVaxE/cAP
rnfL1ZvXIoHEHZosLp59QLv7jgTCBqpHRZnv8n7MOKHSUTbG7ErizgmxHJlB5MXZzxWyLc3b9bLt
9fU9MGro6BSf6CS9PH5xOvOWHSL9O9TW8MAu1SVvnzOF4/GgDQ08YDUqjEo3v49ukqoTQ3cL8aZF
ZZ3TAsmo5C9+bB06EhGtoD5w8giMp3/myGnGDywFpcPrA3lvYgDN/j/GNjS/SDmYz8k3PLXKoJ1Z
fcjoepEzCZ4+7dyzMOoHX7zhK0S5VyZs3Mnp3MnQpWs/Wza6ePgICoxHOT4rpm6gopWK1bmxBYSN
ndjBZGsH/oMgj1beWkNE23FWx4uP2O/2UaQSffIYA+m/kVTlI+GmBI6VR+tg9beoBge9mlj0IUWk
Msme6VRLQ4WpBuSGWhLwKCUp8B9talFQ8jamLA/uaVnmUh+hTPNtCNpxoIruEgmLTlP9Kpkc5QRY
NnwGAx1BxMRtKXYbzC158jdvY7fX8HCYWy95x6a4s634u/u1DnbmlqAxMCCxM5JnE14+gAR+BGcU
NblBs9jwku7Z0KijmXMpQ0bmvsdoEuUnHf1bBHR0jSQEBz080T2O6HrEipV0fua6KOBz/Ec6QNzL
CoJuI5gbVzAtHHS8xbAaU0DgWYKXTi/pzRgrfzapKvTDbZQm3tzeG0IBmWhOWZiApPQoy0VowxDx
UbbS3rdk96Mdb5yDqkp7Y1iWfJiZL+VIyS0Pbg7zckzlgXNvlX1axAribYVlhhhReea8NmWufbg7
5oR+Jp4pBR7BOCDKAvuvii2ulCYwEHoW1SKuB6mxA352Et+iS5p+fOagXwLjiYr2mwya7r6f4o8m
ViqmgZgHig5JLuvUVcZzp93rAm9OJtBYUreRd7AXCbD6Q8OyYAgsvM7pcSyl27SLgT86D+RDlgca
0F3zRW2HYperHCnLMG+FQ8SLXYZK+TwN+c8m+KCGJUMv034qJGPq2MsG6BMB0jaxLrRhGOF8hdbt
OwO/65xykwKHBerZUeJWsFyDl0Oq4isLi/lc5rAqXQDM+3+T1JJr9OlU0tWLNXjk3wq8erFCrULc
z9iSLWNzvRivvkwsfW1hn7dyPQqJgLodfnzXRuDJ20vwfwRauz66x/K2G8fFwLNzQHRf+MzuS2z6
gH94c2wLTiUyBMNnumcf+5pIks/W+N5mUB0B7AUpfo1OhOBA78ROBvv31oim/QX7zfqms0StOi7U
2fPAdGkyceLoKFAuDpr+zKapzE0xrZ+OZ0gftqATSrhOUtyJG6W8/RMhmojhwaFJefdF8R/lOffU
SKEFKKHjT6SqXc+O32pN7nTVzKmIGDQkP2hGz09dUoA4CG7wE4JuX6grxWADeXSGq1WBw/cTZbEe
jZt7nnH9s+Gkk1LQbe31ddzj3XBEnILhmZtWDcGcehT1wUIAvcboKQkZ7daWxxUsUq27GkEnVuMN
vXdFZV7/csw71HNg4tyvGHFz8lnc9UQEZbdW9AsAj4qR1Hz4ifhFcORzyT6W8rLhu3YFV5sMIx98
CPgzw6o2RsK0wIGCRJ3W7BtuGe2zp4m6CU9o2Eo/AmzbOiRQ98/3W0fh5xki/gcVTP9hx1i3IQv1
05vJhPZn2z2lsISZVWLzC4Je9CVfnmDPEYzuz7KXmIoNuXptAe2jAcHrDt9VHrOed2J+UbAIeMvz
wm5qWp7Zfeea9nnhMzwBhVp4IBSLuMSITs83MFV+AX+vrU3Dplx8/9j/cXSvUucmR/cbpN0ul79w
M9sLamPB4WtiYLipmi+7YmKZwiYfETPwJZJaO8YGo7LUteRuHvqiYOKGCUdeLCZU2gqsKlUEg6WX
vWkai8SwC3kCUj1n0+znKgJKK3JVzN3iSSbt+D/lzFQB1D2YhTzcQw1TEM9jcx3+X7XTpM9gKjv8
M26yG5SA0xW//7uESMRpr0POE/zg2hgJ/itD+HIrPGyQDDdkpecgxflP2oPEJWVKX/UXjFIdb5GT
r1lYVcu8O13Y3KrYpV1kbkbZ3gL4Q6wOKECVdXFD4erKCQs7mp7pqoBIMX2042r1902biOgvDKrW
MzSX7UPvPvGT4NT/vdLSKQAh604YmVPQjAC2bggoa4XMkmr4qqejeP5Z0FGfHvcDxTcbvcWRDQOD
9snpUVqu2sf7dGuifOuTSxTie0Ch6cPHsWfmw4ieR2DgZfll0beIdgmzJ4V9R4rTNXXCZ7wIwLiQ
L7AHgv6ZWwEYm8k7R3aYHOL/Nrd2WnpuM/HFuacTLK/cSJ4zPibIIi72Dbp6gZp5cPgPHx5DPzO3
4e4TIngLwNCW/4pRKXMzT0zMV+Fp50cPmJPF7XCmPva59JI9F9v8lOz2lu10REGrvQKOw68t3h54
Ls6BGRkYxN/dxKR3wD4RVcGk9q6K4xU2wqnNOlBXRbEWwJK+pod0gVNKFNViqGMwj4wcLDFihCUB
Csab8YnhIM1dPHeztBoSu2FiaZSjxb866s1Wyv4yD6mB5AXQigdy8rAzJao0ZN6ONC/ivZ5sRwE4
uQoJ2ShvEtRZ0BO54meU88KA5kFDt8C8y8g3KzkS+YBC1EXbRw33b77TVvDjb/u72u3rrEm9VAYB
r9kwUgHfWj/bsUzDsOQ1loDBrcEwoI9xXggqEC6iOR+/3yj6o8JFTqQiCRaik7bdAk/ilp+Bf5c6
eYSxm7fcAIB13d2fImnorjmmngRT+cOFEnpNT3VQC6TzhIqfV5NO76EizoG13qHt+3FJGpj2LXfP
4GWFvrGqQEKw81cW/CnyCt2+Gl49Scy/dfmR34TU4xXBI7vZKuUjMY8swkDTxtzAGoLYhMOMZTDa
/vv5KJjxDTZF03yuJJtP+PFL3dhD7pOSn/vKL09GPYDfVRVkQBSRbfjOE6Rzv3b2Zty41TKNGdnK
I1kmJpac175nPdq/XRvQ1zHudxn+EHXJYAhcbd4/4ldqSYf9rZajOFmmPJjuLZMyPvFWASaXQTsU
cXrx/e9QFxK1eya1uVJqMlA6+O6d4G6LgGqsUdV4640HByCs0wW3fcBsqbhISCBlwXH1dqTnNSyR
nCNPJErOFQDEDU7nHM30tlR6UeofCSavg0mXj9NmcbDah3ApHFz5rkKM0rCZsEhkwrwLcmfaPJpi
tJajNi7tcgBluY8v2q8Dxd8lJiPe3NQEShe0n21e+vb9YJjdF/xB8ZVbW3VS5/4QZy7OAyCtXT38
dUqcJgh55QnFiuc5qTKhYXfzP6/wTHCney9jTsNwTCBdlTxZB6jilRwbg4Iz/rA4AGjc3j9JuzM1
Lgu1QVAmgntNinUA4T5jup/pX3Ht8E8/4jmr11ifjvAS5TSmQb6sAcbpnXq0oN7VY2XfcTyoz0lK
xBcwBT2IQMhHbt8yrfnAxyrCaGEH7SDvF0zGupFL03ilZgjHnjy0hp7i7HqTv3+3WcjVND1kVXQZ
27dpZQ9aNi9jX/2fCnS3AzT1zxiIp8RG/RodtK4AMhVOHnDjVt00OwEcTTwQvDi+2z5LGzgSSZZH
o1NpMOhNie4OWudpLaJtoj9PnmTlDxrUXcUtlDVHqHM/k6ylfJSWDn3+xXaz+4bzw6ifvwIiY5A1
6S9kJTk6fSZJfxDHWTl7kq/TU613nqAW3RmqFXAD0+myIc4MN4V07NUgbarUf/X2vEZ1QlHMVtxn
7GFYSTolllr48oo8w1WZY/MnwuxsM4tzSbNYmxgHqbfobkVL3BMBXQIhZPVGoMnROP2MtOucTnSh
OM2ghdaGjLZgI4stJtifgtTWMNYeFrez4M1GFWVQgo2Eti8EUF0a3fwj1cZ5aB0KG4XUzIIr4DW7
B9Y9rAKy3L3wjw521hw6qpde4sZG5rbATBtiMWd+2zTE1WgEjIt7t0XTmh0wC1sWlxU6XS7LCMKA
ebrPjbgiDn8MVpUVs5nuRvphTK2f/SYJKo49Izn2hXKERQNmTPS7gqFZFWQLl1F3+SGXm/SPkLbY
Fl77no0OKnHx+WOAJuG8Xa3Ebb1W/PhmsFgLEmy+wpJsKFqjuQEje5kLju1Dg05K5uXxesnsvfhC
YsHKXNMHvjGrIHKANMBVb5UMyfULWp47/cc5CWlo0r93TtD8FwILNM286snkKvoJYTPczuQ0c+eB
x34slaTg4X8hDGvKBA/MJE+5tfjAr/yNx3EjyyeKyO42e8BOFUA6QO4LCKKUbSLvbNprqW8SscDx
0k/LzQhhVIgJDFdFZifMBJEnuJxV8jPAbhSkWzzNJMX/KIntvGyl4UqkxJ+1lc5U/bjsU57agP9s
3jVaoql3cPZ5AIdtxNeCUiKx41AGjH4RjK8OQpQ+aOxkqSDifPVdPABh6EHPYnk8cAi4AvPBi1tv
jpxROWu5q3QRFN6ZF/ujcqdmjtjEiorLIMDlymcHUIFT/YMXP0iRJkJF9SHgW+xmRtJFJb5y0tOH
c+DCgq/feCJZLplpRiIPXtrUu3etKjWunW+kVvQ2U4cqoul3EVHwUBmIW222Z4rh108SImZX/YgH
M4xWxtwP/55Z107FEp4sHVtpjh9LJSimqhEggaTkFU7XMcR9apR+F2Tzi7+4GNj5QruCmmn0AmKx
l3F5ouYhXaeV0zCRefD/aDc2F2fEgHa8H0aErr7/FGPKUOb/q48oeFAh9J8kvIU4HFIvDzjaq2wW
3NLzsUQY9GHBVHbAsdAmm8tA845tSKmZY9iTQBFO7weE39SEZftUxRZsVUlst05KI7Srx46gpkHV
sbKGcI38YeKZmAic4a+8BeXI2BBGc9QgPp1lP2ppbm92XHrxHShWddlLinlR30kDe4FKUHOtyFQI
hrRYN6wboTelvgB1Tb66aIK50Cau3bGaHstLkWKqZPhuq9neCCphSSbxRgg2rnenDW/yqqOzcWHf
BLnv4/UrGsED0Zoh2/3DRZTjeH3B2anZ1xO3RLlSSjtVcmlC+DlZsxVuN0i8KyhlYusMRN9qXPQZ
uPT1YC9ceSbkCl2918UeKhniznnUlhCLCKER5E3tiMrGgCLWEgGymMyp/BzvXLv86bXug4g5+Qqx
DpFytusbdAcosik3jJ0bruu8VO2XyqSENfp2VXIbYhEhGNUrdwOXm23ZhN7Yeno7ca2ocFsNRddH
UyhGEa6rSqea6CcohZtOFN8YQZ/+/gEuOWpOZJHZz4p+kNlf4VMJ5kqqdiGUGYS/dyBE8AMaha0U
n53YFNeFevdqLCxMS8NbQwlizw3dVEiaFNStFi/5tVypJBEyH+E3/7GZ/wfxxYEmjaIv2SHBohG9
p0ECOEXwV+mEZkGR0eBuc5PNhUD5aE54gtEi7ZtpgmgcMwYjf3RXz6TkidFNlpf4LqweFQr5Blxc
Ch/HtLTlDfjXfLMDAKAw1VaroFvyxvwnlupPAY3ADbDfOMy2UXpSCM0iDo+XmxoLCCzVK3ozi7jN
rYI+zMIRXP3ayiHJVtYyhDz6dtL9xa635RzV6YMgEAIMv9yatpcLbGvxjkixnNIE8QaE1hDa8UTc
vYiwx7HKCZ0DZ+JBA6SAhakp9dHA5dX9cMMwoCVa0T47tUF6qECl6x5EcztNUtMj1uRzDurphsju
pj3ZJwZO5FGbUcp/tjo24BCMl2Lrm7qr+n3HPWo04IahwoM1LOrHwAt+ocKyej5up6Gf7L32DltR
m3bNLPpYts3S+D1lluu9U8PGG2oXjQ183XWGAC04LZ4Y0F1GDFBLZ9j7vDqSWAp32Z41szPyQYyd
7zbNlxfyTiSrslg3YSF4ZHNZVZ8sYmzePGk1LH6W2BN/xBToDcVKxgz1yiy1qQKaUSG3rpxLW/OT
86PIgZgosIVPJyOrRnpZ7Zx0HevyjQlAS6CW8Zpe6EAPiAMZzZIALIxpYQKmffxgB6lvarQBfKyY
Q1b8xeU43Gbvv+QxuZgyAciHtfmRbFVVzS7Bnk+nUb9kFh7pmkT4C5r1QbuLnNsBpUjGGiv4tqqM
HgvO4+0oXR6IO4RVUtSZ1jxWvb9XAS+tFLHVNl6V/QHKeOxMWu3Epkr1YU5Swf45mh5g6h6Kew/W
APOykrxEwVKJwJrrEba8s5jct1yciOcTT7kGWCIL9lCLLJ5cQwzePqzhYds51oVDghj1ketOg4cC
yAuJQt/0FIoOgFp4v/cygK3bkQ5hdfCaZloHkQIn/6MBlAk7bYzROgKg7K3wmmVi/rE6NT+zeGlr
9YJsopAAjIFYs5C4pNENojmdv1RgudrrS7Jg5MABivrROzytJtsjjLeC/deO/x0Ht+puurRE/K/3
bEB63R1wCVazZDU5xW04gh6UfPoBZI+rwUN/imFYfDq/VtCe1Mo6kLcQaWhLaFGjWSJPvVjJPTTq
6CTtQWa3KjvglZLfYDstwNvLoxox5Mkwzaw8CSupvexcZZxXy+9WMVuAhiVUqdiFvO4K6gapClBH
dpXD+kzhBOvAq0Goh3mh+HfQ8c9JptU12g5fwkx48+nk5Pmm0kIwP+crSKBW8Th+vbKR/ZwVACkB
v6WH6loTsQW+kUkI4+FcycxyX+8xEUvHmYILbx0Qf9jlJfmv62L4kwo6yCqoZ4yn/Y2Ufbj6Ybz0
RdcrdXn4xEYcUcR4skca9AUS83ntjDkbslI+l6vjWifRYjNVAKupfXNPt6dzktCac1h4FfS4Pkn8
avH5BSxuQKbbeLytyZLkBSZwS/ICyqF/uN/waRCTAMZ+MEAKXBU1VGNXxLp12c/sSr/odUeclG6G
tSNIxeJthlx0w586NUz/KiNwOQ52pRdp++NUNdt6cf9+ZIYKSnHhEUbsCPG1FUT4W4b47RgSrXH+
S1jKntIYQvPjcr5o5Z51BhTkaXAKjYA35fNOrGK7kOJz/Z+VyAYOuQd/6Vo68OWG5Moh4DaOhAMg
9ZCio9GvMFpcYOZ6Fhn4DpV5W/9ne7NEYowXOwshi/g5v8O82heQK/buAjudKJY4fuD7LM7ReHWf
gdlu1eXFgxA/ThVOr7XzWDHwzTMM+jdu8c88OYvM4v0caTaZPIXEgmF/lBKqmE0L6QSpcWQD+Qlr
Ejge1fbtPrHPAepfnGgKZhE00QzIMSzv0UAY+IdLLNXdJkZWE79m2LEc1D/0wElk9OvSuP6z2ZNh
cA7vpT1CbjnWmJ2jRWOoyDu5B7FFolM+PPsWP69S+RbMd/KCg5q0W1h1tTOug0KfEOrK/DZ1Nl6i
ovfbP2GX7UUvnG26LwOvjIWnV2HRteLtqWkLOM48MFfg2tHHgRgrUj7IAZOX1G3VHYbS2zz7KWs9
9nGZmJE0KGPf3qeM4NVOYnv1BGp4pXOULbyqHmbfWKta3dlf83rPtKthXuIkiGCEZ5x9LBzvTjb8
V7e2qmH/+1I00Kp2ZLFIPcNHFRgDrqpWMWpOh48EmBDAf0jt/Dv1OI0a2ze+XnZt9Vs0VAyG5n/I
5ipWXxLCyPNjUbDcf+q0PZCVXeJmPQY5jEzQ2iutn99qGdtGdpMvV4P1pjKyywftMlr/O5HL7G/h
HsCzmhcYifZXJohPKmVr6rPsEBQDNUY634nX4/T12M/OfciGFbdlmXaJsmKfrApI8PuZ0Pxnnlw2
tVuKF41auV4iOsUT4003MeulpKb8HOliwBmkjWZAcju9ZvF4Tm57yxifYoYhGp9GXUs4iyiLJl+b
fyWfjwnlTNctNrMOAyt+ruXZ2R6JePHL21lpglMvSZ0iMh8KwYOTXJ9g6ADxTXFv6SdfXMM1wusR
YIoh2l4tMCkzoKAv+NEURpEUsKk4WgMhC2i1cH9Aolwpv9+ZiWfdJfazMZBMxTwZVb425EDT/Rs/
49gopON+ZggUYER4C7RnqVN7j4NJ8XkU7f23eLIHq4LytP3h6z+Ugx73PLOdwVMRbnAKx9j413/3
iG3Ak8YYsA591Jo/cXqXef9FA0slxvz3IxoK5JyUPUt/jR9rqsuJJsbjbtidDBqQCMgFBvglMot2
ZQItMdfMXur982GmS8WbWFhvfhYqZ9Ada5by9gFOOeG0gZ/n/XsofSohNcLLG89usgY66Z/E5b5Y
Uv8fg4ZteajJwqRCZObDu2rEOgPiokqH94dQWTGal/uO0bkd7Sgty5CGJbGpkY9ahYBHDmmVSXsJ
J2iTzgyF42U8lHRiaHVt5pw4bln3UD/jKOCzOJ7ejNSlGBdhGrbS5u2ZuRFPFjGS1aCh9zR5tcaP
3zl1OkcaXFBGHUL0m1N5bmzr9MjGT1lzUdAIec+ZNqRUyWAlOFpuFwS4zR8k8M1wi+y6BbA3zbC4
RpbVQ2PlI0NCNz1DlpW/ANeBjsppysoHPheqw49yYdmYTwdUlOABkJW0vEvYAwSheSPC8mrF2Zl0
6KgNqaEiPsYb9z/YhcSFTQbUciuUFUqByRPfxU/TQ9jGQKxycne6fG83ykfwAwgac8UlfFgB7MXL
F8eWS54Og7Hj0BlgVw4WrZydMOFO3KfFntNHaVNMHpkjgS4nfHO4PQkyBIugEoc25Yzw1P7XWQ+I
MuSe0vY18okXKmz7w/qi7R9BPH+HnzTaH97bs1bWMo99IDA+vSuvoWnrxpv4rPmAUNAHO08NXSGo
2bF/AqJ88jHKFVllXBQHGocFDrlAIjhpnzT9lf6+U2gSqF4p+nNpUcEQ8kjPfq7svZARh3BIOGtP
/sqc6ejdqdrECm9kLo4RFNbdrEyWHpPt7vIVM32ZIn3T3gZgX4wedVzr+kVdLA7uMgeZYJL93nuA
223ZFLAZCAmiUQdyOfwLkzmIvjp/1zJL8XXG9awZXZh/mkHnqkW3elckQshL252P7MFaYTH5rbw6
4WY0uNy5d9G/ijcGkTOfvSTpJ8AzrEXncrQWsMfnwUHdDGFRB+yOSanl/YmQ8QXzjnL27PIXDANt
5t1sPCpW3bZi+wEwfPgvc+J16Hu/0/shgCLXFEMWJeLG/zTcsnAwM3vwYfGuUQ6dgNmqeACpSQaw
ehqSimq64bExnt4Mv54KvYlClQSOKqLhk8RQRxxwOpYxKFYsDEElphGvXUvlZL8ugloLShcEcryz
/c8hR4ML8mGUxCxHMkH6WP8P8MVqiiB8zpwJ1f5/zoItYGNFUNPXTpFjrQDUVgmBZu1Lhq8C9gaZ
/JrCiC/NkBEQT64w+py5+rE7litoCjpLlkjAc+ad1EROY7hyUirLHXXb8hOiPPvxQvXuZi38LbSY
ktK7+1eeIyqkPCJBp+ujaJIGSICd2fnRETAzRu42H1Iey5oJ6raCsYhFICHsdOZ+y/bER2QEEImV
AG6aTicqn7ie+1kZRG1XGdy3yEfqyFmeODTnXtMwvRZCyAAAMEDfJB2ZHAgvqhAi7LK8v1bjAaHv
iYOvZeeObavSpTtYscpjT+4RUiWtKbV50mDxZH25L4DypGSSl512E+RlskjacGrFSWNriykVAsfC
T3FAcv27n1pj9WIU8nodc0t5WCrBSBBpXdhlkRVSC3tdxun9bbCAGZRczrwUz6XYBx5tTrRbMMiN
ubcwiwGH4yMa0wRFwdVi5/eBriIuUA5EeTflDM+aQk+26TILrEtsAVGJwx5BfQZjN7Cot6Vq+qbK
IkxQo0tQS5j9UWAQJ+72x/6fEWL+Tjrsu536nGFU54gznk0a8+tg7BpWBFJdHLYsLzgQUAQYmm+u
d84RC0qdcji+x8VKXNpcn3mlpWowmn4ECJHfx42c6dJ+sJlYKqNgvCUwCTBHT05Mm7bgZ/+BuvDz
BChmmi/AvLgaY+PtPI4ODOtWvFLSg523rLH4MPpMp8QxiI2+QO89r3C6Zc+1lqC5c4Lij+bwgDq4
2F6uVbinnAItJutnko+emOZT4JLoy8NQBBkhsbuoeacPgPWaRt2R8k23HDEHXWyCxO0B7QnBWXT+
+2EN4l7an9YMG6phTlKBsvMLkICnqCls6C0YjRinruPFJJ913//N3wFMCwRneiekzBDTsjDizOOu
Mr0AXSq+FMI2R7z6ElzbqTPEeomMa5toMrc+AMhmUOOrfmNxvewjA/GXn0gqetKRODlajdyyr+qo
A3Drvv9qmtFy7XpB6VonELVRoVyoQBkDLfAnDvTXbGNS0EQscZh0LMBTl71B6JdPPvBhUdmyVw/p
pwp9DUrzLIbAQi5oenTvsbEq4gMAopVIbR+7cR2c+wB73kZpMtjxhwUmOXnytlQ5WhSo5JdnM2H7
r+ug1ouxbxyTiNw6y1zyuU5ZCxs414Sh3Dyq9nnXYuBTlDsV58nsDqnF4k9pHat91DRaz/UH+ccr
MJKZKCqrovnUSw9DgVM8M3Zd6A3BzgR20JuZCo7FeexZ12y4TcUWZe0th6gtejj2I4zG8jyjy1ie
WHRA+bEcw+WjImgnPeGdgOtkDe6DI4AxypbVIFQi/R16mRvek4ffXFgnJVuDBN6HdM+k49uttOzo
SBsxaP0KaOWSdAX8qDpvN4+/tEHaZCEV5R4dgi8kFcbsCoNEvzke2Iwn7wPuc/dG4Rucyz9x4jE1
Se7ubxPsMPueCjI8kNcNxUpkJchlME2p7jbN8j6qJB15mAA3zIaFDvxCIBQf2aoonslbS31OIZJy
2az1I0qBCrknxZot5y58DkAJLd50oEuUYN9alCELQ5umlvQvunwutIpfLC6AcXUo8+UH3v7PcNin
1J4iwuQkAzC5HCjG7CYwDa0InS2NFVXixjAuhXfkPuL1E3T5Xgf33dDDo9eyTGvgf9gFZAhnWM3y
IywDBtjEbitm/0PDnMeFXnIFcyHnLFWRWYn/AYA5kAXrtIresN1EMS/Hr0H7EP921tAY94rtx3Xx
BwyT7BNa6JXcjpikRi7ET6OO7SIB+IeaL8WSAY0qy9ab16T4ADLVz3mZ91uuTdWZl9iSO7ew0ySG
sZeQIynLMeMoChYOzfgFT5MCE/3IakjI7jTDbYSAI7oVBxuQTQakH2PBl2TknQTYsBN4EohZbDCG
32gbSfP7LgPIBdTBVeM1WNU0mmQSmy01H+zKw5aEtTPOy9nGS5r9DOYMx+7QfrQeMkA9W4/CZlxz
F27gsAmE3bkgJwdlBSyNdnMcIhu4HDTIXLWt+ZJJCxm5ovEtogM/3r1vcFu4QLCHQ/6creiPEP9f
sPVARQwOZukGLi6kbQemU8g7OfQ8WbVRNkW91WuexDJSb+R/UMb+JU1qi0vEp8IVsH8KH/uVCxyM
x8AonGMxk6TctSC0xcO2GZ2+elh/ifH2sB+hFtrBcvIb7ZJZTLP9fbgYl42AEW7bc7PTes+vknE5
QPqZpP9HuWc3jbJVMRn2du9k+lDhXxyNlobsJbevT1RMpE6yXcePmDJiGi/o437rhTUrd5MPclWB
z4PPFr4ZOzZrgk7NCLXmHmFjJyJfMJTVk0T+Zx+aHePEjfTmg1hR2KWlAt0MJ7uEJiPtGtIhNkDS
4BrwG6o8xx3QS0fsdUnv84e1ZxNW9wAJqObs3wvG7OEmdFO4X3pfa3Xw8tBlI6N4mkwpsF0C8RoG
Zg6Hl6uxQWnJJJp4DpSwQEcLqPG5tRKXw+VInhKR3UE0ry5f5mW/vCD8FDXJ1WSNUlUmnd9fXbOx
C8+uz83jDowzcGJ+BICDFsDuX3ProkjkzYTfCK4rdsY/ADSVzR3LIIrTujFNTmm0ZP/HiYxvTExR
yuO0V45JGvYkZ1+OX4Ygm3MV5HLU/JVXOxOb+7KQrRjTZrWtGZxDyFFECq9cBTRZ0uGuHvvKF4LQ
t8Qw5jJX7JSWlbfozuafL0K4sSg38itlHIkpteLGQDmSKbzJ2q9B+SMmhmFtJ/+mU+IH2JCMRsp7
1yDrUqaSYi2UmbjiVLxJIatYUTpLbawHAtVrh4xKW1dTPndoyubU9Ecus16YiOyWFzQbw9cFTsI0
uWFWoWf1zhuLbK8GanCOvRp7XHk79/lXHjX2oYrcMJ5hlNh595sj2XVcqyD0b+BoCyZKu9PSF4YP
0Z8m+AR1XOuWyBipEsH7WMBPIVuJ1fPgmrQHLkBnPiHuLP/fHGPTdAPfXLenBI7auwQg28psJKxk
AjVQyqLlGzI406UP3YcVPz796za+WBPvLmB6MOfNk5eO2+SnTJVESjbVo+tHlWaEfH+OcaoE7T8c
C8YdNbU5BJEEfjgxmoaTmTzVnb2f3TPs6gIt8YWVqfYUgOCIhq/Jvs0WYFp0gwqrN9wQqvpBl47k
LkKDEwMvowHn4d/P4Z6xz35eEnQnyPv/M9Ws9QE6HB5jF+sUw36RscPChSnOQs/SVJD0yvn+LMCh
m+BnqRaBNcuK4dgHdCYIK8KTuRV6GBDT6Y236y09useSCVBXTvXHAvLLgaRV16XmIOdg/EeXmwXz
hZmJA0awk23PUfNRTBxurhyUh0tg9y+IByyiOm21jp3Ipg7PZ36osryJrt43iJsr5o6XGnJu47DV
elh3mRf23wQWA+1LmGC6jdkMSWOYeD3LCOhyb7tf/pM6BdctqkwCCRDnUx8MGKS9vHVyBJEilcjY
JZs4pOunEtvHkMWBK/eooEYgtD/I/Mk6lm3OFe+uFncKFp/nrO6ww3QPpnasA9p1L7uI275SAKaC
QsbvMH3g88etYWi9YjPNOz7+2+31HSDU1h9x43OfJNr/jFKp4hmnstPxfDrFgspD923DIQcI4gG4
7KvplfkAnNLK1N6u6929yunixUvdQs5aiMLVeNn7zMhy340cV8OkV50kHRQzA134La76VDOB//AC
Vvm3rj44y7rdTHTn5WbeaV1YyIfz/sj3Pxwgm9kOFnJYptNrCiCWppmE267/6cWdlT6aG9i6eAFS
Us7/JdzsDYqS8wG0IU5mp+FzMbwuhJqKING7pce8kA4EZjcbs0eZW9kBRm3vYLwMSITZ3/E51OeV
vC2go5Rs5pnMPg9C5nNSQch9YvYehOuCP0CRjXhFo8FOaWEdB8Z9HiwR4zzfGrU62xT7m44NKObm
q0bOk8A5qaL6iJ0ObGwqng8WVJShlBNW3whef/w3cD902vLDxzxW9BQnOK1xIyJjwCNGGoEgmE2/
g1UW/Izh4YbwNp67kveqEGsZyB6C4T1RewH/G5fzxbELmEbT754mN6xwuPBfTRT4YvYdi8E8y5D1
LNDqzK7hiS2/thPp5kaHHfXzvoxmBXQCnTQea9IbweoEsvjISRI/C9JFsLUjdzpON3ezt9jlwSV6
juR7hHKd3ol8d+VudZJeFTxkPAAX06gQfo29yWSptSfSXH1m3W5wlunHeYsO505ro9lHrDFEao4o
Nnokme0TbjbQGiOJqMkrO4+E5hnOcvA+3wKVeEniPazYyOt9fM4tPrkt0P5gXh7hjR8MJnCmpp/d
p5JsfFViVZcfE/Fa9o391H41eL9XEZ49qwbUBPSlmSIAYVJM3UCenzs8tSRE1myg7VSGZdmbpBbS
N8oN/rwdVWEcQV6tW8H3S/QFjagisZSVkL8a5zhCHCM+1k/MnmJarYQxa7YkJDpMPcyEIIYyK7yX
+yPcvEuWgyr5W4q6NE+si8vB2QzkKwfRwSg0Xiyia+XYopakZrMWAKTlhpepeXx5QsrueUTA76fe
2k7cyjtLZDhCv9yC/1UlIXVsBIgeG0oa1LofLtYZHSLU48nrNzaM4PSo84hzpPs+o92PDP+EwZrU
qCakKtoEvZJc+xJFIkSBW/LGMjsgjwM/sy4lYjxy7b3oBjONSkQTKV5Vhv59qRMA01OAn3bL3YEX
sLLnhhpbUOohVs78rs8ygIUIFVl1/yFBSEIMI6/Ka+Q63ErIynW/lL/+qyYsyb36IS6gt2qKNa+N
KKx3TUNAsWNMELEPytxtV4U7cFSe45m86Zev3DK1q6trStTce5h4E0zvtD9D46GP9Bk50oPYKBZj
yYJqktFLDHg/B4jak6wdGW/i8gnGICSxeQQi1yzq8V3eJoxP+qbJDfZmeuNjpH9RN6VVgV08f4c0
pYbh4py2TwkqvlJTOfCRABib/NVe0h0rRsbtLx7tZCE5ymjdDDrUwtRgGbS0UMDE/l1WR0STbE1+
xyZdopXRIfMW0YDtYdTqRb/0Irt/h5FehztVWceyrrqxEv3gQZc9eeWZwOyKcw+xYdbtRV2hhDvJ
hVAqsTOMSKnCVkwy0ahLexjpa/XBfxYiOEWOs3Iwbw2pQGwhn2B5oYPOCjvKbaAPVeV+CHT0+amv
BJlojdL6kC7Ql9iJ/Vc7qgVsKJoh2HlxjMOGwNqRZ/p8Ta+jBBCMmi+z2Ethuv/QKLibsCbJIlrb
QjKRYSh3MS3EFABc65yRqErbwSM4TclvZcbEuQF1hNJbfYkoMzAT4i3ZjNXzsUupwObEKgUPAv2H
DndiDxSutOGfeQe/FEGh7vR2mnlym/9OxytapqSPa7f5fLvuRDBLInldaKP8PYsOWt8n0XH/CA1h
opB3ee/hURZNm7Fy9DUsPWIXhRdPqYCsP2Cpzw/ZglEguiZH8FPZTDw7zb8tgPd/iVWlAkJulsnb
Un1RdypYldu+afTUsnfAg9Ld0ZijdmGIMvw9yVLLeybZConP9FK9TuMN33w9x3Zm3Hr9Ahv4NOTI
E+zoo3hkSFV0Oz0dvdUilcWnkppYQhFJxqrS8uMLiZcFdSZy0k2vNQ1lu9NguHytNlJJkPgR7A4o
uEofOYcnWbU/RhoZ1ldB7LjSeb9CdhQ+jjS3pEWhWm+10f2W3trYyKn3SlzLa2wnyMAdJtPLTCoV
OXu/9yqukcgWE5F7NJo6Te/AWJI7y7cAsVOBAfgjeDpY9a+q+40mJ0gfJEezj7vS2GzTVuXd+bTU
LOxmFDRiG29ylt+9sTlwTMfFdWAz5hskcy7puKPfFffzNqCxpkZ8P8v94eFKRrZS1qwuIS+WM1di
9RWXkjlBDtCIoNf0R8sl21tIbw8uxOBjd6Wdp+G+vIw/PmLTYZRdOlyIkTy2CR5ZvSrS1qR5eMiZ
DgAKZqGEc2hoQbggOX2qHDmFpRaQhaouFcWGxCBorHY5OO/0VhNaJxrvXk/XYr1dck0bsPv1pE/m
QupZEq0kbO5zh2qoY39NNJ+CpkFddDJy9+BF9ZKfYqj6yanclluvrReJvlfXEetAaq/EZx0udMB8
OrowjLWgqK7XKiPFvYmXtts5djI4Dq+Ed/DDb5FFzs0SWL5qdht4U5LNCL4YOQYWAl0WTYE/YgLH
HrvuB9mOJ2Gjy2EB9A1guahd3rvzf9Cd1EocVVw+GjJbDIO9TdmbvTA/A6zIXZS1s+9suto5bWeq
AeEBPFfUInYjqkxVLe3u9l/Odoe8lS+PR9eb46sOs+9mGfPtrMHp2+RLLHM8EDtkDxXUwg0v8I/4
kUOs5y4dUC0we7Qqmm2auNuVyAbChlo6zrHJfpoGNSL/Oze7M/5S9tPfvcM1gNim2tRcksy+sDnm
1/kQ7lzkki5lWIsRK7A9cZwGyHC5phVHT1iug+f5/2L/weAEoXA6MWmdvhR0kXc6NnCJYObtnHqk
YI2/oe+WnRrEzNZTM4Gc8jXMo0/M6GEy9UYKsxZuQao5KtKwWUJGyJ+DYBwbAhkR3893kWS8XieB
i7Vxpj5LU8TfMtJmkCFdODuqAWPQOuPJCYYBYjkbA9nL9bDNoNKczYFg8v4ZkpHXyp7Jj4USRY/1
rsVGDuT+nM7MhVsXTuGdjvdFzro4kw/qaKkjTiwJshAtxrJSbMBfT6UJ6O5eutwOuCEctkmcjlJs
/btK4ulDgCBj1vKA2pI8qtXlIn2rVYmoWFbY+FqUAOZV7oqD50OrDZpTqETpcnyzbz0WT2yEVX1r
8KQPVuVbL+CRADjbMsRKj3XylPotFs+o0j6kecZcx+uH8eAwxZzZP23XozxQEfV4RDlQObZJGJwV
pAfW9lyrdK00NMU6smvmnZ5hANwR3Cy648DCJkDXl7+Z7EUCf/yCg/mzb4yRDGwcCjloBIG47Wdr
qqMlDoWikzl/5bDd8z0bNdpC2QZLtQRiDMJwmEJq/cZVTCZsrI15uygZL83jBKeJwAN+J1GXbUEx
vEtR+7ZFKSRXTKGYAqdvFV8eVLgFd+bwGtEyhpx6mPsIYdGIe/CTvVxDHom9cFKcCHS+f/nFuPIN
pSMEjBB3h1VKfMH+GAXy1gXZcwyhAqDFfdYqDkFAYF3a7q1VbsIARZWU3+zJyvMQkEZmkXxLIqFh
1A7efhTzkcuFZGSQqHgccEbIF+Y4h0jN5iIKErrRt/njAFoR0Dwxj+RO/Bvk93rLZEhWY6daTmX5
wnb63OtsPtKSemGtd6jA9E43biwkZi/vzEY83HwNdUCVj9j9r2dfWIgFtLp/hPp01Yb6v9R+xV65
2LF3gtLsEnBnaR/UbjxidWAggGITM9N2bVeVb925ttYmjf+a+95+B87HP2AyrhZniWn9m6q/hm7z
gIBz/JnAM/Palslw6elWbSJzVSX7ThIuCPggtHvdRmdkfl71qJ+BLRb7NhgcPNR2RAxRs3yVVjGO
PzgDShEbOSNim7zRR4IgE51BQ2WepzYZu1mHkCjxbBESCkxlG4yvjjocxYfECMpwggzLnUsUslKs
3JhXBqJg1hcbYEjM9wkoJi8wPRWh3Q3Ft52BAkAsyaTHBZQzkbaXkTQGXsB6AfBYN6/dwCz6n6Gc
DBAh0OlrCfTZuJMNmpS04NrpGDG5Ti94RHT0P1kbOl8sOD2E3MFlByIt77vGL4H5XZbWvg79Rvp8
ME4TP5mwz4GrU7S5O5R1aT27S14pH44DmK2G6ODv/x7BShA2undwDm6J6XPW0NMc0dE+EQqM1rQ/
FJivM/5nKMfgW7n9HYRxCdBroHXvc4p4rITcfMZHSRb2owJeq3D7SDilT3kP5xe69E0t3OWXrbBC
jrBFF2ItJUepyiCMe8kG3PtO5c79VMA0ZXAJKaqr454rC/pfRUshZPJUHsTArxsJZ639TYbGhRnp
jD4UCidT2wyxcZiDNdc3BEu6m1BgzciGlpdc/IfSUfB7MjkWRv6WL4uAkXMXijnZ4I7rhacmUhIR
itN++w2ZeS05lE6kwH+1uon5IKXg642SrCMIwunMYBMkocG//vcw+lYBA19kyitVdax4bBTRtMpY
wjggbg+VsyJuUL4wDwDY6EV4grMzYNvBztEHHv8JaEcHbQYOha47kXI+RSoPt7EsZS4NSMfrjm3x
01UZKM+JTnHgd1svgLll7oEHEBfmMOvIp3xDDMChlyLulXnhVDPjwWriLngDHADzU+mOCPu6G/eq
D5YhGCWCkBe/KR9vGAK4y4qiUubnP4p2Pp7R0kMIr3cr+aikLdOK6WoFtCexrnGBPaI8yJQQfZYi
5LCsu+fhxJEunV1qTZ33GVZFOj1Wgs4T9/m13PXXbgmlAZlw5Jw6K3DlnPNRcNgqI4avAdvHrJYw
7GEis0Z3AhTxwsD6Zj8APpGtpsCB64PxKbvsXZmjdBlOSVnrw/BSISja28HngMcYEvTIE8490udf
M2XRmKsZ+H85SCiYw91KcQ7ukA54MB2Vz9FYB1hLlyARSw7XrEMYG4tgR2tKu4SkDnBXM+pHROzr
B4P7PeMMjlnn7OTUgt9zZLq85w8WtVuwTRvoEsb9G79KH9X9xzCv3v8QhZT5cH/yq/eTJx0Se3wK
PKnsd/ZNLYJhFNhD9/9TnYJ6H1kprtFINIhyrRKwYehvHbO1HA8INRbahwEmAY/fDcJ4mm2fXrap
PEwnpmZBdhyFp5/WXbyfFyudmIROqGp5syPmYUnwyaUwMYyhNdFrrDCvkE7uskr798HUw4MDJNnM
+DCPJVA94pL2RrdD4NwInfh8xqDhT+9rToWQq+ayN2ix+Qf8SRaQbSHAIvnYFswmmswgsJwVw38I
D14yJWNhe/im0GOpI8Yu9GcLgw2FeVMi6kY0BH/zq37Xbvq1S38hxJtTQ3agijNM0zkjcRTHWjyQ
GJ6NYm8VozXvvfplcwBxSVH7VOb3Hu2Mn3QFbdujx4GFSYOOaRfmTB+7ugFBHxPWxQOe4mL04HCC
4bGhAsboFub2LZK8dCz+XZyjPI4gLdpz2E3OR79JkilMYImR1WGJHTlBLGag0jUAvrC8cQnRjk4s
gpZtKlWY+UaSMTSeeokSkINQe2sy1+/wjMMTSORhgIRdd4vUQoV0T0+/Xs9ZsMXOzzGkbtRazJ24
XLlmOEpCgdrpwLK+gs4z1jprZ9tWicMOw0tisEKiyhgPaonN02Q8v6eLZ89E2PpupIIwbmH4CavW
O+uXgU25HlQFvgH86oAuA7BwjBYLDoP0Sqev10KUcZzdcbe2TIaPc+EvN9pvDz48RAQ4qzrmklFx
5wiFglaxC0TjZ1d2sMRYbfEC+EZ8pVHwlJYjjXTcNBZEjIEXahxzDC0N7O7vogatN9xWoZXq8AkI
Y1W4pph94LiATc4w3mLYG7CBBA3ik8DUuXJyIMBja4qvhX62hzfqZH36be9YGV8Kcl2BSNIv2e1V
sxZI4qVRjMjDFTxNig8WOUTsOgSde7qRa8Zka9L+2P8iMc1UcYMThytwMWzGTTkrirUsTd0+4h7b
Z1wefmmMI9dHf2H7TYPuGQHo+p17vRAkISknSg2miNEKFVBC4s+UQ6OkcEA2MChyhGae78CWGsp7
OgjqVLu70tLHoN5NIaBHbVpySNM8fTi18I+zgoDGeIPSOlJQtUFns7ga2n+hy1+feR7iRl3WCGS/
kbgTzUZy9oL++mAK9T8b5cm5HoAeOAh8mwXCK3f3cZ56TPPufEu/LGr6CjDGvc+UX+xbaoZOoDMv
5U/FYR8K1mGqpOD25x1BH323DtDlbrJHd/psIeSW+yxPg/VCcXHn4SMZk8v+7xDfGmqn9yKGtc56
40+e3DhxyHJ4KhBmYLrUccfoaI2V6vpORMYp46GucES8RELGTNFr9e91cjCSgL4znBMUJcd8W6fY
i31JRB+f14meRWb3HDrN/qX/FiBqaBBiEvaqR/r+gsK18cFRkJ1N32oLlZoCrJGDWJct7bygSTvc
JUhoemigiqTUe9RODnDXoZQwySi8TmaQ+l467S0HbvUH7+pQbZe7xmZafDsuD008BSCtTugAxDOk
eb4+f0LIvNesd2eOweZv+vbvPrCNUrsCL0uZtRBj59VhL6xmCm8vW7reXJuLxp2++xuaYFCrzcRO
w4M7vZ+xl8lgom+LziLEe8uB+4f2nskcs+VQKriPn7u30b6dZAXdyLblBd15y7FbIAykGuqOWkkL
cfBz1jxPmfegOIh0Y0HlN7jEJpwW0h3Q1lX8VmD1pr59y84hSuKQXh5yrVdpmTR/c9phRWgd0KZW
uBLiV5l09+AR4TelusgOZfp5ZrRkdGXgbfjDRFOhtNDsH6w/7fTqFFlvl9O8iSJOIHmrdHpzGSuM
wovWcZ+jlzUlrSO4LfwHWR2m9PeeOcesXP52XPgFOrvceNl5hxhxYt0o/zSLLmYot8wwWCcJyjuh
vojRF+YcQLxBBr34ouyHsYJEB3aKwZtAu87qntGD0fSxTuNkCAMja7ZdGB3ySFBGyGnktiMfZwEy
c8fFRZeFY3DYTUk4g8aV0LAEsS5Hd08rrF6v1A63/UEqbWrux7baBKWiuFygWs6zzPWiWyuoukcx
5g1UK1PdPEvOx3bFmduFyu1obNs2js1lFlEIIxWVoUIa2c39NkGPOGw+rXlLTe8snMAo8HpdemMq
osw4G1KZEjvcZ9tBTFgmeDkekyK1xaK+9ZhHko9fu7e4GzrtDL+rpb0w7wYn573I0cELlgan2fr/
0WrPY2OlvNaHL6xkQ9HSL9sJYpbJ4I30iw6wD7ahcYXG/zrak6Ju/MqDzIZs3QcLdCN5GJoGVVVA
j35VNFca3JcxEi6WMmJY5If4kgHV8LBiXD/m3nrIG2at01MXqc1QSFvUNSm6NHyvNKO9FXzJjXVJ
5bA6SpS48bC5LG5kYpJTWLU55hT+qNr4Ad6/fKwVrmJl5bvDhdKYrVemYxj2nSFbUGW7oraIuLWf
MIw8WM/16WGLhHxzGMDLIzxAbYgO5sl00/yXSuBdQb8XokDXzqnmtESd47sw40DhyWLAMNSUD9w+
460nY6OayMgd2wXOA7xLOOdG1Qjf5Dw1iE94z+X1zxJK5cUft9pFALbsm3doozEkq9edko8Z3P6f
WirxjxBJKTx/pWCigpmM9ad+G9XtqVk+6UlrEDBEIEmxRKXgRWKVBU4rGVF2MEVUtR9aBTG4KLj+
4kv1VpttQVUxK5wIYTjtiI9x/a+72G48wyX7U1wuOPrdX5xrtVpTrNVvQRxsQ1V9XZxb/xPiq9nS
1GgVU4KeAxHPinuUcuF7VsLes2nYFj+T+5rpt5jVDpwAmX/ImcwRid1CCVZK+NZGMfx4eAnZpbub
MIdVqP7YHPgSyBI1Kb+1Fxv35oZfdUhM00Xwd+xKxCwUcnt9K771y87JfBqJsw/NDaGmvc/K5dfX
1DkY7l4VCpe5rrwitEz82RyL2dhbAyTFcPkcwhlJtZ4vE6L4N4g5XsP0PrgZAXjhV0vndpXgLbsJ
gqs/nA8RSZQKuPxtBeSFXt90w6nlcWYU0Q+EZyIlDLl1ZWkGSe72i+8QZsqtQrq0KG4XdWJLUQut
pfwUMAGLkZeriKftXS34uHJ2ioKtTZZLJy+wMAf82GYkoCw/P6d42F0zdsUyFq6X/GHqp95WuGw/
6IpjowuS3RR0OdLER2ZNKWVYJEHSFPG4GM+1qzfomjZDoSBdYtjpFb4vYZcxdpTBgtF9olfrGW0k
AhFZGRczCuR1tIWkOrH8y2ShYCp7VkA3nj5YfjcIEq2DPREP5ArOChCXjIc2ux4ARotxwzUBecol
ubuBC8DX7THv9dAA7Dhu5tmw/UrI24P1DvXOP00DYXlUjglWVUHiTYWv057uI3GZ7OlWdT3Usitg
zqYBNmywgsyoDJC0qBtkf3Mw8bTJlxADb9tsRAvZuXCVabxG7xW933EKQ+pn6EsHHAyc+cthJWst
0xIYDXcf36IUZ10kN+Oo4kII0KvgUDhmKMM0jYkFXzg47Y38WR6dnhGTSLmq/ClXoTXyI38WIgwc
j7nsApDOPaYVozFmc093va+ZV0EXopPsjS5VH1zHLsObQHh1cu5kcrv9LPn0oKBU3M6XHyWRUyny
mLSJSmhdQUCD+9FWLbJuuNdzu5Frsld4hrp3tfvmyuA4B8KK9wTQeAwoB7rkzbcWmCR1KwNI1V8P
0WF1bGC6jCxsv4pujmyTtokYa1eFtLtOuaUB8BoVVycQmUr5V5tWP8ho6Y3mHdTra3XHb+dvOOW7
b0MA0w3W0vv4vSiZTV48JD/Gup4zft7rkmS4pgHdnvoaEFu5jkfpCaG+fa1IuUIZFNr4dNUtohrA
3KeD8pi23g54635PG+1S7lOhbw4j5gbPzEuMfOJ/pcMN3W+izIyquqmQYoJqGUxIr8pLNorEPJAG
b6JY+vzZWDE0HNp0pxZSIXUyjSTL8nHfgUQISVWNqlAxXPtUlSjrEeGT/nk3AOG2ke/QoiI17hwK
zz1/NCvacnUf8cqQwmeLow5HsCbwcoOkUy1wJCx6KyjZZGCZb/ggNaFoGaAQmYf836zfef+0MiGi
4WNzTuGUnJ8gn0EDnhrO6pG/0VbNcpLXZR1ERDQLTIZyOk+zy+/MuQp6ov1A6Wm7PEyvOb9jv9tp
POzm5g/CbRrPWtV7VymUJ1rQZHlyPLuEfspcoWCwLhwzNoBMxlUjctbTkdFzr/lOV9ftSpvSyTi3
Qoyz9VpL+l0dJjbvSSzBEwbpWxjnFU021e9Qe/hrwTF7khsz5s+WEZmrfyUajpp8LJ3l4Y3J/KMW
4CWMzySMcgAp2/avtEVfudj5NWJVVRjtUUVXin2r3smrSMxhThI+0fYM7MxA2Tj44BWYumMIsmjp
W40nFzSUaf8appXkAQtUeJybJlFFXVXHlB9fsAgg/HuOY5NPMGE4V5VjsWMbpVpQpXnlIJ9N+E6u
/iISRIpB8eUdQc4/A8uKPmCl58UbqdmHXw7Rl5farxX/am/2Gmi3dmkwUVMSICqGkt1Hmc3Xeqk/
3lhjLP9e72/H+VCIiL70im+dGpzr2btw8CQ2o4sEmzR0Vf7ggmSdChSTaQuJ06DEnPOylDO6Odae
USGWeKuxNp8pYUbH8YyWZfgQ8KaKG4tkzAkzWbyJb9O9Bhs2iMmbfCnhXWJICKvqvf+5BAKDn3Q5
vy5NDHDgRJZwMoTlKIYhjCAIK3Cf7RzslICUjbXECa7rqPDYTFKvsxarvBRIw3S8iWxpdumsdH9/
KoJagbHUWHtes/5WmpOlqM8yjWVXpsEM8641SE5CgpvysLWjug0Au2sbITbrJmEOHcOCjftMi+8+
smAREofOFBbe3UM1bKqa9O292ZKyl1reYgJZQ4w5MCkuisUJDay1GgUMacCieVqN9MXJ6VgJQ++l
JkcQJdvihex7v40QL/7SUqloOgv2dAgJ1jvTAdhuA0nODGURAOzZKtoy2ldy0KUO6r3pO1rwngze
R2ubQk0fTCqNHfqgmjABKrD4yOIuc6gFcBrBSH78prfAOe/21CueXpgj1tuKyzEn4WZNkMnU8SHe
7dAAPQzP7z199MWNnLfzoWqXIMQJIML8qRFDZbFMcCpMTkkTF7/byvoJbYyDDfr/TX+6tFFP90Sz
1GX1fWE1YKjkyoUVRi3kVgmyh+Q+FN6jWgtz+QNjj9UBa1hOqTFGMkU8OSIbnKno7SShBW8iTMFh
9fzrxjqkuuy4iw3R/GOjRoOicKVQ7D6PODcyrrRJs9bSlIonHMwDo62GlP9dSn40eYy6zUJCY5F+
JROVAORWjk9vbq6cNGvlzVi5ZTd38gZfWxpI/ibTnEERZaebvMPmudyasliYc8AqG7njZtYw1dWQ
YEFDVgEUwkRdBWHVDUlQ/xEa/BIKiaVFDd+P55gkEhsgypE8A8HL8pmd0V3/24PFNkOOESgIxnn9
RvxfMMnFUjbeI5D1OJjqiz0BvIANNyWE/P0joU5veiYZExyLVqGiNPnke1aCSbFocYhWW29xAJq9
7/cxtglcfOjP/naL4SuuUP9eVUlHZneu15s87vsVE+5Seh6D+kR7uNw/2Hi6Y0wvxHMXCh3KY/J9
BAdoY0vEEn1I7Pr5YetAycmmpxvyRnt5EMAIHefMjhVAfBxmAz+Du5zDCeY5L7XDyE3Swq7plY26
keshs4EmDjBgi/2HcVLkh1dyYfAYCHbZ7QZ05GZQLl4m1loFEuns8rDs/DoTxXHGq1dcuQ6XbHA+
ok3E2TlI68bhrGaDLWKaRyK/+6rhIu7FIXwJzV8lOw7UAV/lhgYW+4QXCxA92MKUPs/WDK3iQEZT
Gc1S/V4C0E52wFR+u0Qea3S0DBoageJI18XxF6i0G0qkaVtzxHwuU+DB17EyBcvF2Lcb2tnIcDE4
TpgVMFGKE7F+eK6t9T/hsUS5ZyvZsRWoB1R0SLjMTuCKNiNKZWNFI/uy5TncwO76UTcpNethM5ZG
916+XrL7TosAPGttfSKRIQUgvsp/ztzKColoKC/1Z9FcfNgMjvlcnW0N4QKGBBtI8R1aDUTUyrrI
qU5m7HljGlBbP+iFM3upihga9X1lxtKvkLKm/1LObEu8RKnWmx6d1qH4q+cPPcbX1oG+cHn0OPbC
xtkK3gkgVkxBi7SKT4eky3pvUxAp8NtKGmF8WzhDWEh1zu5SJrVXCcEYDtgdgkYdGOQAORdKTyqk
plEqb1Pdb/NolegRaiAMz2ndht8ONx+y/zhrDShxl4krUqQlHHoASJOqLwAa5ZSrbh8zqXUtd3wl
haQmse8BKuhbes7YASSwwi9vRx7kuQCaMGiw+DHSEx4s7tMtlADxRfSwk/r4Boe5odDORPlJG4Lq
O8k1rqxcwZI3kJyEyIzZDRIg5oZiEkiiYOzPmE7SoxlXrQr4WtwPbJvjKErBTsTZlfIyG3ZFk7PR
M63L6CjAhYbXgT+lHT/8AQqMHY5yk5yZe+4p/O7xik0LfS62OIoDCGpDXwLsdyAhlcpGM7iUGkFA
I16C9qtILBgvPEjDniBxAatxYwOs0uR2OrhQ5VpZA0Zf/2K4WbTJrOzSjgafu/U2R7TiXxgrvZJw
+tvQaTLnWPj5qZYEuKD9kPS5eApdyLCqiowzWqqsWu+CGzbEiyeW1QNPcmpbT/PPTaGUd8OLoIs9
n+/eLIKOFZd3Mv0BwlDe1HLpgEpWT1WfXhqYQVx7YdcvuAU2WhclW/p2Mfq5tJapTIIG1Q6TFOHB
AYZ1yeAzV94c6RwEGiLuZGV5WvBfCzia/bjsXQ5UQ8epavkU2LNMv1KWonDQChEonfiOm39iXzwy
l2rIy1QoEtG4pCodHHyxI4OFyYsvbra3/FeljllxcQqV6ppkepiToLEcbppCFXxGZOEoMce/Z7bd
kXwo5ONJun0LFm1UdNm6wQXn/dvsAt+uQUaXYnH64kjkgocMweaXO7g2srSWmDxT0P4GL4ZwCjWS
BbSh9gnfCFEioCAGXmwZzmi17JgTYlJITg/U93N57XDs+ZGul8wqKwEjHSlbZ6Q0jwPGey/DKVWw
Vt2l651izpsP/sQIIO2JGQmbNPH3c4FLYj6hgBE/7LeVndHjQXTcHut64oIsCYwaiG9omEL0UWuV
38HhebFN/66yFqUjWdbYRICKXkUclbar6flnlsWt5MTbCx6iDY4kI7p13PA/i3fOMbP8Ws1+RyOV
3s09RnWGGLbWiDC+hfwIrIxtGAWvkKR+8i/V2h+JDp5uoxzkVjio5MSXXb380HCIea6nkRgrJZqO
V8HmNqwEujgHhqVjiqx2nitq8WWehsxNJw7hPkxF9uvSZ2Vnccf4aTiTqWPY2BaF60NuYpbgOunp
62ecyhNibzbilz3/g28IEHFRdQGvGrgAqNUzMdiSYZB2yCmBdyC76uQ0dL1qMKWYjOyt5lBlkva1
c7u4D7/ipdVc6I4o5qccL0AD+LWQQ7Fi7868/aCFMWMWbirnIXnqv5lmRkrr81D2Zw7zgiHcPNXN
gQSV2Y2mOfCpO2us4Va7uUQSD0ogBYWL9Pnh+mmO+tiVDeO1q0nG4Zx+jo4Z5TLpvR+WvNODbTEe
PslxCjh+QoQszWyjJxrxXfjR4Wrc1Lfi6/wuxbgyPmDB+Spt5GXnIZR82f6m0GYwBtGWrcZqMBE2
CGAKdyF6nG+cIDlop1EUbqojgbn6ZuKCWxy9ljKUWcKPCOzeOpszqSyLEoDCROmbLmMx4FOmmoq+
JOgcur1yiKpnTsY9FlpoIE0txnO0OfSaYh6BA7zDZ4fetJYm5WzhiQM3/0opN1sN3S4NezgLtOml
ZOu50fhcfEEw1CFLhU1AZPnfaIk+nmjTseo/t+9tL1SuGj/cxNdJP40atd5RdruePj+Rq6wztGuj
OMbdYKPzsZGKb3KE2sv6qmosX4bF/qHIzNtbDY23DhBVrNjC3/wqLpUTKTkBjNiCNawG9II321wY
v5S7/tMGSF42fFbEQmzdt2CXmAmXZdeYDW0J7yZTJtTqiS/LXgy+6gtSzxzx6AxbigpF2jXR8J++
TpgxQ0eAegm2zEwAEmE6SaltfBzMxib0FeBDEA5Fz7rb58n/bsoAkoKMtYa75QmRAnQa9f5A9CWm
PRmHYgnjG7OV4eFpmaWWWhmKR4lVFWPmooGbpCHDumaw9GZtkky7/+YiS3bbv3aqG7EhwvZS7Q2s
ZAwBSj8h5a/p+nTe4NBuT4zLOjuq5zGeqj0t14d5WNe2ji+IBoPfdulSkfOcabB4jNrj3/XRR/56
cohfxZgzFZd6zczfzrQotE0Tf+71jalA5RwXvGjxcmS+J1Cv+8N5rxZ640Y5Nx2PtDTZC/0+Elwl
l/vcrAAxhFx9hqDRJJWy2FuAa+iJ9NXnthz5jCmpD4h8ZULig6fkX3597UlxKPKnW3CvLViwVnY2
kssSNlp1CQJcspem/3ogbjad9nhgIjztHmN4OxvSghpjQ7eSucH2ConWx0GCsbQ/aSVJKFZ/vypC
4vZbIIHRs7wkKjC3ASNjZzOky1HrEMspQgmJ3yYa6sMCyoTHRLAdMT28wNjGs3UYPN5cNs6+bsZd
3Q2nsqVZMwAhrirKiMOot0E1XLxFc+Mzh9qOQzrz40LTgdab4GNa9ievPjM+Pb6mRHJSkbNdkZfj
ZWdGsV2G0eC2uoO/yzZDOAXgfw10CLknLMOAEOD0BjEYdSFNomyXG9mwTLzs//oxs6KiE0TPP26o
JDwqvz1KqKg+FhlLU+JiqgN+uvzfu2XDp1cZOgS0S+9kaCXODT6TDKpqFwFvi1Ct0mMdeE8d3JOm
rr+TSMx/6pzB8bQL2DdY4Hy7sa/RnswDlwRDjkro+wk7orpdWtJu5PedlhonBnNA5Zbhp153AK/b
LBrYJibPEfnlJtCQw16Or0vOEe0eBYw52y+fywlN/cYk8QBGBQahOqM3jmbv4QRN1d6BYImjEmv9
K+z+Pr47WcJzpvrZnPzt52AUBhyBca31c4GyDOb/6PsjYxWs/LXBkeXee/rz/lyQFK87J1eRcc95
hzoehc6rTy2vuuDyto9cN/0sF823ssmo0K4PtUjLAGExf/7I8Hza008CjYzgJHeyVhuyFLJKZ3El
1dYwO6KoU7tMkcz9AMJ/0rx81WY8M6mgNbHZRwSjBsewHnX9zM4oGiFXqeKyI3icjH/5uSP7uvB5
+5KT0cK2vIVa4hT80w+UKTXB3zOeXfwNsOzAwS69NEAh5g/z72Y8srj2s736qMpWYEcoMJOgy7Fm
TZ9fh8MYgmrcthFLWOJWYH+Z1tfrfjDyMsBOUD1MOrfCBaBK6i3bGaFUEn0wwlzckjtt65NIORF5
QQN1Q/w+Zf6q7PFoVwnAabc3MUheIVHuFfcv9wA7sFMQe615UevkSS9B93SnlrvNDYZDM5w+ie25
xGLPSjDu9z3RfTl+/evjnlRB8QkCZpfIgBuZbARtnSijYneS2/XlPuFZ13upBAlAHsLAyAsGE52C
/T9IxYgrS30tdyxRRvRtEuHpK2jHr6Kllso7bQBylSlGnd0mzz6/D+slPjo/CQgciqEz2QeClUdQ
GHTpTlHW/ez9NMWNHlhPss97aSMfTA/wVLyGljg181m7fvTBgICk/XwtOfAxdkEL201lh0ZxRLB8
6ElIjKHdEyROKKRgZAyaNlsgN5QujD5hRZhf9b2Raq8/BzyERmmufwKuttjMgaSb6fdUJ9Qr3dhO
st7z78UI1VLONIJDzLpvrSyP/9VYfKRXIcydi4ZRpx5FL4a73nqsqIiXdVD0lJFSvVSIvJiXAnAk
2WgQy8TyT5MP6lvbN+iXFjGhG7irOBPKj1+b1bBxNA3Uk3f1SqIx4LFH/o8hNnNWxZrIeiWWTuRK
nB7nunDSB5bQxyukLiCOn6CnRp/1TRYCR8hkGqdBWSV+b0NHmVncHJgUoippy+4JcR2cxy9rzxxA
OWc8hJb+hV22edLvW6DaovL4FZz0/P52oJtwWmBf/5xUwUKf6ghz0a6o5BbJQt+Cmb9947lJClMA
KjOBNzL0BqFeizdhQElt2qUA3R/bKYxFrzclSMvLaZh5qWl/W0Uon0cZkgZZ3hmVC7dLoEf0SC3f
+aEA/fPGXZzxsQK2bioMuPjiJ2ewcWD0Oev8RxCIr6FdQYpg1Ai4gZysy1USnlPCAxS+WhmC9GWF
kPvRuT/XmsjjmVlkh1SNElGtylKA9NOxiqwkcfDm3bIaxD0wwz79OHbAQ5M702TxcLMD9ohUkLTq
FpMNt5WSWb/iEuc6R2NCwXX+f5Z4C0VlfmN8kVfIIB0A60Nn1WXhNz6qMzA+V2O25fGtVKx8Wths
I+e8/AAUjLLdbP3SlQO1/exxMFkYnihZlpfMTfU+PNRLDlKYGVGNIJuiqt8wIIY8kUJQdkTVUYIH
PbYqYTeXnHyzJSMup9aCHrJZkPLCaXuOF7ZjJZiA+mQrpeKYtePdHXbqJKJaVZjV5HsqRn0xPEAU
l3lTeV9ACtd+HQIqfH296K4YAyVyeqZINJHmUE66RYMz4qtfupRMfW3s31PUeqHBYnnB2yXzaeIY
lSpGyNOulvkHJLi3x/MxAA62Q1f1bFf4hX7TB/qSckhBt4bhrH8FIcIc3cjRrE8UPH6ZzN8Ck2io
Tcz03I7JIe0n8tVMtq2aG35FTYae2AqrW0o7l7n9kl9gzv2ipTLrOME0owwxlRzFoXi+cb5kl7Si
5hIW8aOP1/c4jxkdnf9TUmHIPXr81Fgoq6qQxEVELmtRWMlt78ZvRIzOmiAxFli0J1KKXafmySLa
QiFtd8HShGOdwXc0Tf6viYArHrTB4PVqbR6GMQulC8mySE/yH0ypUirLwzr0yG3ydiKHkPEu5qxd
Y09A63hBkvF6YH/SuYn6Rau9VP3hnz9UAY4QXdObYJLlr8hAEFQ8n5LMBTnQliuFT2DkfBHq+dMb
dQQkNgq9jEZ372FERel9hhudZ5vqjkwWoiQgz3+apnukBgl8Rd+0F0HlOTcPie88LGIESw4BPOjO
VzTgBzrwmXrXhKZYMbba16asvO5F88zTAt27bW9kHyh+7mbjIfRNsgHFHpfZVZpDlYjU9cvqGDFJ
jhSVyEa6ADfuL0GAwPSsV5ktoFF1ZwEKwyqZDe5dySADZfQIQlzvpvox0YVON37YDqOtsScFf712
3r59VKnxGVxmz8um6nBdnQxiqSuYazolA/ZZBjCSnzYvzKrWn4hY26O/tURSDmYDsIChDtjP3b8m
2umQp2BueItsUWdSNs4NEqida0ckI+27M6uzYlph13zjJfcDbhH0hgadPsi9h5XqPniC+ngRmWUA
DxESWss95FWITX7dPyrJeuFY394/TgdZXdpZZ6EsGtK9rCS/zNF3lF5964w4XgkWsdku0ouSj+oV
R2bi9mj2xYtMs0AdSs2giO2rCPuoCnfiZc52+5EXr23Sv5+oFhx7tXa/2mdHFxuD2bb9YWP0ICpV
6+Np9WU7vi3u3XkbCoow7OuSPRsIVY4W5VMqkG0hrTkGpxh+evCD7tOGnDvpHvFuShSf3yatKaDX
jf6DyDqqHd3ZGulBsqi6RYQUE6qH5mqyft41lX+51yAzfr242/Wj3Yxb5NNgdJmHo5W5miJ7iBR6
Gjm88Sa1cz17BScuh9S2Fct64I8a81W0js/X5m8vCUriAT7rG5fFsO9S/zIcBRx4EIncHAHWn35u
l+SXyp3t4AqAY1hohnOF1vX0oCwulk3X+wJfRzglVQxIoTeeKIbe6MMchrv3G4GkXzJlbCENeHQi
d7wlZgFDLhhAEY3scyAjCkoIlhuiVZXj/46Zb9UA4kPJbqvk7zdCtm7Ri/iRHIoWouic8BLDNsXe
VgvyH28HwzkoYzwA/CexNFrMZ8D8PsrOfOabOVI78kZbbNPmky5b37NgXefHVRu7gCHbpHO7epVB
6C0qqOcBhAS87Q/a8zvPLTYmP6Re088JzcHb7jt1vkmk+Pbe+TU4fSWbAAsIHKK/86JtYXqwq5Yw
10vi6ZtfwgDG/hy9pog8bxj5x6bxgVY1sCRjEfdn0QRheNzOjpxVbetaSXQilEsC+bzyYlgi5BPr
Qn7nMTUOz4Qcrx7EFXLbrp2TDvBigKH0427Y/pPFoAn51Nq8XKzTUEEksHyPfpns8hhEyFYP8Omp
WXBKcu7teUDudEvi7cfhmSX/BfQG6dbQAEeLkhla9KMmaS1EDesGQ/W4zW7J1W/qCnu1bC0OI+r0
YVa0zUnGjxBvAvs6k9TSUC3Ny6+AGJt0veMGpkwKqeh7W/mAsdz7EoUZ+8hyhxfapxr8Lz1o6hAS
hsUX2wmbKUvCOlaomaVPcx578hJdwYjhb74uFqk2hAkPIwTOvZcEELEDMb4IOTNGnt8M5xcAcVD6
mh0IBuffDWjCO7o2iZBgIr9YPUQwQXnzHgFrskIS28ZxiwDH6P0gNigkz8j6dTe2YvvzkUEdUgoi
d3I5z5eeRNlEceHNSojh2XRyoRk48zBUZb2KY5VMvwPMW05M6Ilje+Lr32GMUiBasP+/vBcNJbFA
fCfv/gzkIvkUQsxqiPFOjXH5KdimjrkJhkCHlua0Kc6Rm8trLB4h7tZSXMgTNKluL0OBNaDoRjEG
F6VFbHcJgmOGXlmIj7CfCmiEe5m+hyZbI9cEXz6B0RaxHVNt+88m48NOuPDgjOFhlKdYlhW+ggeK
drYbhzQgT+XxOAuxZW4KbpZFkgwqSfQ+3XgV5iK2UD+1elDbUpNHctdgJaGUhIoDsmtYlIreofsT
s6uvr4jXiFl1U9Ze95ChV+gNS5vjHf2oHxVFY7b2RNZksprk1bRaH5CLPr57FYjiEUf6C6ldYb7G
tkkB5lovBSDd+GqQHngm+TOuiLYtRfW00IgwrXKEnUrS7yXZTnxYfFmMkNn0O64FcgQZj+Oie0d4
gkppuh/zYPWvi6tqSgmSqlPqubM3Heqg4reQrFO3lM4det4x7819QMU75x73ugdTXvLPVDP5NuDe
Bewp+72mkQIfNnX9K668as3WUJsYp6Y0JLl59il5caIMsOHfy6QaMRi6G26KwfWcJHoZetXxX6Wz
1I4KhktG4ErEXDvM+Z+H9VIgJ5UYgRfHTItCyauSy0KVvUpWnX1yKGGY30ssEuHEDdDKuWXP7f9D
UHJ/6h3Vyjr1201zpfksJhtG3CmKlQ677hyGLinAPfh+AGMbI2e1K5kKBSuJYtf7+Xlktxt77Ffi
Twe1WpvO4h11YFrt7/+33ABNrsjWbDWrIxunpVjIiEyxm54dyCigRx6MOEE7axq+bZsWgBpHAm1G
pr0288hJciyP/EekYN8Mxe/mpwUBa0/RJLUxM58gXkPXYpmMTTLJnglJR/RLH6PBBWQv+r6DpzGY
uwozEK0fllIFhH2El1WHxpGAn3sWgL1NLk4H5tFVuXHMeZor7EG/oyn6NIab/3Y4Lb0Ovjl2XF2Z
C1H5SBjtStDzO1KFZ7Sq5YoGO1YWcYr18PPUbyWMJGxOeg2GxJ3kDKl60W6YIsvWTbG9D41A7tx3
2BftzmaURv0V75wHjTd3PErzMyuwVzJ4hDo6c7Z2VUqpCEk3a2AfYGKM4NBZ39ErWv57F+am0hyt
iN+SDbJmP3RPMsaE4HSvPy7NCbeQ1ZwLnjIfgR04cpR8vEalK0QiH5s0uyQPMFcUFg7wECUaI+wk
QzlYAHDJJOKNtF0bMnZ16MCVg73brbAWoww/k+y0Fq/+j6Do6hSv7HoA/JQm0ENWxindPx+KSDuI
SAH3iuUt3p8j2FoICyW33zRvHIaeQZ3QUxnQM9+L5mtBPK8CvuCQJ2n1ukJkWZwNwayBUA4TyyHX
+raRbJ3uwEiSznboPkWxP2dpuye+yeLxawc6STm34f0HnTIj4vdg1xLxPFlX5Ec3qdUs+IyjSKNE
mhtHkVdyD/BBpnF/areHCam+Zd/flAxTA68DI8rj4uY47v1RHCUs2lyqSduxBrbG+UcDLLrhVot3
VzTY/5cl23KQ1EfQDLgzLXUDr2JLzswvTtAcHy2VO0GWfKSwR5U1SWYz0SvGrL390VowVYAaaHsH
I3LSa5ZT3cmoqXKmOB/0/yPibHig7/4ioyfhi/InKXab4TXWyJcU53yYLxAcE29O+fktiEmH0SPW
QA3r8O03j2MydnPtHhip6yV3Q3/ZkORCdJxlPtObWSpUInnxTo7MJ4n8sIdOzKgjn/51t8im7rZx
8+AlMgX73ErNu0FHjBbSWk3vLIcyVER6DphFn9dYwQ1emT49RtFy4r+85tZcx6HE+77Q1dXgO8Od
9EVp2k17UbndIG+2NNCqlBHvirv7LQHz9vOIgl7hU5A70lMdMaSWaFOdxd0NU8TJ4q9j9pySdDAC
NQ3ZCStjenIRvwALawooMnfAbtJbf/PLQyDG+aTWlrfJsJYbuKEOMVDtH/tHuOxjp63qlAE3kRxM
P0LXPtSKp2/t5FF8shyVedjnjXrmNBdsVC3FEZsdoLL6t6DWJnW3jF9GGLceaXu2N87P60nHj8Yc
dCjol5zZsswP4t8rU5zjU88mwvHwj9AQxGpZvVBeU4X8Dox3EQ3fAj45xJI8gzlMAUQY0/1gSOuD
yzFh00e5kgAYJ3VtakqAPzHGywKbYF3DDiwtKjau5oWpofPcoHya9Orrb/mNVRhRTs80I6s4RPx2
rYJWxJcBXXAGNlTKScO48tZMComJnJhADfc+i2n9Jz4ewmvR4IYZp8SzftMfHbbYnv05ENKyqqhD
c6wRtpV13xTwKZuOe0K+kZc8Km1qs5x6uzPt8UVG4bSjtw4xc7bhjf80J3GZYf4pmVO/6Mt9BOfQ
xGFW4cdKzrLF01pWY3onx53IFKnNaVRBJscXF73lHKgjcQQ49iMPY9LGyKOXLVw8k3YvjvwxaPI8
SjhPLjM1Sb1d0O47WMayp8Td0fvQRXtWTfaFiDuy274wByIkmRc/vidMaBiclnkzjfxw+4tlFdNL
gG2eo51feACBK2vMCZhcSmTMOs2TCFNBIzHRKYirNQmgUH3T5+QavRWViE9ja4qvz+6bnhjYJJIR
BYCDl4HgQALeY+vLalKoePXO0SxS+sA+ogSXGC2BDuvBUxCguC9PPgkysqMvrkZhBp0yHuMx5y9L
j5x0Z8t0hJUajy3lr6h6QLP+4W9iNIH+qMk/iFhmgNAHaoaDYOUrW0U9/po1FMD1rCeO3s9z9yyv
x1P2r+oXmLTFXZuWDcdDP2X8+JD4FLiKmzbthxk4BN/KDE3e6IXzLKpCfRvvCAxacNA7Nd3AxWOf
k0Nzi4lkWX8t8+tRCAxpGBV1h1QR58zHkBM1duA2u1mKffd9fb0J1oZhoYeOiknLyWFj24xvaT5Q
Q6PJsi2vhuQwsOJJGyCkVBkSlt1Mee/8Sjw8VemBHw9XqQGOPcaeSseNfKzrJ2UnOhxntsLskNQU
8q3qV20gQD62OZ8lwYiciEqHdc2B0Gx28+8ngZyFliSaEoDX1Q3F3+Cm7cSJYyWSLaYiFxtqsSf3
vA1AKOk5sUFVirV1ubrU7G5ufC/scQuFhgE7MKLFV4VpoQ1G/O6u3DKX+MMup2rABvIn8291SbcF
TGOs2f8goyD3ceHAd4p13Ro1quS3+f+ydkXBt6RRUVU6jTx2KKaR6QGNAwq6QEyVFNYB4JVOH9eU
vM/23SJ2i2nItpgSXR+NYznyiRaUXcmZ524w2M0i+E2RucAK2o70eE9kb+KX0Ank7o1vetYUXmiY
FL1DhFPg1VnxN7jtvsQFgvNcuWLkCh+wQuP17jmAzMWgLddk7h4U2EjOryHLpFSQfefJ5EqDn6OC
eqoVy+OR1zMZEM66JrqXxSmQUQa7kyfT9/Fyq+QtKAJ3QoWiM8Q8QTBRw4yq64XV4JhKgfQgevWC
xTw9wX1H3h+6ABVmDoQmi+Q7eZjhNZFMWFWgAEsWJhX6w7ovpzlow1Uozmal7gdPh++898/le6Tz
4iVLnCO0TewWzpHVDGOBCGyY5pW+6RB7VGV8pc/l2Gb7fAO1Bu7SCwOXTFJp3WbeMyMRfKV7CD8F
kExSD/RI0vhGK5S8Hoq3VZ1EaJVLhN9a9MkZcCAIBX/VzVTNXCSspfrlDwNG21ze+IU2Su9/2D/y
tggYaseCGXb12pRmyzQWMdcMjW7NDcb5b0a/pgJHq41itqHS3dfWqmuQ6hc+V/fio1xOYuadtU1t
ZDy2FWcVXh8hM68dUMRNZa0HscLb1e4tadaxGncjSEcLM9NKDVTsf7Ke97r5MIqXxEKASRKFnisb
DQE2ZcjsGGVQrKM6OfoSihDMt4Xe7Y9JsNBJq8u9nPvIWJ3nOB+22/TSshGuEi4LocmtrQgyaioZ
Kp0pGH+oQ/aq0VcMAmgeun2Lbn4D2WH0HqeX1AnizD3k1EDs9kuCu9yDJ3XsZtXXGzZ7wP894hDc
E1nMy48SmwaX4ybn9tSSYzM6YMcIZHFPHajEc1QYbEXX/jPIlIiYbTtuXlFE5XPjOxu2GWvtmmIP
w1uqlyX5JnAEjt8ZZfHKh/bdKMx+oZbTKPL+j1ND0NQGetYstOERCZeiILGu/0jfJ5cq+Xoewk8r
F1ls+OjFBnTMgjd0SAupIxAvhBFPJRNJ/hsp469GurXVzpsGJFpMuTaCaasqoCHuKPwQxVX+pBLx
SG7Oj45RwcJrG0SU7xU/kAjSODLayk2oqavsA8GOidNti1b6SiZsmYsfHyS11IvV21FvT8eB4XXD
XzLMng9mJNm6QrOkpDZ3DFTLunUFUxpDsIkgngKWfhlzgzHT1fvbWsPqcKOvHr6tQQZaVsX5cbsS
oopnatIzAPiS0hstiA5b6vRVAMnMw5BHb0LF/6FuvJCboa6l2kAPnNZGbGVi3VMFKqfxW5eoLhZo
zvy/PLEuoRsSUY1TV22naE/t4Kgesn/o4pesP8DkvRcFUmxJF18K2qNZDmyKn2RlINg/I+A6qAOx
MguR3oJ+ZhehHdGy+KzaY7+TDE628EY1JwTVPqUx4D7WQju/GTnw3zMCaP1PaXOJiTalaYk/2tsg
hFimQXXqMmC3H0F6XdiGivJey1fUR5PH+XcGWeD0CT6xBcgprB1keX+vQ75ZWGCX32daIx82IixY
q9tukA10AGaXNk//hGmbJcmZI9swgkjLcZrFCBwJasaYL1gw9GsIZnVzd15cbPyeeDC5PpQi+zvr
W2PxyiICxSwefxAs3N8zb32uQ/Zs3UcY8YvUieB5X87Wf4/vFErj6PozxIBKLvJrOPQMyN3kK5T9
sSycEYZpudW7MVfStLhvh5s3bSuMCvuOU3MLSkFCr2N7vIBOcReKJpfmiKvHyA8RebdCf3AuPiHJ
XJngBn/2QEbiO9ewps8pJjzbDA26f5GLg86Lm2hqnNGZtmT6n48USEFXpkmOPxidqL1tQ1ni1qrg
JzfJ282gW9ePkzygqwlqdpDJomlFzGG3UtoYV2YEP/XbKFrRKHcktVjVCJfUMM9TkjJMA3GoapeF
l89D6Hu1LiMHr+GBKWjAp1xYmW1i0iW30CxZ3e82kyFt4uk8Li8lhs1s5WMCpJrjJmza33lwMe42
Xs+gbrJpHYMIai9OmETmXZGqS3Uav6qP4eJE7qSlglr7ud6VuAn2l8mH8TIMmS+EdJVPccmLi2zj
CWmVWORt7DFY/bMRviZQiNbMa32Wob5f3D70XBAbmdLQhGDBL3cprwh+mC/+h4IBRnuQV36B4FVO
51xpSXuESdgX+r4kl5BV5eXF4cn/wpMWR1Z2LuR/j35vK2nBOPRxIDltmxuwRhvboEzC+TXUFEg9
gGXx2K9khJ1Jd4jJXWOqZ+gN1k9DKTH99MYuBOAEFr7Rv3qablHAwX/zbOi/peMH5Fefful43onV
BxnumcQCg0wNEuUWLTl6cNkjsoJJTO93btoJ1Ori17Fe2A6JTmaeXZb84uQLzzQJzw2UpxPG++Dm
30U456gH5dw9sv4TKHJFe9jEHN4dNkMUERDkCjNreY78FjyOPTxsrmwdNEKEjhSwmy+tWqoDtyQZ
ZRjFqbs4x13IGSMpyX6ghmlNXaSGyT/ZXX5DfMyPp6HQ+NuVmURJgFenqgRrzskhaqMg24dvK0we
Sz9/+8S6mS8/7xEsaozkvdM4pfIJhB3zS+ekO3KanHTyXMZ6+mkwyGoULPww0+az7NI4089yX92J
QQjb0/XW8n6srhuHVkP+Itq810BZxgY7m84PudEWsMjfQeV7VRT/UG8k68e8wPF61onq2dj5CJro
HZpvVNWgGmnLAiUPM/ImGAoF7AHGuufpWxvr5ZZj/MoIBkDhfhnkj4HsprPMoCigkoBXESqvH5qy
53Cw0+SADCJCz6sNcHgsKZPFb9tiqhJVDF45Y+uyKlFLi9nXMzhVzgi10nMW6dJI1TCWvSA2T1cd
BjHhGxGDeC/K29/V1jU2eRg0vMAEM4glwOAIFeEy+npV5SA+u/Z7lQ7uEBid54IMkDlymJ3T6Nrz
KzEZJlatzv84Ro1JFooQ43Eit7R/rsQwrCooGBS6c0MTmd5i8KBaR88Tevxp3EZtlfFJvJwX6qHa
rMFZyM/Jw98/kvscbgGLgbmtaO3t8mhLNX6jaZpehJPsjQOETk/6bZADzTiHDmzzZTplPBcEUmxB
gNVFqxC4LLtkBiKu8H9bOx66KKSL+HKbqKQLHFGb2cq3VZHEBWeEaC+Z5T772FwzGCGuMHHRI/2L
2TcZ/djxKWimVgFlT455ELOz9nb+TKvfNjh8OtSWEt4lDzNTIwblQP2TnmCEorJHdzMrXGWCF9dz
IxabrUZsdptNqCvsB/ZIQgk3/Z25ZezSACZi1IupHtwT23IOl3wRabWQbStHebVvW9rSHmgrSbiF
eDd98ZKv89EOEgZDr8lQonoo4K4KV1kY8PDpLE+H2fp/j/9/uAKOgFJ44wYy/MV9yjXkcZp1KpGW
JUf8Z1BZvLucDGLmVpIw9TPIbPdQ1sZyrzVebivIdQmim5U6fuN8+FFV+NNcipyyEoFF4xgUWhvm
a8RIPM3Xcnehs9Nwx5aawzpkeLSIO03JD0Rtiog9Xe7zvcmdIWmyhhBfCuEjOVOC3tlbZzPiJG/i
nD4bnCUTP9EoZL5rBZCvSOJHupSh99/zKDprsCEE9/NyYid2EW898x+kLRBaRMPTmWAweP2KxkgN
sGUHxn3SrMBge6JCABGE0kMIG5yUE4ihU9BqNd7uQCT+QZlMO7H0QZ2Rej1G2rCmMVzDGQgzwyln
eFBmQhQAlu/62eULZlY/U0wpiX6UxzKUdZMADbp3fRFGAoaL52gFNm293r8cWI95Qrb7y61irZe1
Fcp9iV5Y0w/kCZEwrhHIilREOgrYKa4+VCp5BtYx0IOUfJTaYRzwe+qVUh6hQCTr/h+SGNSoFYWS
P3Yp0toocwjbePYzxfxV3ESUy0uV43JwB89jA27LQUXRRAKUYAyuLm2Z8NtKX5DZbgFcDjMI731h
u/YKaQ/BaHkksL8ec8+5ATmfd8oJQd+3V44W+x71qVEP0EDBwTEcKvFovHtBi6G+PHGk9V2xUWVO
yzG7ySQlTAoKHFSQjBpKl+FJwXjFpU4EhDq8TiBJAmFj8Ph6S6/0mTBbo+CGCGt8jG38WUgwYNJk
OCMO4GP/CRfGPGzRXmrPpk0DXGaZ1gDfuKjRyVeppqeSlR1dWO0sNyNrVKw8HSISW52JTtIHQ0vX
D+nSQXlA2smBYySalPgE9YgPr97oPFlnNqBLOAu7AR30IRfuaN5V/2gw/cRMTukNbQa6BDe0NNWe
2emBV6vObg9V4BbQhS4ojWtnlqp03aKYpuB3tKPz+F/xFUrDxJ03HXGvgw0TzvUOcT6zVds0rzl9
lnk5YhBmCSX/lN6ZyYibculHNacd7LcfJ//r8MLDeK7vkRlAMRpsZy/oyAnPxugLzU6WkE+X5X3g
F89YGq2kSYH1exbCrqLJWXIdQCp/3jCV5mrCfrMV5XkDl9zSUFnwkV1mivzv07jND8T1af93vXoE
RHXkAzNiV3s408Nj3UYoXZginlgKnV1aMyO0I9RkQdYdPH1KRVAnyd2YbzeZCC/o9Hof6WBUbgEu
JSzXpbIMoma6bAMqwzkoDgKSJaN9HbdPuvTQvIW1cSdq6SwEfCh7Pc/JCxGKbLoS9j28tPlhhXS/
bY85OA0M1GWFUDW5puAatM1rGXULcAWAvJqH76KeWi0xjjR7UojVBItB5pRpvMCC/cGtsrPQ/B8n
5z6FJq7F1OOyFMsNcEiS1rshlulHgwYGkQkiYftyj406H0KF68cOU1105WX1BhseEv01gcq6McJe
Ashx7ceI2YKV5ATPVa1CCbNJYADS7B2qIGxliQf0ovt2uqW9dPVFhMxlwxaK/L2RVdHWzivorHuf
+j1V9u/GCbZo8AJ1hxpnfZNoVc9IdXC804ctsWf1cXGQ/P3ZlYdtOpm8GmTw64JfgLPSJJWHNGfb
s2Q5L7AyT3/kJcXItDyFr73rZjn7it8Z76WfkiDZLC7GPFOjhk6vIK+cc6DA40uQOFkXbtSlorUC
RX99XE7p3gWzgi1IYzst4aP0M/Ewxb5cWa1Al/klRNtsKPhXTTfRe7wMAn9RnHPggjwc926qiG1c
XKzNgbab8EQB/Wl2ghHPFJx+3oTihLD05SX/MsNJwtayMBJL7WncPyHE4y3uL6mPWv9Fsyn2mDOm
wlHigWWcaq7srGLZWqygfyd4vlfn6NfTy+sgX2NHC3Nz52L/A4UGm/WdCIsga0xyOD7gP6BmlG2/
KzOeezDKX8viysp11bEtwMIvzQec36SThkk5di3IiMPkVIw4xx36L7lDfW85VStePsy+q38V/bVM
jVWunwGUrYmIIY4srlXg71lK+6Nr9bLEKEK55Tpenfs1UkY8n+XZyn2jhBYMfEf0Tsz+WPxB6wj7
MJFuHyBXpGdqlOlQM64PfjI7zTaiwLU5E3OPRPdCMuSFSwmalgSHvodlbrFAWl5Cjp7Na15gEk3o
m91yvkeNGEKRkKtcyU2KqlaS5Oe3kQVZ+n/54eSA8sg8DRLT1Pia6NxfpqAexrmZ7BfFGxHrJsPA
UBiMJ5HRizT8klSrPWH3clQ29F1UEVBKn4N+vcCORqekrLafuugLRvTtS6yt/yLvt68o9sIv4QWJ
hOMsit/2hojzVGPwgN863F4OHzsKbVaWbqtevP1oYxaryS0m5s0suRB15KxQUIC4r3l5bIhaybAl
WxDVbVM+3hJk1VdA/snFAX7U3GW4Y9/Z+PdZHdM/HntFNF0Op3UF4xIYCYpPCeGl24lDsqiTBJ0G
aZfWlJCeRm5qslKV3rAtkpPwXnj7w/pMCuuDHAFxHX0Fy25dk4EBsaMopBXPVY8eapcKBGYWlsE7
FilacFw89cgU9kUHKUp5L5bN1tr+88PnTFK7BEZtyOqf4iGq9TSVwc+VrxF7Be/NFWYoQC4lh+dD
2HHNIife2YaSDyI/NtshFwgphzxFoDzhn+hOmxvgQmbMi2/ywKEaQUBtbAU4tkbb2G9EjWvqWjQ/
1UBpIOxS9VYhyTizBEOpqBybJ9X3tLrr9zGX2YZ8+rqLKbGwCWFu+3OMDIZKIKDG4usQjMVmf5rf
qbHh5LSkxzzSQF8xwg+lYI3REZtuNT3NSBL0r8s0tBBzj9LfmFNoDjnIpTBChS5Z9S4IauFlsPcB
mrzEMvm//1Qu8WCq1y1KJAoBkAtYYnOQzON6w2EcxNPCR4fZanIUwbeQdwr4kzvPZxyh+WbX/S8C
gjQgzYmvCwkNIoiCsXiMyN38b2ymCXb0pmYEPn5d/yhV4nuQgTW+v4cXgiMhXsF5A2iE41pVrGrt
1LZKIbHUK77K42Z5gLH3N9JcxWVa3p56b41nnlU37d85dAQicFPuLzrTjGEGb5TPxjKNlszlENZA
M1J8v9AJxqqi12t1wdRo5wlosncfG+zBmgNIzjRbPg7bvlVSzEOQ/SZXcAilSWnPZhvwPZBhqQv5
mEmylMWi8CCzYqwdOZiW+gHNS0kByZJpT87TrkO52+gWXG3W8xsm58urfV99bHnDuuuTNDF+mRvB
tppNiyMgxxQviQj44eHsyqqRMJE1K1W0SQirEWekLINuUflpmQ/Sx/iTVnj8iWrNnodAZQAf0yEK
cQv6ZqPNKtQgHdxxgRyVFeOqGKGZEVpLwkctIclVanChZ29+F5N7TU7FZwerET8LanXyZZgkQaUP
DEaIO15XEJkd1evCzFC1pbw13hpq6AJaSPl31LTmLBtBfp0Wqd7901Y50rIQ7U7usgrfE9X7cmEt
pISKMJnLRH6kghkprJEVwNDDYDqsjiUE2pqJGYpKH+om8D00WXSOI6ZUPmF9vwpmxjftvGLa/JbM
53D0uaKiFaxkfa4Th5nopYw6Ua0Woqg51DADRFIk+LPCQ26jtpLHPZQ0ikq/q6D/1mi8q0LoxlTv
SmZT9HkTcGlYsY+u3RXaBpJnjWPfgyIoArrUHOfLQGlHySrdgitw8/GwYLwb0Ga46iV08bLfjPEs
5KwW9vpL7xKXCytXppSQxIdaBKjP/UbVmG1e+y8edhVZUL3JC+RRxSgulAswA81tos5lnB4sh6oK
FWdFYSMrzPfHNpRAd7wOStxUeKkEPDf3+tkRa+Lpb8cN73MrvXQ8vZb/uoxtaARZc8m76y7HitW1
hYVt6r59bCMN+9bYzBdxqkeIaCMwc9eatkJIvXPpq70dNx/qTpW6S4hjKkk0wLKdt/ac8DcdKFEO
2b/1JnokOwl4aE8TD7c3m2xjDsDjI+/FNIoDDQT1/imFwzzDyya0TLuO3RbRrsW3Z6akYOj4KSDO
Hxw39+eSotKQE7NYCyufcmAPizDVwdam10YPA7csCFvpIo8y4pWf0SKD5Lc6SlyicGsnLqh4jG2Q
CXRoaq84xvPKFIKs9MOte1iJ3I2QXNwYLX1Rxp6VbSs5OrWZcGpQFjpv0LcG5mHQufaKm2gnZyXV
n/hFu/LhxvcuGDpV8WzryPcJwt2Eg+K8LILfiWSJh1TY7MMtAAuBaW5wSqvwpm+hbd5nTXKnIfPY
xEglsMqxYZVMw6sP1+VTBs5jQNCBzI/5plmHABVi1iww9/sxJdny4Mx+h6ezOzRoEwg7CEyxHPbZ
h1kPX9Dc4rY2jXcuXJGtBaHYI6lVffAILkLv54u5pMh27LTj2yJbu2VR6NUyuBTeOFH2lQYHJvmm
f5LJklUw5ZqYFEqbY88pFPQd7AnQEMruUWPlwJq7RnDIGASCmsdJQYvqcHa7lgxXQ25VS4gNRrBE
Qq6uqLvNrZtVSBttKmQ5+6/aqMwmoewp2lS3GVuY7pDu39wrkxT1junT748NP9SWYeoTv5K1ZDSB
k+dW1VZP5Km3tx84EsB3UcRWqb+AwJveqGzpYNVQqI9hkpsixiOK7MlWcX2JILgR427cY/Abxpsy
FGh/iboPLzawgmnbhzCqxE/ETZp0FGQJgRepCb/fEl9d2QZvkRJhho5o4ZH+CM3N8e3hbqcHWM6V
6mPql4HfqfWcP0g2ujtqbTS5nCQS5aJUfh/jNG/nEDw8kh88wVCaS3/OOmK4gp4juZ1akK3Lvjqr
yN5zPxtrm5nB1jokstMjPOGeoPHMnFWthmAVE2M41+a+2aC1qw5q+fCCziaEoODljRi1DMD3lblF
syKhPYyKel9VI5R4MgDPV2Cl4iqAecLudE6EAyXepK2jt3woTlbd7Y+9AEjI40QCSxNRmtdE54eE
xI8O2lQiXEt/A/3kfLW8pPHcbaX7pKl+DoWFbtECuTskUm5mbaZ3WhvegtuV1A8Dtod9AvpnRexB
3bQFmBn/GeuSOUjBRbtpX9wKyZNjjSxxdvvVsmK6363EhmjaJ7TGdizA2KDNPUTAoOMtrbXDd3ez
YRBzWwAUg8xozY0mR4H3oPBKb3RIRukEsvn3IsE1lm+37b8mSnMfVSQySnjzqYCgZArWyvR7R6nY
H/2X/x+xHuyXmJ6ph0xDcMrg9n5//T3YCglr8WL4eVs6YWLwjK4+sI+3mBzF8/UX0s56CNhQnDHZ
gq/OMa0LDoVeSwJ6Xs7QupSl42xIpGjA7NF7lPSa8IjyzN8p2y483YweeT0tUAtugvm5IaoSEuEQ
kVAhez1maVpTOz1+fRHJJKA2kkeS/SEEQylCGQwbIKRM02n8JZTmy5fv2OTdJukueyM4Kq63RE3/
Ndm/MDFDsMSzpiQo49bcDQtWaPL1wU7a9R58ASTvpS6pk4X5QV0gtzX7U68aoNjAwjMHr8QLpHIP
c0HUWVPjxP+hE8lStU0HTYJcL44ZRdR/FhZWCbnnEYWF5qPti7dCKcK0m/Csu+Qh82VGY1uv++3G
oLUAqJoY1hkP954SC6HMjiZiqXS1McntK5Rw3v2KgCny9WBMUrCd1/f2uai3YutjE3Kk8o0qNnOn
tMhezHwfKbBgaAi0D6HuGLgZo5aJXzwL237L2Gm2DmD3BwVlY+s/kroj0u1xvMtWwBby0OjMlRkX
5Q5BOMAc+gVXTn5MQwfVlKKlnrus2H8ZEFybPAdjZzP1dmo2S1cGKgrnXsKGHkFqmmAL3Ttabwc9
e2Y7SsMTGCh5xShNzZnsBENnNo6oUzcHM+dSYwbhMfH+4e4qtNbvY4tKVvEW7BNUO0zT1aU9OQ6x
4xcfUY0v+nPnDx9o5ka2AedmARSxad8WWBm+yLVPftNK8fLDlSwwwjGAtJlLCPtCiFroYKUJLacy
MLazKdMmZ0iDcFbSjXY3GF0rTfA2zdOXTNIDHVxwMv5NzPxYugtLFOjsPufRwOvIbZeRWyYtMN8g
boniuuVyKETy9Q22wQFyLiLunNc93USBc8MIYGdtb+OJ2qjhRD4xiMZ7KDT3I/wQecF0ov+WPKmk
w74U4zfnv3i/e9jgPlKaH1NSCkDZK34udaZila57xhxrI6tjmHacGVeXT1nWd1rL6cYQ/rDZpwvU
SAe/XB5mEeR1fsyw55jRIEmcOPiDcCsmW59GN9CyQG1QagIx7jkOOi4RVLFJ3HI8iOdwgfAU7BtI
ogPwADkebaNQUt4SaX6CZK7dMXsVVYVV4hD7d1a/c34Chj2QDj2GBO3UQA9lu+3Z/i/9oCjVrc86
gzRZqSwoBabKwan46IRDzYM52dc5jx6iq3J0JkgDMD21nFFZYTSURsfIhDA/F6PEimHg3I45zLoN
3AiaokoKFjyz8SGxgoO1PLzZiyenr5SPMus0xbH7nfeT7jahZrTlGPCSU8VRYgYfSVn+2A6bW6w2
BQKJ3poPBa4ZSTqXSnd/F+LI0IrnBesM4Kv0G4SEiVzxVd3Jek7H18aVCytbY++bFL0Dxa/1bZ/f
xOCfmjMgONagvpG0xT+lbZUsAMpBt+DwjaS1kYbuHUq8uRyGoHTugIFZJ3C/OWfH0ppWmYGkYoPH
Bh75Z1HoMgw04VgYilA13eYFu27X0zrJm7zbBCkeYHTJ3l4DbYbao//+zz8bPK/gCaL2ehxMRfiq
M+o6DWuZb6K1sqDUREaMIu4NCUTjWvo1OBYn5J4U4/JEe2TgMzfTqvxCweyZs7weqsWEkwmjapM1
cCfcF0I5yMEeQzBcD6d2kK7/yQWE1PPyJUe2pRA5cGdZ5bchpirHXvzHwdFPhwQfL0LmSICoyu50
Dw2hsaCYihjg+cVuLhQl17CrlMj2nRg+cbHr6vBtlXyV/ZLv3WaueZwX6NH0b6LZz45nqqwu3nAl
WZQ8qKTBMUFZMys8aawE3dqqjrQDsuXoXLJ+FV/QtItU7oyb6f6N67zFd2u7anzr9DXuWknfn3Rw
QU3AJImPa7UBZC+J7ZQHmFCKn9gS8sidL0XfxcGIWBHrAkq+Im0/7MugOSwVZbUcj4taA+2ol2RK
Y9to5vTfy19RwjE1uLScAWlNiW33kwcTYvZCGvsPrn8KG3k6iXR4yLGo1V08Ss0gglhM1SKQJ9A7
dYLuBQnJO6BCs4Ng8bPWr9FQFcAPiiOkfyhxNxmdF/hocRP5YSPng0ylKUK2vsESWPt0zzaRD/h3
B4K5gdKjYDTFGSlp9m0fE+losSBozFcbHbcfdwSUlbFcY3oqFu3OaTduIebxGv2Zulm0s02To5OS
+A6aemc29XS3xs/eaNwb0F1f4RFZZTfxn9o5xWrJYMcrsna/JR1on++Um1ItfiKT9dnCa0fZXd2Y
owhLOEN9GDg+hl/YrZ1h9GqOCrXjyjg1Ymn2XQRQEQoazbiEsYZp3iIhIhHTWSZwm1Cp9zAbONZx
8z2xaDIosUNSwBB2mSK02p4zIeGTh+DQWd9oJIC/mmRf+hJ63TT2rHYQqpY/6d+a0vF2AbEYaQyN
XIh0uNZrk22w2BfUxlz/WAdeNSWawf+Eck3MgUOXhhorZKniFbyac9ySzGUaCMVmsmfD6QfkrWUj
SusCknS1kY3uQhFQquP7ZQiWlTANRmO6mYBLW0ZhwAmT78P2XVajUhBuGSFNTtUpPm3AfPJEx1LX
tU0KOTWagL4Uu2h3Lf9S2ICFRuNnubj+ubyiD51xHTHolmT11q+kGkROhJANlkwOe79BKQyN55aF
uCH93d65hW9E99AJMzRgepp+W5jJxAWp91k0T94zdOHxbErDLCIVkabj8NWzro1crcGAXHxbz3yc
j40wDGTPCMMbUe0d31iZQCgzoQfXo02ZmXic0buonbuccomFaESAXwuLwRbea6sThz/wnOOiU/4i
qh5U89zTg4UwhBX6g0+rh43iBDMys8YhlScjh3T1HzTN9YUVOgcnjmghyzkQX0vE92zbXoUyfgW4
vwN8OYTtnHHsLb4OGr97K5Medsmr+s88E2bQwgld5f3671aLGgmOvRZ7lbjpCmjOPTUz/fWnsR1U
cgiM3Zp8ElfeytHovlAYWPTJelN7ItrQXxKo5d67wkGDRLpzSX3t70UWnheovf1zmxl77yIyRaCD
tt1frXp7MpSJdWi1LkYWcF7W0VdZO27Rpc4gjJEARLzBjsf0UhRBbq7GOgeYtBVol5qD0WjSYeL3
KkRjKW+DhGgDN5fBBm+LNO1PGEQqN3MQjlPuy/7I1ICccLjFnMlu25sFXxTKD4qV6cYOstOCeFdI
0PP8AxJ7HWbArxH+9NfSH/VYDoB3SWlyvuolk6EGUUiDgbncCZ3trfmGY4OSx4Ank9UhVyyhtYRF
DhXi3WmWS1sddvD8OdgXBcVUv8PFJjFByfh0pYq8XYRKo8flMW6oM/casKqrQn6lCFAUxa9B7uAk
P20DvJxatI/aQkNSvYJkez4t50h0erhpwmoEtGNrF+OA4gjYTyYCdHxKEPLZmU1sFgZSzgXiTlqR
DsTfvRSexrT4rlanO+xnJ5wScykmhBraXEigUWzXTXb6K2qcSvHm8G2BaxdR0qXhpavZN0lX0Wsb
Lo/jXtlnbhkElwMPXVxRL8xoIcWKI3GZsYv7FWgTWqpm8qn668as6dlcz1EjOVUFy/2hujKgpDq6
KGR5IyX/XjM/bqQ36JwnwhOmVtwq9E7BuZMCAvsbv+OdpP/YDrUiH1k7/wspBL+efYW2dzYR2Dwi
SbB2EV+q0vkAVQQIl2N4tBOTdLKQ05qkM2xlbwsWGPbbdWOn2nfO7Q80vVhESE1MPZgC5ZOyTQEg
Zz7IFbuNjBhRYOOHkTwiuGaqP9D16Vu/NjYFEbAHA4ItSzkz8AaQ29I9FmYZdG9DCwSyP6FGfdvh
TrlzfNbREHUAcgv3oA+mZPJ72sBU9oMz6y3nmiAzLI7tYTa2g9hRv9hpkWMRkZgtAdr221EtsrXi
EqTdhjwhlEXnFOXMe058yY7b/45R5Nqu3ieSGs/k2M5svS0sQkCMdJkrf89aB9cmbdNfo1GO7LOI
IXoDHvZhsgjPsozn1fXY75lmq/1uHW4W3MzJVONX7lKIJaAw4P0BNOHsLN7XTp+8t8K/Eek73w6y
YDMoSahrBcHk7B8S7VLI+LPpOHfajQThNKRG9VWqUdcf6U0jJuJiI4OY9+wcqypbodJLdRYtuV3F
Xum9WSMTJEBlOFNhcktbe3IabawaWVRaY00B07DnzNGtrRsEzF8A8i31yhOV4DNNFbaDbrgLElun
FqatsvksfTSGs3j9NVQpoVuALL6yi2SWxYo/n5KPAWdexbPj7peheBo3v68JCpfaXReEsStSFL2F
g8FRi47kJD6t/OxxXShO1iZgJNXRQmdlaP4LRTUYU49KczQbIC11tik9qN3VLJVXHnz9GSP4ycQM
d8wYy9mciwXVNxduWU1Xv0Cyppia03m4xwIQGO7fb9S7CwDYjh0o7j3TN7A6TcX03XlA+iBBFnHj
PCr3W1m4FoeXFVQH1buzEkg57+HdZdLAzjw4TJFvFlQYUBsstloJp67rjl8hEcP07bDGL+lmVtN3
CLaDohztqSsmhpJB8MCZWnDl1jHdpF3xVvX/hU9D34CbwE/RJls5AesjXS5mYAx+6fx5123Af5ve
oANxrO6S4gIb+qAOgjn1w0X7NL6KrihJ5l18pPasNETkkTCYQxQ4Cw1xwIcst2fI3pV38b+7MQL0
Q9GbLsvrgKNRKMge9RPa3UcgUSkMl+4x+3whb0c0LY54yUUUcO5NnMZEvBSqC8tvUiNdeW5uOreQ
05iHfVIWm3wgos9PZaS13UNQONkfH3F69DcCpYHmFYCrllsSxSaCkFhU14gWqNf2jNQLj7KBAQkJ
PQbp/nbrpK2H4WGarWEpoI4zuIxAZSWc3XMjCdFFBECc6pBnq+aXn/dKQphCPCr7lclqEIsL/2vb
6v20ifVzQMNOKvWNJ3Voux22fOFxPI5pTb/UUY+sWdFLvB/G78AL8ScDbMOBVQ681Z7O7RWtqaB5
298nYp2R9x1IL0bYRe/MABP1W9lOVL/zI4tzTGVohg352AhDNjnhj9VW80ur3326uTJ66CqATw3t
fJUXnWJe51m+9I4IB3xFrJpfEH6GdPWna/ErcXIL6Jvg3z0zNhrm/ZoSRuZW1SWVE36xzS8gkzfE
ImGbHTetk5djVN1kIGnWRFYZ4VdvJpaqTiN8nEQXpg13uE4rASgSmrj4Dtymxnr898hjsnuOZ8bf
3SFSP843JrRD0AUvr10dR/QdudkpiMYe7sZYEuaJ9eMzpBzqkfWpfeHIxJGVnpwfAdlN25d+XBHE
3lrzTT9zWA9su9Uy3vnU3rzRUyK6ujue8VwUcScqTnj6zDQPl6bld3Nr3EWYyCU+sYxL6JByfQDE
hhjGOg4AkpmVNyurtmDWh+WtPqLpu/cDyZ4zQQoVIUCY0+wLmErlXQJEf6jg+xO+73Gjl7/2JOvk
5OItIqLt4vvJh3dvb9GEh8GEpLYJFn6XJB7QkZbKJ59ZQ0nqHPO+jiozFnSeM1R4Lw8/KwujfuGX
Nnd/pZOFtkUHL0Jpd5/UWxU97kHmhqEVxysi3cLAZMo+3sEGm9IaZ707KBwxZ55jBtwJ1Fqr6UCV
KuZS2zCwMDO2QHSznE76hG61dLUUMFVT0IX5yuZhz+QoXhNZGmjK1vEhf3Ya3sFnZ38ANEPtoBIm
93M6RZHwvEXmo0SrbA8lF6Hrnguo3mxt7uCWI58y1xHY0fUu0mF+Nw19dwqMOi+wZ5+XE8+s51Du
7t7vwO0c+JEHbIjYeGjVwj9F1XAVnQIVfCSrbngcshXYFPVp5a3jPsmXDVhJNqm+wPg7F8pExh10
RbFMXLQLwPbYU4aMykNFV+EKK+4jVrfbG54erG9ffegV0e6S4CJmIhbiEGDya1OJfZrXlQHUu0np
NE4OBwx3eluVpkDj9DHJT/L3tSmVfFnHcrlOodG9PnmeG2iu37wq4e2QOWzkYoMkPZI6E+DdrJjv
0KGsX33RmFHbUmq0534E8NM6f5q0SZDr1iW29JzYOteFUfUljR6WEcwplkcuuf9KzFn0IBMCJ1R4
c3bODAS8tuetxuX+pRWBfe9zaaak9o0YyrAhqwsN3xbA2HHIeYDpU+xSQHnui2qfwLmd2ZXN+JXV
vINSQBEUVDYVECSTn8p+fExjB/WxmK/FhJBJr9g6tv4obzs6EVBlCW/vE2GMAAm36WstjL17ITv9
mJnx57+rEQ3+yatcezKNZ9v4UE1v1VgkYzlBcTY/o6PlpQAhbmdBj1bVqS0niP6dKDxEbwFewiq3
raEtC1VtPZ/LTNaa3GU01axDN5acNSb3Zd7AZlQWYEy0vaPLcvO5h7uudMrsclIml7MZ2CeoI/Lx
X7GEG5uw2GWh568epwFAfAo2c6I4AKnMzKSDz47T8CvJcXuZuGQzLCQaibyqw7b39z1/3n0HA+8s
DNkUCcJZZwOAzpE4QE3/Q757EsWdF9UHk8rHWf1uuC169V1A8kH7kB36RhIGqhoc+D92NIHqgXfG
waikkyYtL3Q8BGXO/Rn4tob6EDPg2lII1oOJT1FWOfJfN0mD2TFYKj9z8a1etm5wYZKnftBPHI6f
9CCWJK8cIT2LF+JI0GMv0D4qnd0RcjJVrzbd7uAeFuQtYtGMyK+NlD69k0EEcdZegbvwJF93knq/
KQ9khQWU/DssV7QX7k/pZroHemIEg+7U5YOJxJp7vn/MNRlCCjG99eYpTsnt57mLyxzg4qGvURmw
4be0uql1niz5JCihySu1nCAWFZXhnXjGL416sVBoyFF1Zdn4PXPXbRZGQbERwzhro9r53p8Ad7YQ
NR5p4GAV0i16Ps1uU6wyT37+sWchrEBBgRrzWKXtcZKzSeAfqyssTtCwBdpqbS8fjFtJ91eoXtOe
KBvU/HDTVXFMdeg8xR8FwNkQpnfidDk99+NA9iueyMKZzrkCe7/Ej2Gk9hMk5zUsMe6SyIXVX6rJ
fzCpC+B2IjUke0AhC2DpXgzdD+Xurprr8GiteOxM9SNE4jNaIMAmQjGIb6aOYXTLSbSVJ9Gz6K0k
Wr8qQ4NLyokgnH6GQWMinYnG67/ZQ1DDi/W07JbfSF769lWvUHEE0g8ba+KiXom8TVcKT1RQCtg0
60UOWOcYumDc1Eeni/SHCxhEGvHALcWGD5aiTWmFC5d9dKSLZnTowtVKk7UTjCHYm4rchal4dVQj
x2W3FCN6XFX9tmGwqXQks2CHB1J7E5hePUPsmSvcarKqhd4cW56nxhoMODEn2HzeFjfjyqVglJ+j
gHM8sGD0l/QDvoaH8+bZLt0pHSG6ZuEvsqXWoALi3/SEMNqlsb58ZX5hT1pph9ECbhbNh/hnXRRe
pQ59QuXmKgO1YHcXbjBMIJjalODa5XZ8W+yUMDQg789pjaj9Q8tWiQJc2jcn9s5J1U9tqBjac+Bz
WNSwxNT9trw3oZyoGip84uCyyrecpvoESuQHfTxzZZYwvTjHysRXYV7LqBHA2UQkDmqro+yzbGG0
EuRETZ/1Wz3OkPFhGpl2d9WIpcWJkBnWpFLdpn83GgP9N/kHZYDRUGw6m4Z2onohvJz95nsWfhlK
q7swREt/KHc0gSSLRDEroCVf2l0jNJIR5B1C8e0Xmammvmy31AI8S6On6FyM31qsAUfsmggzVvJP
AjUK/+ZMzK36Pp5aI1Q6UE3WpXLwKAmHfoDT6w7mMmzSsaEd3JsYK4yef4MCoKnqGSDnm53487M7
DX3iw/RY9Pr2fbbKEO+x24xMnNnJz860//CPsm6C8wSsFr5vR7Yg6GNzLMFCftKLvPX1dCR44RWm
Oe4oYGOguqCZc2pCLCfHi/NTrUUW4nclJSNBexkb8hXfJ2uwIryFOfGvAgCqLckMpKPfmBQIZ65f
Idn6jt1geF4NOitAm0H71VO4DrDktoRQElanBTaLpirbwMsppqG7lpOThqjMlMSfg6XyDabGABs7
gu0pfcjcUKQTCpPEEgW+X6YjUiHVJcRjT0AG8QZH+9j0t0gUZa9Q4Uf89FsJYdW5EOjYeNyF9yr5
lVPNCnX3Dw44mZl4kHsy6BgW5DYC22OKZnuexkDbOk6DHzzujKnk+Gx7qIG1+fVtaA6/Z6tfEAs5
uF9Eo5K1iY8qkzCSkQ5uuDydKJIPhkVk8EZtrLW0IcZ0JoflNLaC3t6xRZAwLLCLNqoCDoNfUwWr
Dge0MsNl07aVrLWE0pBmdeIapzZMrFI6tEuyXQmoELBsMIlgc1jNrnNDGCpNSrasJGtSgCbHvjjm
jhbFIIf+wfvzVeAf/muqBapFFwvuINyu5O2zrE+tlgfYAdNMAQtKH3/+UfrKvx+9zvn5qZWStCJ3
ecKhaF9vpe7UN+RB0cSqdO2xoHk16scTE6So+6fXBR78+n1Z+kjMfiXJfUTJTD74rgc+fWhtLyyb
6N9LpuZXxN3KT3Lt3vXCqOFYwTQhh2ynci9lEQ29F9LA2WVOyA79V9sf9jjA6stLdAppngnIwdcE
XH0qHGsrKkGoh/O+peEYsVDNXz5p6SrM5sKUVrQG6hSwShzB6BFpjBsit7MHcE/KeYrmYJMEUyxp
DUl8/pEGpaet/Xe8cyE5gV42iq/m8wCiZcw+PUwxXWiwBLyT4LuyJSXw/WyEy4s0lc7MViO5Clgd
RJJCgsK35OSkXwUKtTQ16fG5gew9anjRnYSSQ0chc8IQKiJ9xMZK4XHx5XouPKEV5pQLH8847yAM
CdFRgCey/NhL7vnx2o5IM0Ng06x+vlpx6ImpEJoY/gWY1BQPvTe4UrTV6IsI4PNmM20mg8VMOcFH
RvMOj6P3qM0/siuMTQZID3kRILRvknPyi+HrsRD8VwL9TPVgUHuxKCO/1iu6Az5v31hhj3kaTYC/
0+ebhBDtcZlZu0c0InR9cbqKi8nX0oMA4LJjU+5lg8rVefooFPzLyG9GDn/vaNv4BAx5cf/dx5Uw
V0or4todjtsyqPgiYGxIKjddYiViJX2QSMqoMG6RQHtjFFHwNqQB86gq8YBno23WWHUlOIjGEiob
ERFmJIZ5bPbVxlI9KZahfMdBan0eEmnNj+4K6rqzjOKcm4cCT8bsPDFDhKce1jHeFM6Qub3kGCtA
CLh/H09OYYgkti4fwkJP0QB0QO2U3RQ0K9jYiDXO4kzYT8PaHHhjRGChqT1Zf2RyEjly/9O8OK1T
b4JpFs8dMRawrOD9FPapTFgxHvQPtU2rTjifZhzxwk+m7HboG7U/ZxP393cnXp8Ua5ZbKlXtQTnd
G0p3a6c48liIQO94tEQ7zJECbEQpawBnBZ/icGtout0HB7993Dd7Ft2uRlXmaOZ0YpnnlJtv1BUp
mcvvH3TFaHWyWgFH1wxtI17QFhVdsVeXPTJNX9tcskxt7kW5zpHbEpzDHcmdKTrqjflBF/M9rD8o
byswRPLaWRiKPmM5F3M5K5/o5foRWW88PAOT+IkF7UkvH/Cugj6Z6vgD2z/G+KHEP8aL16A6OCJZ
EVhqCNGusHj1PChH+Wpz+0FPQPVlv6MGGggNwSTUa/C4i7tjUl2NRupxALH90KkAGMISMwBXSpCO
FZr5OenfILgOlcqxVm+W+P7+oC2Ax8czFUzfJxCrAOkoSZ3l1WbMPnIP4gXR4TYUc5LxwFBveO1a
SFlR4OFE9KNrnK/2riNFoZWJWrTVYlZwjEnpKXl1iZz81rfnMlzMWNJnS5GJMk2CfSnCUcZkVYXi
3ftflKbZ94qqW0dKDIR+WWZHyBONhOE+3NZq7ho7eOwnJm3J/4fKqLtvJ4R/PsQX9aJOvol3LrhX
JOLByIBzsQ74JZOGduKoqq9S0rpTz2Vewz/K3HxgGAQJ86FTVzLe/YPznI48WELBcmaS9iaJCpx0
UoxjI7IVUT+Lht4dFURHC8sAbCXPz+dp3LIsYY4Toxnjo+J1qTR53O4FELB04HElkrFwxmniXE3P
6eBRmUxUpnqTn03qm+qMUgcJ2cbGOQMJetMKPShi7u9dbimfvD3ZiNrFwNoHwVam25ITZYDcxUaS
8sSn1MZWW5C7VykFqdPxsLi38yssyttN0hn5qTOTlQ442/c6eD92aQDU5enn9LshWn10Sf6T54uR
z6Ae/0/cAMdl52M0iLwtaGUQi6GsusoDAfnzPKeu3tC/ViEaIQFDhAgs8+7I3Wy8wqtD4bkVo5VK
QP3nkxxKN8PdDdFfI45QFJv1N/MoPks7mnhFfGMMqlgXgcZXG38lAEWS38totIusD1e8Oh6iFitE
r0YzsLdeqwHsGKR0+ZDxOoM27/BddMtbGbLNI2vZPSP2n5fIPN4417wWVuEWg8+DJoJtVLCx0909
3crisGh4rwJvO7A/gkcNelCv3XW3AsqSMFK7pYUX5G2qaFzo3kXKaA1y1jZXrcyc2L2al8krNEgf
TChwS+IpmRCGu2uD7C+bd5Ht/+bkM5oZiuwlWDRIhCUsBXwuDBXlL0zDfQWMUpsosNl4qsSO8B3O
oxEW11uAL2sd4SR2F/vJRVhjdEiqdtG2EYsm3K61m/SVK3mcGSyYcc2mMLzuBl2SAN5LbFCGZBiy
IlPbsVKAnGFHg9PDbCd8Aw8J+dRUNJbs3ATpmBwnlJIP+PojjI3L4aZDnHKPaogzLRCgzb/uDDvN
Uus3TDyH3behaXLZR+MQxldO2aM46yAhTlf47VpCWID8T9y88py6D1s8uMS8mIbo+ATBstkF6IPc
Vya0INke3wUqw9a6QcKmBwGbnIfs2JKtHFosFU3xU4cyEZRYblN7WXxFzSaUY0q+ob/8cq9L4Ofz
EzxvgC+/xZq1KTqUS/sogFkurH66wegetqL+e+NLOynlevEA1Ykz9It1bNL3gTAmKCcIfnFYDlbO
s4oSr0hf/Bq0wWJ0sj47QwSVxp6wcw9AVTki8JRZvbQzlOZ6hlKE6OMOo5k3LGMXPI53ALQGWbMm
ofL03Zqwf2KQiOyaqU4eGEjx+XHZgUfaXV8yIgW4/gVWKayR1bQaLkviG3JRXx5k2+OLOA1z4hIE
b4dPmSuW0tXCvw/9/SZTBwKhxIdSDeyAp+daPOY+vmPu2XGISE0c/1jXRj/f0fFZ2vsWJapMyNU0
gd9X5J4hshZNIQHptvp7fWIzAnktzefntGHZjg49pjgHO4uIdxH2/Y6swUQeGdIwoifwWVUuub9x
R1ctHng5ADIyYhneqZr5eOhJFhS5ZNjA40ziGtVKxbQ+WMrmCK3brXTMQqckCqac9SFma62GYLgP
w2PYJEVBvDpDgJXpWkYOrOfVyMEPMEZfqANS/aWlpXPZZw2yinVv9PmcXK0pjpkEFIT4ClSJnMeB
g/IEkiK7dkdRQHtd8BAGti72h42Mr6oCsCZdpKlJb4ZVbkto7Ok4ptB1NlexnNF/BlFN8U+HLJOd
3upUNC5orQB5Mdv1ovKyi5QdT8b8DY4gLHFDe5f8QTHonZzqEAhdIv3bwCURxp5UvmYYyFvDTvoq
zJUyDqFzfLzkBPtwebQoGrYfKNy9PdMAyXiBnU2HM1BwSGtdlkK9JG4TQ/FO8yAmSH4lbQqHunTO
/X3nD9tGWO7TopmB/fnUM/has0bCnbHMvaSpvHP58nqmj3xs8EIi6JG+w+Q10nbksEWVr7xp/k7V
91BljDM13SZENyPyuVmRnQrFErHUv/2UMtRiRCfQDrlrMDvJlQ9OrYBmZbHZMiPpjfqZaY2j27nm
GkBziGWgKfHkyHrutri6MGoq43aLyO87rMBtblbCUoOtPnfJgi7F29uXQrkFIimUcI6NsCVKPFg8
IbiF3dE9d3GtcZtLBDBA4LTj/C3kKmHk1Xko16+3JPnUG7Sngigs1BOnDXoyhZUVX7n+nGCyfk4+
yznO4gDExYunQ9AA1OolA0Sh3qzUIEll6hACxfOlTK0TtDrC+VvuDG2Io9i1XVJkq02sPIuGUoAY
VylKOPiKvPbyBqoD3JQn0OAFymIKxbXEj3TVr3IQmWsa9y91Kotso1JtGZiM2TPYgt8tS1cqVr5V
GA17/Ca5Lv3l69dQDVlFdHxxSG5Fjjaoxu/n5ISuEp57ziNwO2s7vtalozYecdxE/gvrzhEKt+3m
3rUDRK5aW+3Edv1oZssSCk80KI1xQCD5xlKX+gMi6oXNxOxJXMv1jdQALLiF2b5wQoa9Rrbj6Izi
SgTJV8haJ4em6BHCpZORcAx9QyTPlt5CmRMTEyb8Xv4azj8N7+8RGvSL3TckmlsXHDYJ4UY4ySRo
vWfJIdKU1EBokn3qgfAOTquO2wK56SiFqIrZS8vXD58hwtJ4ZnwB8ceuS8xQ2OrCNHimpbfc9rV3
e9ZySCwOodjczX5fNIMwqlUNeUHnWoQaQuIvNsdoHod2S4XxLTc8UKq/TA94NOVoLbiuj4qOA2R0
cmAq3kUFGlitSx1hVPHT45xhq1Y3pR8wePyVGinMU1uYtAD7DfEeXdc8qXiCrcXCsbYnAMWRqkEV
3sf3x2PYu9R2JVhgCdKmnrF6GZsRdPHlMYV4Bt6LsnuHojGrTEJkYLRYGbjQMb9FueCNI+UNHDJA
tCzgjLwI3hm/OxaOMNOIGWe9u5zoBQuBsPPzOdqh+ahGacUQpGM+kXDcfQYPGdJeu1+gU9TJgJ/i
3esDWWMEEeeZr7wWJD4Krwj/HgeGwaV2LxsF0JsBvWNRry+p/gOiIMvPqxg8l94efp2WkFdB5dl0
jZhgYhbvEoV+QiqNRR0Fs6UdUqnBaTbrIo/TUk92wzzzuJYjArtVIP2JoT3srYqHnu5VurLo0scc
tT+lE8N+woYahzvaJr0WnwpwLCrfUrqy03lvdexDtMm9bozPORr55nHK5y8fm9zPFUjGjM/lptDG
kSbBCvhQJfMPd036Q+Y+PZdIdiaDjFG18dXZgtu1cBEd4tSwnqjNw+W+k3sPAESNY+ZwKIcsw7Nt
g/4NO312MEsYAsWaozXYsOnYvdZ//6uX43nYm9VGgV4FeIgntLee+iNwHftuzYzcyTN2Sg9rfP2h
Z1Douu+Hk7KyUkB1rWim9CXxsxdNUuEQ58SH6KlcU2DciLW6Fd6Ouj7j6cp4TLD/n7llD3Lk2lIS
8XPCe7zILIRkq7NaaOccd4qzOLGFrcgYhGoR3gDZpXq0CiZRKOx8xUaDve45sNbAE1FNMsKof4Ev
39RY5jhv/OJnDqhG5LiMJ+T6dPSpVjbfpG4bAXr/N9zmJGsTQayPOFXHGFhQwRR3u/B1ztrGaWJS
bGICuCPLijZRZLyVWmnTrxyk2h6cWxIhnPJkJ4iktjdzKQwmtmQYRQ1qSpsMLJnsdxQGNcBEnxGt
PeXNCxMAaV61ThNIj94cUPp5jjOTb2KMpYMoi7VsfS9wML4lwmr1ANdwAKHO+fou/5RO2j2Kbboh
PmqPf8k5+YoXOR1TsixeTEGxmY9l8KsLj0Cv5dagkqm7iTgakYfPg7wb02Q0yhM8pL/F93rQeqja
Q0UttDaCIWYSth9eoTdna9kLh0z8Kr7Fjxl182vcoCK01cm3YBI6M2qY2RYBFI7apnbDorapCUwV
c+EX1yypyXxZlfdqANbzcmmQpYjMGvQX9fifVBce0DisLdbln/8NFvxaYf+1uSA/j117J25z+gYb
axrLYiX+z7ggqqU/ZnsV96xCTcJMJvRKJhNC9dp6Np+MbfkSPRtcBdmCRLOJSrmIF/k8uIVs15l/
kMiiHv7bRWL4/vRjx6XGUELff6a2JGGPDBLynYjbziTRzb87T2QVf0o1FAm1i1vEQaGegNwEYSOo
vk5a4u1ujMQkaDzueT+lqay5tYjrFlhvPBUTpo8N/zQdZTVby7/5Om8yqHWu+UUhmpGq8osAHyOg
Sa5LOJSZuI452K48USxLaI7c9SDRCSD7Lly8ccTt77VBdIM8RVoZUiec3Z5/OKvFZ1hqlvg/K9/m
HqwM3DXYBNhqqL7ia8hXOG2kk1ZeWnDE9qrta0BrN8ggYrceZlqexEY4qXE1tR8vm9iU/g9r0oFY
5oNWCg43w9MevY28BnzYZTPix+vZgwHiAit/JD+JAILzyvA2xRiugNiYCA+mwcojiLjnnoTmA/ky
4p25bCtC6GRcYCK5eS/rM3RazsH7pXafv/S2ku77mE33c7afMWyN7bQ6oE4fghefw9+uCq40mMs/
fpUWgKulG8tFPlYurH/pmvlWP2hWu6oS5EVxg4XNKO9DnZHu9ujuFg7fFcSLhXfQF7xmFc7SXuJd
7f7h+nXCQu8dHWlyQ7qi58OibDpadK9n2OVyE1C6Qpyg8a8b9a+954ILa/yVXzCNC/9mxypSdNoM
kd+wOgY1REpKysbn7QFyrsWPjmHmKUl0jRakXrvruU7Xxx1Dejxs5BjAayNfuvvRROQDPbnH9eMh
CTdw2IKrQ7B6GP+XQsPEyQwyr7knqOh5h5Pthnc4YrHGOOtRi8JGBLEjMPvtZHJGWOMoiOwh/6Wp
cWGSsbEoGYwCxduypFK/M/77xhiK7ChwIvzFgx3d/00IHMSNiCM/FXAaL63nhn4iCmW6/y7xfD79
VJcXNrpoGjUxVwZd6K5xPpIvsi4rOmc5nnXdZxEyrotG8+OyuhcDXRADEk2jHKw6FwRppsHU065Y
dRfrE5tJfKWVmN/EeTpE73Ao7ZPUDm2HBxkp2yqnsMZ6FIn6Y2+2n60fOismMt1ZlmRRZuzN2QlH
o9RmQBq/YruBtoh7/Mpyno7rzqV730N0SH6v9Fcr28qhpfV4ZTNVmrqB8BxGsI/GFMPDrMfzw0lp
YWUQf6V2acxKSbSCtEwGDRlHLym8M+oWKYAzCSXUMF4G9UsAUypgcmpsM3THdpi8KOkPw5kD7+vN
mgPWnME6NR6hqnpWuKmNUGR8v4cTCRl+GQE051SBdQj5ho4gHeHvDhm/gS4/reNEAfpZPPZUMKbn
iIgOrL++rntZgIpu6KK1SHgCaaxy9rDUV/jriyPwpfDsyMTcgm3EKQJ/Gwd+QnUtoOaFM7gAW+L5
Q9sQAFgNAsR/gf1mxhrHa8MS23gRKlW2KkAdLjv0ygzheln45mPoePnzqIhhT+isMjSLAbyB9gT+
bl5RJ4oaV9GO4Z0kBa/n1Qj9P+tW5Nml0OCgXbcikhdvItRI6J2cKpbu/jdu4tXbSIpRkhsbW3n8
0TrmL6NDSTwFsnhzHj8HLtUVARqTAChVWW6/WqoZf/UKFiiPAbL1gSmG/bA9aymzWVUrkVjxBOxZ
dQDJBnItTXzOCv/UJd2Yzjih5xBykF5WmSfXQ+rimzZQ3dZ6tf04wP5+StLLLJWKUEppCSiIGVD9
p/RqepnK74xTjha3XPb2mk1ul7848KifjSjwg0p2DUU/6X0gFUn6FPw+TkEjSx9K2XxkR5I1tVuV
2dCK5jLoYNMrg6fDWjjMubPohSSN0YkOnsZL8Ogx6KyFsGhaGTDTbFjqGAdHhPBYlQiUTJip8b3m
uHFBxwou8YOpxbR0Mp9MgtDHReugY+3eEv7ibelDyL5D4E4TBHKu0OpUsqso1sxWyFmBptCQOKPg
ZUXmbKci2BG3YqUjZa2hNS7ghMfDOzxt6PG7YBp+vWYUZezlikLdw5RWkH2jAqszJvSdK/hevSid
FHJAMGkA1aVLJEmcow58uuGPxL5F1tWgnACggAMitVaG45whf4nEGIKuioJ5FB7yeBxbWxDXgjxj
bZNlEh/TwsfRag4KU0ufeLqMRSPoG5OdVOjmkoP2WUotKsNotN/CFD2Exm7B1qHoGm0Ptv0i6lkn
7c6j05NtfH/nmj3LlWzlOppXW3IUSaYcwohDCwF+03GlOqFB6NBm6PWjy4WL188UFO7tXkBa7+17
C84Dpde6WAJOc2E/gzErxI1Q5bTZQkiSAsDPimQSBldrIqMIzhkPWK39FPQMvvfSDc2LHEPkBwH3
8Ti/pC/9JfIaavn4zyRVqaeu+rshFmpv62fBQlkV0LToA0mnmwMWu8FXrPlDy3qyYArEfTYCZ6z+
yyFkVJb2cZ9vlJE/4PbrQ/RTOCzg9Q63T8JD6GDMBYUb1lI2PoKssdxpYq/0/4YuQgIAhOx+Woyt
qLs8TIg/8DUD8vhf/V+IL4lXSUDH21ukM7W1Cnqecp4vJiAXC4CbWuPqCEX5hTZwj2KaLmQ5QsMf
cjRsPn47kPwrfKUiRzCCtI9uAyzIzlECddnYQJah1ucHJFM+f72ksrGM3keqz8+jnYMuLR4H+8Xo
tlCskRssevcR761IMfajgIvl+F6R8+mxHtxDFJJ5XAlJW2YaBqrC0/rXRLNaojFmYuqy00AgQZnb
+lZoQfQV69m/KL9fr3AdpuYObu9m1AZDb4npUNvyi54rDFHmY1vLiKxQ2X9daYwc1rCcBweE4iQQ
co3pEBNx81UBLr4cNLQdAXd+8xRfxHqviVRa4sGBYKEpK7mnpYBy1TtgGbw8dI/2hVwz0wh06sA2
lo+qndjvc3byvHZ3olOyh4lz8KUu+vAiAtrX4tUMGOR6BNSW9MlqeO6ccRx3Ke48uEnUGDDERdYl
Scw2ghL8YOUWoN0gNPmfZh8k10GUK0cilr9PgDBTC5lIfi7gj9OWOhl0+MdN7zIr/AtZvPwVkPxX
o/1NfwcgL76zCSg0kcYGv1v2WFzXaWZxIJgihFF/lfvJZN2N/2ByNgrj74AGzqhSfUQUOZFO/ty8
YhZfelSgW8tIoLDp1pFM1SE1/lm6tGc5h25nSwUJwNTDDXqvvEusC1lnfiF+DmVwV2TOg02WyfP1
MDo4vRkgRjiSM3/SH92eoCTijH/DxuKM3X9s0lEY+Oe6Q/ia9dZSTLpkG2hhJ86NeSS9L+jjGwBg
2AKbyFAG+jxPBKTsr3C0jnPyVdVUQLTP6yXDq3ELO+Xuk+BSPAmiYyJe9sql7EDTFLdHav/M680U
mCOewIkBMOMfe1KeGxt8bALxRBJfoh9bkMlcd9fx3Yhil4c80/lvHSbsT1yab89H+TjG6VDQkrN5
9sMLisOmWD+b5mI4qZU77ITgVgCoadpah4Vw5kUjmd9MGtwfDMyAVsPghCJpWak5fun473DPeRBk
xy5gSSgNkIJKYcXDKz8JAd80izajf7/v6Q2UNkzNmKlOeUhiwpz1qOWX8WIy5nhLJ1SpLIEnziFw
I1pKlRyFzme0fOzO2MQuDckix4eJOpXQnvKvLutNkevcEJ3K9Rdzz3J6sAdWlrF0euhiHHcNVn+0
Hg/LvupMYhjYAvwCg9PAdt3qkB0+x8KL6lB+hloeLulKysFBGeXEjGpfL/u3f6+FnHvhKQfUqOyn
r0CQDakkW7CNBitjZRq6wh4B0OjZvZ3CHEQXeSjqAzCuoUSpZ6TMejxILe7VCNmUlkxjxAYSHfSt
cleyiT2ts52gJa5KwBmuMHNi/GAVt6LGyHpIWMu70BirTX6rz7CAsRmkU6DjYitvH/cJxLlojFCC
udDz8Ku+4e+gRTv416pREBB6GsnRtpcEcE5BEQ3KkTgN80V13JRiSx67uwRY8/76ND3UdinmLhI3
OFulwXq0J/BHN2vs/+K4lsxbOULD91A0Ip/xpLstQB4ohHGuvYIkgRaEpfq30xuBDqUHVkGnMzvd
1Nmr4AL28VvN4ngyYfATpr8ni511pBxwdcEbSEyolLmNKcsPhTkMpZndiQKcPlsbdHX0gqNv8QLz
c2F6D8n+5EGtGcpmWhj5iZdsOyLw7fzRZSgX9yvOKtJCDUWYr346jdwU6KuJ9qf1dgqWZoPO2/MF
Pk9qXMU/R+nGOXtGGaOBXfqKBT/D+EmLTNTenJIu6r1HUMjJaga8o0ZkdyZpEa/6KN+Nu0lcM44f
mrbM05tlFt4l08slW2u69nLBaWEHq12YlxwJLcOwtrD6qzO1Y10/xS3JN/3aWoX8muRwZfcF0dr+
YW1Xl8TFXQmeJFaIxqPvb7A5F0svKQbe3y2XWuPtT7IxItXOqGWHe+qd8PQ2IQGBaKPkKNfMDV0/
OirthTbAvkUmaKyKeDNjgjW1H722uA+hlwnebCwlXUyx6/6DTzJuOfVRf5KO82sQxC5+iMsaPwaB
1hAoc8hXtmMxeMmizlrnj1h1Q+Cu2V1gpDu6r0T+X/LRGx/ZzLkcsDy42SDUgYHLOCFDJ/5IK1hG
8nNuGepDnqvvCUa0yckVD5sgc+Fw0DnlUkKOBRQKiCwJtZhdIiIjiFsBW13KhPzZs8uS/usHuQ5i
7+DsSHsZndL/HNuRMxmWtqhzyJ4ut9rbLsLpJf7dDOTI+78dqAyImvqUQTFumqz2hubm9OfAlip+
BNtaalXPfq08O3w7wnUshbarCWUQvqP/wVyj54K/TaUuAUGSeDfaoLI8SSjdYAY2WIQAI3xDBqdB
ex2wp9roBz+hDeB0ikz/MBhSsA0/on8+zzd7U7DdED7UpODc2AfddP47nfryJvO9j0PQebcgKRAI
DNAhlSHx1jfrtjHBrKOfVDb7Ke87w+lgGn4R/c6iUV+JEqdDh+mGYtn9VxLxG8y/FX1AyRndvkyQ
APpEwq4Qe/AIjbmvB2oYyV6xEdfrSUquIFzWJJnl6XL7WVMy+b0qci1JAX/G7EWNH4fHeALyITnn
GsYWrW6OVqXsMuA3J6++mRmOPa/BRI0TviaK2QwERGkxI1tdUp/zoP431wP/XdFA52Se6d39Y05s
xhkZsHCXldrtUqm5zDtp9JGzJQn9a06CeGYzla4RMuVdIslTdSDf7PT3NDzWa/ZAdMz/urGwGFZp
KOv2o/xxUEOw64uZXPYsF/mdW7afDSl2Zy3HjaDEKuEtjxnGwIubR5oxgSDMUzZ0P5iaDHSIKIQ7
XTM8yMMA7jNMhTRPFBiqL23eQqnRyK6kezekRQAxIGeM8Ipyp8tDvxeYHtu/4ZsBYYd2kB+lqFtS
LnNW2kNzUd+3E7UX2xpPkvSx72R2djz8XJzAu6/9i8FR5kBBHr5le4UgLXNU1VEgXwZWQW/swdt5
uxGWjALWh7Ex+mAxqUtC+niui/cmEdGgN+8gQDj4o2RqgpU5kw+9wKl9InFxsuAUvZFO/qgIAVvN
BA1fuDf19zd1JdUdlk5rKFvsn3Kiyva1TG8+ODH8T9xQm/sUUSbFP8b2YNSY8MqwwDRB96gaQLOG
0waTNgeG7MHM6Nl8/i+jszVcq6pGgWwYg//R1yY71nUqQixWBupbyQ1OPrU0pk56FcDEMczLNocU
Nry90HatmFsWjoWN+iU8S5j7p9EcsZSmvPitcx5Kpn4TEiLSbQEuTbmCx8n2/vhrDLuqKuqQlQ06
gxYYL25d2ecl33rOsODPBojQKxpGvMe1JINabteMS1qUEmIQgI6k+7dqNFBBCMPRdyFF1CRuiIND
oNYkSBuzlEQWvfoCge/M8sM9+NjhSO5m5EJIwMizJFwo8aXnT6d2/9tRVIi+ayWESQ0vUBIA5XWj
KHZfvX8ezWdg67vZG2dRTGXWYEeoexnS7SFJDDpmiNXZo5KwYw7KkmBlHWQhJ/KRNiobpx4KMTP6
mU9EQnbhVVotc6273U/IjBUsP1srjoi7VAqxwDtp/zvQF7oD+rr3YptcPXA+z2K8mxwnW4ykJGSq
tauGcuqekfpCVgXxd29qV+P8pbXXhLsYp1nhvV94rACRA6XyQ1E6LhVBrWf8zT6KL5+S40g8ldcP
4KU14BygIFeGZIH3C9u1Dfd36BN03mN2SQsMc+0LncIq0eWe5JE9aqdFHuUkfTz8HhwvYgtSIgv9
aB2Evdf1SOZQe/Qso+fcB3/PH4LuoBgYe+iX8EbpRVmR6KK6Sw/LfLlGlcifYwJP8WhHEtr8toFv
LodolC8whtpUs90jc/ui4DsIRS2oyebp0tFDqgPCe8u4dD3ytLI5KrRTB+3AgoiAgjRhXc3XaHpI
qmeozUoJpoXPHFYvUOJMrmS/7rX2lMa63o51AYVrvLV0v8/93uTv8KukMkDwtPonszJIpzQMarQM
I6JPrKAjP1leN5QwMw/8YhpUTyD0tyLhh9eI+L+e6JAYbgV/pD1ky7VHGnPf5kiXc9HK0Q36xZfp
PUQWAApHVVCRJil26knBl4Bx/D3f8Cqc3BVIx9OLZgfZY5OqX2HC1I3whF0BXCO7zhW/g99ygriz
GzXVJ5fnoEN7s4LWSeLf21rNGmwdGUnvRSxdzTMJ6kbf2sbKtDwnFKlyIou/hTrkSRkxP9plkQY2
0HMvE36gb/owZkx0ZhVtjJlD+9qTaPN9ow8B5dCCkfszdnc5aglIBEbjVBQual6PRz57G/XEkv/W
XEfd7oVUtAOkJFid6ibFtCASiP9EUZczFlIr02j9O6jFtWp41/EN+o/EG6k+KaOKGHp4Az73VTaJ
9ur06WnGDW1/fo2XGUQDHrLGBA4kC8I8PWwQkdHUEPZq7yA5zxL7p3gC60IqspqtZnS/zuEcT+41
rzWXimwTu0gnBQE1R4L6dcpRqG/jArqzVfUKVCK5CnbsGRHcmsze8+ojrNTLg77R/woJVJjdoKYo
QvB4xAmyGLqbmz1QS80U5Baca9fw6HgTA+w3Ahsv46BPGrDthFyYTkDYty+bU6XAaRXV9G8LzAKG
9H4eYinscR9pikb7CLkm0RIeKy/x4ZgY3SrK30DjbRrk1kLYfP4vh0zdAGwkRblO43gXeU9n3cOp
Wl34ZEQXLhiIl/zntYL2aayVgLUouIB4zzTjSf0Rm0V7Ui4Pk/TGr2N4Pzux8JRAnLBPOKxtsUO5
8MNkul0N5f3syCFOG7eVRPRpVtvRnCqMCS3ohF0bbqqkbN2BFJ4D+7Mp06hFUM/mDOp0/a/VEkwR
eLrN8+M9R3oJgxrO9/DJEWmYI1Ao1M4eRTOZg5ypsYtKJYhnucMGMl0xOc2R33ilut5hC3x0FkxG
ZHGctes4BLmlp54/nc8mVVIKCFMBhHbRzBSdmlaSzG3nLaxOIu2lOKJ0bRQvDe5xoReE69jHgoGU
9f4zSAbJtmmnPjRtj2Kq9wKnfAQPFliAg4nSxCe6tH7knMqkg9k5C790pZWJgYir6FWe/QyBsnrf
6U7GxS2EOR0jlyusKhJsF6DpRAKN9R20NoXocbnqO8OV9CgC2eJouxNkka+Lv/c0Mh/MyiZwfewc
HFtwpNoqUg/+9N/CZ6l2zwR6pO0xut35bp6yl6B4NKBwXeqR2KpsyXGhrovyc/aETa1eJO3yAa2H
6pJYRwY2ZAVE0fUtGpNvuQ0ArUN7YqMcW7HzK3fsqoBF/h4gf0ORfK860WqK0F4Za7zMljpM+bH7
Dv0wer1Ajw2yJMIj+8/5jZChAkGrZaC6krss52Jv/Z278Upt53dq4WlAoy/G+GDv04JObvBl5e2W
JqIGzoyPw72lXGXQQ/7FTu7Bc/5921nUXkyZ+QMD3rvugbNSxzrelREz3uJ4JVuW44ZQ0Qg41/3u
Va3NEx8yHeTzJHa1lVFU07a6hskJfXrI1B1QtmlTqyVCJl0Oc+iZyUol4c4e8ELDpdmK/QhA16Iv
4KXNOFUYOQTnu2Igl6VH1iYWb/9kvCQl+ZkIA1J4tgFUvf8KfcKCVY9cPXPFWFESxhYMioo6axt4
WKvZ3K+NqWKL8FNIPag44/3UBtLd0QPYvFbE3/kQ2s+s6r7Eo//hVadBOTy0j7MywLJBsa8YgnzB
GWLXYlbVi+MnJVRBhYeMRTqfsl520OkjJkqDHRAc+hry345yWL4Jeqa0DoUbnrzA3c/WZHuduCz4
B9MI6PQEGruINtnggNFoaCxT3/T9LbcWbxkJm35thdimVtYHrHxjR2DSlc0ZVKgTjPzn9WI67uh4
oeB0UR6oC+PRjcP0sTCkiVKnKzfvrgYoB9acaIc3RpgXRX5/427MUe3JXN/uFxJ3EsSXzHQfYLQ6
mvALwoUansmKOeUXO9WPnF0yTuTQfUPTMjhuaVr9c3/M7Ud1LiqYQFVKG+5HndbLCZIHrAS+g+5P
1W5w2YCDLnoA73rEz4C3xQExJ1bLIBybo2m+R+BGRmiPRmvrjEekwcsF0zFoW6Y7KNhRefHzs+jM
8A2k6f/vLx5rR1sNhTSm6kzWuYafx36fcrjclFFYd2O2WGSOlSQ43qCJYNnyqkS8gbqHSxSI3zpA
xRs/Q+7g1uiRtQN1kDvTeakF9BsGTNveRDOcvY9WW0jT9pKBIEy4B7zPL5BnwYCIpWBVK/Nh17BH
u6I7ChCoW7R6dDUml5PvsUtxA4kmfCsJJx/w9rvQAzj9Io2+oPgeioIYRBbnsSZWdfnWuLrUFZAT
OKTTiH+jQz0DNQ/B1PeGHATvNElt235TIy8IkGjkjoJsRvQrR3hg3/5p6u+M2ycJ359LfvY1RsR+
nzDiuR5deX4UbVoOUATS0Th8tTRquxu2iZB4DQgV0PP3FWOsv7izZzfgPKHw4I1SkbUmYmKwTywF
jECko0UWuLv/DkVz+zt+2h16bGjOyLiqQYHAmsGXPjMEmlRq/2oDUGSvGw+smPnTMug5WpjPDZy+
4iQxOhWJ3xpsdO35ZncMVZz/hJsASRHW6Di9vJ3l5v2dCeSydobiBOcYwK+1xfVyPJW9laqWzehz
cP8WQzE5Crd1hPPDVv3ElHxbYyj2r5iMioDQbZ6ZrQimVAfhVL314FLFifyt62vLcCl429Al5NK6
Bj+/OUwgMVYHJUbfQbAwP3vtbfiVkz4EpR+8lcpZjP7xW/ODvIzEw9jpjBhg/yj0wM+hq6yyaDZn
hA34Q0wKExA9giDNFw6jsPHbkLh/d0HFwGD3YdGRhkx9nlTDtiOQ6CXyezog2/TWC0495+FZ6bLj
0KV2QGvYkK3BtLS43zeWhFacpBGrnSVtlCboV7DZK+awqARQeKEP4FZ3vMwxsoas1YzYhMQh0d2d
JtO3wIAuHkJrjuBjd1HmgW75VlSgR6Y13xzgIzHNA3ou1XZ5MbDdgXbe1eoiq0BU4x2PDuqeW/v1
h3dc5h+3FUL2IBGC5xxo1elGLvF3+jOcfr8SZazr+6UdCt/78+YiqGhox7Ndd8b3qkSv5zZj5/+r
uTlHMOy5Utu8mG3pECW3zBrFn4J8MJmqZ0qXOHhRSI/0MfhRc034VZx3f8/89EZyQJ0GHDTmatcp
u8RLugaov/G+e82EZXKyeM9DH+7qmqL7hq1pAwBHN7J6z/hhdNpV4IRm2Yczoqi4/4JaZOoXltgk
gS6T9YYAI+a8ZaJt9RGOJVsSnLxMkUnYIGLswQV8p5FkFNMOjzJ2erxgV04AEK5vimHbBws07bj0
UvHWEGW2ujYqPRWEO3RzKTnVokrryhHQ+6Jt/NVXBG9Lv6EsBqXotuFhuNSX2KoWuMwnuoVLbIUq
59bu3vlWLzS+YHgj0eW9A1KHQ8n557HR5WrLQAuazRj/osSOjt8QtpYEr6Uvl5j45MdG7gbInXUI
V6gG1GVTqNWoysU+FxH+GuaKnKUqhVdT1WtmBloUdAP1JzmWgZsKia+2K0PpvCDzGxWjXdR4E52a
mgLK6WCBvEQfCc21Tj4nLIwtA2zbgqLOjPVK4usj/MIKjcDk34pVDDWUvNmBxMMjBdpij9g16PVq
gz9UYPEARXm/SnknFZkvBnaEOg6umbVJSwOJPc8tUhqP8+eRkQS7ITVTufkUt0SnpK7FzkE6ELQp
Z/CsIXzwLGlLgQv6K6dgLs3ahbXBg3PyiWXtuM7i1jFcAYRV6iE+N6X2MQMn8oClD2cbWpwbUU8r
n3an9AcB433k2jYL9ODJeoxmmSa2KAB3JLmQxtbw0ISli9C6h9SR38WRtTgqWDvtnToNtInHSzh7
fnRNsFO4anmcUDqEMopGS0352t43lKv2XOC9EzBu7H7h5iiRcolRiAdxUiUndacEXALY3IEwplRs
lYbcHliDXj/AOT4Kc+C9aOyxhHbIEr8dOVkndpuMpzHv9EykTH49F+eo/RqKLLVMZ6oCtI6TOVf/
NkBf5ODOOyqDOnq/+rbKFTJfXsUqZyQTxw/ZRPHk5gBmTsRAsNY6DhYTLsGVB0usGmAo3v0yGi6/
K2xTaXhRscFObZdVI364/bggR5dVJK3bsaYIGBpjs6/llY+WKa5Pv1v/YwIONETd/8E8x1y3yI+P
wFjdYev2z7hObpSYEZdfEDP407JxgRDvlTx/kLP8T1GUdMa4xcuZ6r3l3EKsgdaz6DFrW7dRqUq2
SSskDWwC5EFzxWDz1cJ9I85MzWHT8bvNLTvWnti//rkKGV4yUV16YOj6La8qnBv6J3yLCJrZ7a71
yQEKu/Y8tYbX13/ujgQDObOsF+detAoPVwp208RaI7d0kozt6JmfHAw7UkcGRc2u2ikoyx3eg+xH
0c4itswsCc8ondv1z4HGiTvbpeOQHqQGdIDxn3dkIpdOYW0mb48oWBPNzfj3LOYmYjfiWP8W1bsJ
68C6avGaqnhPnsC5DSrnxjwpWmnswCD/BhZViZhsHjP185lHveDiaCgLGHZaO9FMkhR0PZQY49QX
jQYmuik8Wvc0FcznzMPQZKiCiBEGdCshBiSEerKrJLeRaggoZCeQz2vGR2+sexvcrRV/XAKy9SJK
l7aGGBnEiei3buP/L2oho6tI2UKIqMv0mdEum5bIxbCmsfy7Unjlw5IbLadRRiJaB02uu1RpNb8t
z8yDIj2elpGz8cJ5GSeEwtQeYz7y30GLlriurmPgEd+ezDXPJPq20PV3B/n6ninTHgTIVPoPVFSc
vGTpbpAy7cHYvohQjwvAip6dxMfRnDaA42v2SSJ9OREQhZpJRJNH8yNUajpT1Wr6ywdaViXGeBfY
71kOvHm3BxY1HDPqcRa5+EGni7GtsYNdDL9eGSJ9m46fHjEqMx8WNkvt9/Vo6q8RlFknS+rWt9Hx
Kl413SrqFfNJZ+xy6u3cHQzSuTnjngYwRjglrgF5tLc/f6Uz3WWqWOgIdxbnX6vAu3nVhp8SYf4C
HHbWxf0BmNap8XeOoo3fPneu5hPKKa+dY3UuTwhgejF9uMi7zk6FiVWba1jqtIGvnXr/Qu6HBQ3K
mCvJW0QduLrpwn2lif2zF/aKtlDF+laLTV7v7wAO9d9pf+/roYZ9C5QlohG3A4isULW9X4sfk6Fw
37grWsYCcKkmRxpB3eA9vWXABUkp3Q3g65hCLTaZQN5smNTiZN+/T5kknA3iYWsckvaT9Kr0a58B
kpX6+P30Nov5DALdYTc45fPxPtfHECFpWvPIAMIWvvqQPHns4DtIcQkJPdG9Slf5CaM+kZEBcX0e
/MWSio79MSGbsbQWPa2LsqLdMwM+8Jp3HgKsbDI7VtsCf4JWZNAcesw4dxlnXMa0S9aoJdSbywpY
2x86+svkuC0s75LWalvLLCZdDnLK/1TYM5SqoxJKdK5OJhYQqddbBRRUfjfdwGa4ivHVi0/2nsQ/
KOf7WCfRq2djI4FmwUEHrrBETpWLhZZzZS9nJGO51BaP7YTgT4dTre6LlQQ2vYXGCkFzrIvZHqp/
NxXhn/DGcOmOf0mEa30dLMJBPDFp1TLakSpvSae/z2sG9mZ3unI0oG/i/RE+SHzq6HJoszqre41Y
/3x7NdJOANCGpDCOKBJsjyBhsofPGF9sySmCw5ET7FCA6btU+i6h//7FHQuYYyvgUtbryIeuMtYT
27q419KT4eRVNley7oIEkS2Fs4rztJW5enGwi3sO0H9yKfNiScbEib4cT7/q6AizqpOnaGRgH0SD
Tk1JWB2YlIz055reiUIIqYWaH6xp7C7XZNpMqqOrr7Socw0WpqjKg+q/OKDyPaeh9Y/4JICuYT6O
vpv8xJtwvGgeddMDTgrBl9msi4Gp3P4ECL3K0XX15pAK7jIY8Mqmnc+EXXke5DRszJQ2MUXwg1wQ
A9KnxrU4mfQN5VB6UDcY+TSCE7rKmk0PqTa6g2nbYX/x9pvbpnbW3GLhV1mpTBj1cE0cF+KZdEWy
BMu21UGo8eASzRvItJVCBzRrWBdKlDKG3QeYB3hg4ZwJSgDp7vHe+X4h3d8Ml9D4B0jsYjdjb76r
QwPsUGVds458sr3z7/mrpEGoSxccRyfuKLPZfRhIRG0t177MVKVDV0YKQ0HwqP5AJZJ6J/dJkIIt
WfCUFdUltUFUXruZYIhOxbsxDp/Bn4P+I6vLJP5SJlexxRIbaSpiR7qPjuC72YDs7G5FRvTqS69U
ezs+QbFp4kYovGNT8Bj+7Ub2A3jAWjWH12uK5STp+OWOYzzvbW6tV3lNg+vRB+E+tj/CNgwMcOvI
zyEkDRfiIuzruO56h2TEkglyXW5SEb2J1YdLLjD0JjvObeRGRipTDlvM1YABeH8H6bsZKmwNV3aU
oR9AGMtrGF9QaJ6uP/GoBVjv6WvxjGjDbbo6c2QtjMPhaL89etCd9+iHPN255gmfKcAIX8Z0VRiH
PKgE0MCcdrqRMt0RW7zpZCG/PI6Sk7aQ0Ybm4DrU9NTcxWIolTL2Cqf7yEcRz6uik3HXqM9//SU4
FMRE3Xpga1rp3Ndqa4lMz7LPhBpv68LYGhhVW978i2cLB6bofBo1me+lWhV6ENphnSlf4JayMId9
34mRjetpFVmxqLVy5Zqrj/1Uprdc/uhQ/WWpwQbXUodTpz5E/tDqBwqxZsqyUdYCe5V7NXFJlWMO
vIDgkvalPS0SxKpAfXegaFqpdrQASDNKUknkRR8noklQLXxniMtwVv73D2/Ew1KYULu/IGzlgYwF
Dz012jNRZwyc+u0ShRqumlQmI6ng9cc3P8N8iUPCjC5yXTwiAYSRzn66ZV2oxuYzfRJDzsfgK+VM
WpclJfSMx/eGKzkenvLJkg+XWNW6P0AI1/m4YW98FNteJrWKg2lyT+UTKl9eSVcx6GPrxkQQgS/C
2pknsak/v2BI7ag0lmipRi4fBxoacVhPeu+4c7t15yefpfqKqkmJCjpDSpburIMNm1yUvX95QSqr
QN9fTwp/SznJ0oYSW2LFLiz5n2nBZkYumr3qhiBOnEbErxkDCJQ+xHNhIw/819CNL7IPoPmdO10E
zHDb7BmI+dOMom4ZRlxTD9rYl+qgILRleDJta1H+KFRPNPU7rR9jnKx1mz4fNFh5Gyj8QgDEJGF/
1bd+x9ZgR7V1i69c6sAEp6OrIobJ282LDw0pwFjQ35dIamusffs05hbqyg2QLPEJ0s2i1CWP/F6S
pmr5Rn63LmtpAgl0e69Aue8Cs8ja6m4VRm1GodU20fHdUGVIWrfaVwH5jHEbaFy2vuumAaQEY6Da
fszvMdMa3P+YMtIV8RCw1KPTWL4J19Q7BspgkiN4rsVSEf5C5pO8lcS3wtGFpgUmK40YU/dyzkUc
Qx/CgGVNu9eieiuEFdX95/C5xapnTJqXOM8HRD7bBmkmoYq3BQk3T/vmTDMPc56H6sEasA3/fxQU
eWvpTW0IHcMT1DqKTYpN382CTmStu7RbKc8Ka9rMUJ9p+FnpomYN2L3/9T331PVV7htnSivuFZe8
zFVy1RGiUXswvqyx9VBIVM3+F9NQE/gdvAV4BWaKzhQeWF6Xh2dj4a5jvPli4Tq8lSicpv/9/Ig/
pS59Ki9lfgp2/oamVgi/ffAvxgDoylUlufqxr/sZsiCb8ryrSYVYIwOxVjR9r5fqJ3EM3p5dIVVL
R04fh48DBweI6yWJPZmxVea2mOYTb6mI5P1sjwjooaYQKTlHq1QHxxBNQB/3fynQcoCUEIQsFMOL
cE14k3u7zjpETVMKxzB38NGbAS2g4glQo64ETA9DtfSwzCn1TR+Np4q3VpNk29Rh2MVuIvI4k8pw
/WkuhOEjQ0Dlfji+FDflEm5bGhBMB9HGA+w/1l8tU0GAcwojjuFdLHgWLYLogAQT1+u2u+DVmmTX
D0ZEIBZhuB2bP4T256RswDeE4nHKMkCwLgpT6C+JOIrW6ddFMeabiOnxW3h3MCRa/CmpmYu/zLCD
+QDVD6MQmvkEWMhtK2L4mBF47Dznqog3f+Z0N9WQPcMtuCTuZsviMIWqBFuplmzD11RiruUtBeWV
26tWAXIye9wJv2Die0XibzeE3ZyXjMNgGYBQdDeL3KVx6TrrjXONSDithv8vwZ9Aa+hON5HIgQl4
siu+f4y+WI3GdiR3otaZRt3QTleGWp9fHAFpqGvVfKU2qegdNVInlH35zjVmhp5hdh3OHK5gAJaW
biI15kZt7t+95DiSoCf3udpJ3eSSp3DdxAOrp1krQyDh37dT9OEvGtU/wl5wONsbS7cLM/pnK/4q
u0lrbbpoub1nY8u+Rh4bXR6VWWkdYcEiU7eR2rPUKaPQQzW8w63kJaEHRmv9c1JEPmzHxpszV/pC
j311BwWP0ChP9lWVUPEL6UqYWRlprG8l0p4nOBi/rTi2nQ4gZuQm+nRjZHgDG+tuzSVNy1w6c/d/
plOwGLoa/YIpg3q7dIVmB9WXyfzUAJfZXwGvnKfq5ec30OquQ6a1B5YK7fh/DY+eLG45+8xIndC+
/67jbDXai2fe0pGMPNU8L7ffN4nP136UIsIXA8Qqn2xiWlYc3JxyWI+OTTZyQoGzqb7zsF+Y9mDX
aoXCgBXueApx5651o9VUTyUzbQacyonOuMdDZ6qOhsUJFHb3oB6tnIMt4+pcYyzLTBrDS7bXIKFh
7Fp7HJapuEr1NSF5RfQysKpJ6wL5WESvo0VsQyZD4YNUCBx8JffNQb8pRhnmemuBz1eKdz3Pc9sr
m74cWGS+LjYtVIhOWogq6sDx87K8FTjOP+zrtPxCkfQQrhfSqxF2G1lv5BP6umvBQAY+eiwlS0+Y
Hwm/w/wEk+pbQax4X1CHpr25zqHwj25OIcQLeSLSzF2uUHbcJho8ksMqNuw9DgooE4tZoYKMZ5Xz
FlWmNXGl1n7hTO57o6hGuzQIxpiPhrWwSAKm/xgBwtZXB6DN2MGoLEvhCWW0D/AfVwJFat8vcvqd
k31ANr5//DyZHn8fJIXiFPIbYQ95iSr0UxIb5jXAGD/Ao2D+jgpt8RmfxR2hkNblqPC2BOkZGv4T
Gyl7nImrUSI5DCqYlx4Me7eiV87KxhVJLGAh52w3oxvhvrMAuZRuirJn8kbzs50efa7x4IPYqm/W
Em0DDypiiKpBmFSXKYa1BvVlnM6zQJQduS3nX7ivZf2c366PFikB2pLG5PRgkrhVIEi0BWOisqDL
AX7rS9SUnU5hFDyTS36LOa7ZlGHmrJDJ0eH3m0SHV2gcELUs+5I8NBkUMCBfpUC/FwX849EL26nG
4cagRWwDWtZbr44Xbv0qVdTTxEwrbm8fXDFApZn8o2z1kTrLFtCWYiopAUbzzYRNooaim4hLeedS
YPaKiUYVoe74SZlmx92P/ZxLXQMGEVTiry9bMtBlMA0Sk/wCnTey1P8w/+OEjvz/tlaicGvmi3IL
Rg8cJroBadKjZzCSdvWJthA1fLKiiMRLCd5Edg22AiLAbkc9cL1dXVE9HgU06a548/UGvygl5u35
sFVVLxq7trOI7MUgbJ/2pkDFlxJerzVLV/MoRPEIyuhEWaYSM2Frnk/zH2uikCk0JdH6iPmWcsrR
tkj5yIyx52kztMVzccDdOMIFQ9bqaVg8Lnh5u6iUgdvJaw6A3nm8t1k3lNFeAspTaKJzV7EQv8Te
4aquoGsJxHuWnUdWn45Dh1QFQCf9/LWbmUmuYCpuo50Kq9R3UkJzR3+mEZys5povQdEn874g5Y6j
E4TkzjeC1UYbC8sDmdr2d2EBwV/QCA2hYF3ykiewjIenB16egecTUQ486Ap5jvGard1ST+cq02+/
fbcDyJDOL6YMjv2ZsoaZAiHPVmTcoMFmWJgTG3/sc095kuwIyXmdKn7NYTo+Z2Ly5pTa9X5C23u0
/TpTYj51HRsOs/OeOCrNMItl1Mvn0CYy9gHdgu2xykACCAjm9LFF9gNAH8ZCl3YRh7FGbTONm0Ut
NfuA88fB5Avs6jUlQfs3t4VzfBWVIQbjisJt1YQmQlBVMWE2tj1QkL9VtRVd5U3XWqgQwPTK/IUI
EmZ187u2ayr4TRSBOYSOLTczzjovh2wodxDNPoVApRehmRkQwZKTYAbztZQSS9kLJ6OJ8gNV+t8t
Zsd4H8B2TzUpbbjSoi4yKAdZiNduuxrlQ3EOg48E0wbZvneT31XuiZSK6FTksczoDFr5C0ZY27xy
YCB3eVSlgJj6NHyHfkjAKrzWgZYhV/uFS8Sh+MhbAv1pTRoY93o/BTFyWKsGbbGoGxjhR6LKChrC
GdiM6i2CH++wewSVrT3UZSogmtvAuhADF9beSIaNqHP9L8L8jmY8Tw56EJMg4IzMsYVNkMraTI+J
agDOgefacq5Yvx8ghgC7uRWIdhQfUNwKlJ0kE+HoK6okdYoWsyGjcgqkjq7FNJUx6uumQqms1gYC
wS8+rMHrnnYe1alxpSPd4A0ENyuUmVlhhrlrXgvh529nY8nfBu24RcoB+6Pu6naWWKuOgxRQDoR0
NoIEwv7NvqR9jgv/43JWosg4s52JnxTWq4WZewCqWuNzYMRP0AMuBpaySt8WYYSVVk0HntxE+h/p
Nee+I9wQWFkRuWVKx5+q+3ig+giHcOCWuQ9E6WrQEG4KtPt0vAherczmqxOA5GgyRtPUIspd6vwJ
Ms6Y9JjlQJ/GtPyHELWDR1OJ/L97kggA2lTmesH80OJN3W6IbbgH69dNFBBr4j6UFKNV6wl3shD4
SotMkIypvpp9s+F3LDi6eqRT//6akbLe8Abr613UK/yhDr+1gmtjdZwH4Ve0JcLS12GWhg4Gpe95
S7Hv4CuHzySffx8XZxAfOa3UxfsseNOOyBx7OtyXHXCZ0T7EsLK+WHTwlN2wppiA1GspkMh5Zok1
c/3sWFaPxZH+P/TuPsRfe2/+cihp9CIZzUwGZHRHSdMW8z21BBWTNNOI4wv1lM8kTsjYe1Wr5Qau
ZIqRba152gxT5Tk6bmF7CcVIJv2W5ywwKp/EhnMNy2tBTGnfor3IkML6TXIgzD+kddm8h7cw5Yp1
L/txD3mSPW2pC2Tqi1ufL1AYo5mByXBx6kkTmNCN3VxXTiDTMw0TLRoQZrffmwJ4rbcZ2IZedvoj
R1vn3sxFdQ0mkEbOsWxTQpgnGzTHJOzGx/P3cGYCDSHRNcNZRs1rZGG0KfeGlQi0N7VK78odCyPH
0JhubduzmmCuA3CiP/E3Szs6icqU0MDChXKp2/L3WsB1kKivq5sHAr439DtGJaTAu7wtn848DFLV
4AjRYABy3L+ZbmT2VOhV34DqSzlJoaXeysbTKksjwQLI+Indmrq34rBd5Me3e0MJK21nTRQiAM5u
e4sl1RUyEnPE+EjH6pvOD9kAPbQjmiZ3ZhG5IHIYEeYTjnoRO6d2t+ZqXvv1BSZhrKzIeSMzg/c7
W63/CHaY9t4lVXVdRePx4udvIja+sOAX7L0aSbgb3p2Y1ehcERv5TyG50FAq9zrUSrhJcOaaEpdQ
PiWEaduz1z4FzhpZuhymczWlt7AHKmhusgRtr2RpCiv7T6RiVmNjNPWRRemv6nP/dN+Twaxazucz
MSDaw1jzwNNrS22Lst+BaBeOVASbCM7S4uTsY7VnUkOKEh+Bi3d04A+PryELr0MfbM/2e/pz83s7
M6C/IGlrw1j8hbKY2uCCCq2noDTnGDGnKQDF80ZkegzEu2/1yV+c8xH1QzLtTlAIhYrYgqfiNztV
qc1AKw8smc7NQ2BZD/wo/d8boJKrDcEO24YJDDV8LeYev2Iscn3i+vWeztIH+R5qmcaLnrE+Reqk
/DiPLy+/6PlR9bE1jtFFyGYvt3pecyHTGnhIGnVGeph7hBaAFKnkPTYuOSKPmTNii+0dklG+XMCr
az9CgD8wgG2iPVwUWJ0E7lAIXrQ/YWpACcsdRD9G0sCKF6jB3qDP7nK9pgi0laRv1H9HT7k5bJUS
VqfVxwOpcLw/NXzPjlVgSdZ/9h8Nj5FEC/TyAUucxfZEeqk8M059keGZ4Pbzj1vTeh70iBdIlity
Ws0bxiFnqrfsrRtfFRoSxsQQ7CHS1nd7AZPXKpFewN4dp84PeIgwB9yMH4XIgV6q+aI1yYpjVKxf
F3J55cZb2/tFY7YFSSHy+BOwPQGSudg0s4naDmfK7jhIIewz79rriLU4m/KBScniURjj3G2A57Fr
NskQ0PrLA2cn8B58MbTB4VxkAe/4xj7HtmLBLzRiGZmcYCBTJ/B+izVh3FORCgB3UjyCqktPUbH1
QnOgx7Uj7/03/UzDVN1etjA/ObpVToRV1PBfM1i88F8u6rm+B9OLGpHK//hHO27HgNKlzilAieTt
RwBcyEPdjO7y27OIiUeGOKn3AL+OmTa1NB0V9EMkV/XB9rvT1VE8iYm1UThNxemWFtvbdfc/FVGP
TFz5LzHtbKWpI1xEgaXcJ+4ZCNON3dO6yOgkaFLJ89ZFBOUf/ONb5Yr/BO4AvPTOftFLf2wEo9aD
S1F4U8zIOIjSNkFVxMyYjXt+7LwJzqO2R4wYTVGSge2g/WfHqoptxwuXi0xJPSM0GLEqlLrPrj1v
XQlE7kdAxgRZZaT5U+SJVx7dfhfLCbY5Jhh0ernCGZ2/7UYAtSgmhIq8xOmX4MlGLS/+fSJkGSUx
uQgQckW0OXGUO76GUFdC2GfcLGsK59BN9Y4T4c25mncPbutFIYFb7hYtcmYzZIp6dMbkCpMVT5Nl
c7fDZUn7w0pDRygP5Oxfo7yLYm3hJS4w5aJBWszoLRsnylcb0d4mggfh8MjT8Q6O6EjIMOkIplLQ
OwHKmkfxCQSBqZ7PEGgDpZ6dilfDae+rcNXaufY3ca4Sk2cQwqf/fXQ7HujGZMzV6GbIsdlTSrqE
VrTdm4sOh3015NRX96KUwe1ZG6rSAiMEzDEIdqcq1tToxQlL9znWr0JlM+VDt72W0RSm0361MWWR
lE7kWYSdUEoZ4mEWU7y7EULWY/NYIcjKJsKSIgkBSHnX025S8okHCr5eMo8n3JVtMVkusl0t9urI
+6I3v5QYQ2lV6Cs9lDukd0gv+U1sfcHfanum4k7qwv50xRigJXAq23oKpFhcqpyrJUAXP3rE4EXI
+UXCI7dEXlhz4SmGZ5lr/pHiH71ll2FurcaI7SiGZCh4IsIe2VNIZElmeWAHZhLuT/ybv3lR5Qcu
WUNaXBoX3SxqfQdBz8UaKHa0PqPN3JiWCAcXiVhTBl3oLnQZKkKHTb/ACjGBEKL8cec2Gyd1VEAn
emYox0OPBfWgV04ZtWEq2hgTD5F+kcd4VbXySLQ3dbeZiSbdQyEvbbn/mQWaEGxJUkHt6p3R2Z/7
hku6mA8h4vc0lEe6eKhYhYoU4dVNZA8pMz0lvKj3s1dSqVb4alhXlAllq6JpTxvE+XwWIBqA4Iie
V5hfecL2kvEVtipBxGPdRkSFE+WSW24rjWuVsL8KPzezuq9slJ6/Bsq6qMDYvx7PZsyVd75IQFXN
0SSfb6ujjdpJudyBTKF4wc8PsjOTVOfkzNKuE6wM4rinUHnN0fib9CRAaabRSveLblq6Y6LjctlE
w3tvBPge8/v0nij+en7yVcoSQShN7Truz9k6CZ1CWljRDeTNdrfBdZqMf0LTcpFMzedcmfvrJ3Fs
fn2+XVq1aTQiIb1RBS87Hry2fzx+zeGBCmIfWifSyKLg4SOgct2uSni4PhKDQLOkCle1HUUtn3gw
PEhYONfIqkdLj8MTCF6QXItVZePUJm4AuwOd+I0Ku42/gjmo+aP6JF+B/tOWGSrSp8WdtrtkZy+X
eE022eSCY8FBGSOtkfomYz4BFwMo0TEi1GdNZxuCVdMFeUKtE44hhC9IEeowtjEejN2GLqVufTeL
2/nOibtuMhb7gA18IKaoEp15E39GiPTC318KAEPNVIltrZDD3ryl9Ju1yr/VvRNSR6uKzNjSDJIm
gXDC4RtVSf1SwiNS/Nkw+INLlP2JYy178Bcm9GfPECIv4RP5us1OMypQHJZ+hb6jdau32g+ecUZd
4ksws9S3dCU4y4LYpAIFHEkDug5UrL0mUsf6roQlw1Wb8UNMjtunR5Q/yr+5kLYgYx8H6Qo9z2WQ
SRr5vxx89cSWGzHCpnjyuJ6czVPt+V7jwNQeaJ+Jq9uPv6/uwHlvkOBq+vfZ1RirSD0QXyCRxOWq
5cP5YXpeEBlUhIk4K1w1N8Q9ZNQu+rU3HqZHKTBMd8GPKl2sqLDD2NYSA4GptWy6ygCm6Qj7eFpx
tPEWnB6Yi2rdO5qW9N0y13mMw9JCpIfQS5m4aR0SAVVBhL6VG+jaZWhAJy2RYGNatPK0WnbYBl2z
uEKDE0uGtQ+poRQkpz59fO/1Z1hr1BlaD9STeFA4pwTc/SYStQrcLetndUivLqPD04jXLbapkh1r
kYP4bKrUASm4uq7zr8t0cnEbBm/2Vz2rwhhCeOAQjANcLF7kPHXoN2c4/zsgs8HwXRMTdbeqfedC
jf/QXEM+Qc0w8K9V8cKAAw1CbxjfT7XRf9TCN04tA4wL/rmqPgWWLnw1dhaZnP0R5/OQLfKHJwdq
X4D8naEhSWCyqJcUfjJzCfQd//DPA+4rnckgZW8Vys9mPsYvWG6cmVpT1roJaEOKv3vCaUQlum75
MBV3MVPl4+9wbn6BxLfe5u0exYXZr0LAgHHPGxN+Z62v5jnEVlAuVbCVmgb+EN8cJef7fOwDtRav
ZDJS7DAbjMLON5je7oOiV4LCjI+5nuxBD0BajOj1j7cPITvX90MJSbsW4iFzubu/I83TBO0tRbLL
lSQnI2r2Q7b1cN4As3imXvPtC3e/VXK99dByXguX3MykUMAp2sLxgzpl5gQSf9rbhSqBolxfb5zd
nCmqoLNRiZIQc95SFrlzUsR3PDuepL9AcgPfVCl4iG8r9NbwMZmBCWJbzG8qZLltNCKBFF5Mikpd
79xPeSvoXRtNPM6bJQ5sRJf1j5Dni0oLZnAQ09T0SAHVXItT7ZHVKrZ/bRjnhQA9dybmHju2GNet
YNW4EliZOLa+HAsq0126fCzkZRK3YLoGmotdVxXgNi30UN7Cc0g9QsvAOWpSlkEkihqo2R1aYkrw
n/HPt3/FHQvzJg3IHagVYOrW2jSRVbg6Oua4FAk2zvm7mKJNRaR9157qZs/qWftG5IMK9Qy1SmzI
XcalPq72c7B+m5A7GJqqfEylOwTW3WhUUJVF3QUNAcP2OLMoTdhoOAilk+g6JJAAlfygMj/gcoBZ
nMMEyovd0qZd01Bn+rH8Lzk/WideQtV/8AoTvnZiQBo6cxISGsvyQr1sfyGzZk4jq/7YASITS9Pj
zt4M2vVojD5jT8y3thfMrPF2tQQBi3+QFkpDHXxbhxUiwSNp0U7nigICg054msbOYY2ZzzF6pqS8
kbeiSc2Jtbb+Hmkm5nXNRBqx7b5BL5U5ZN4GaWD7YX6s7xZpH7bWksO/wtMUxerW8G2+lrXjB6Om
X9gacqWYp+txV1KbbAZxwAxXd8jqxmRTCFnD48DiS+wsaM7hVOTR0zZqt4h21iRjtrIxQJb1viP2
+YWzDLZH4Gi0qL+Z4uibe6s6Y/3onRT78zvHfCwDamxd3OuBtrK98WSi1o1O3jEm28/MX8y4jsmt
670Fs96/aNTp0OB1bdUf8LaboxO9vupn6a/AWrEaAhMaAvrRbL2+93is/jnwLUPOEE/Wy953bUtk
ux4SwZCgvJ/Smogg9NYQjrwdwxEwW8L8inIJqFKhzW8yj+sd68g8cc4mAsTl3Yf4CRIgk2vu0S0z
zcqEAaetSIqyp4K7wiMdSeNeFga3/xC9d+iRqSt4F6U0MNy/2AuO5TYFALU7267jj6a4grQq/LSK
WksTMhFfhveqP/gA4wbm4hbwxhdNmaSfo6sO7IttBWur/TDzMB5s/F7mkIWUAKbNYBnkEs1angLJ
aSt1EfCr3Y9gZypL3hBZVsV+hvIEeiwvCJ6nEIqJO7lTlMGBnIlsMzqiOUL0a31LkHxaaiv1JYmq
lvmFTWIxNrN0I6xuV3Lnxq0h4pWRnZSkzUnJO+a/UyMn8FzwaCnrQbTO3tDTMX6PGf7jgOVKKzHu
beh81zSIFkms57pTRAP0rvi7e7kIrm0gEMwjX2TUK5EDb8NSt8Jgak8pzGiotXx8ZN/OCxNYxVjW
eHvIEnXbGPQI86HKawb0p1k/dAglRBt7AFYaTpMLer+BzGxundPcbke6FXr+JLfXMdYcwstwnpbB
yI3+nj5BfqhRPL3e7Kz/9hRJ48xQ0xob+zJo1+7xhy2/PQsxM/fma+3sxmlbsXGtbr84YcX/5SuG
mkb3WA/LPZHWG105c7JnaVxhZczIEzFo83Hf0UbNaA4zct9YZOVGb3RtVcUJkMA15QdfFRcOYIeA
CxlXGcWnoDQTw0stJ1i0l2M6kzQFOWQmzh1UN5JUBTYJDzSXnU6vHDXWSLhHGAC69sl7tX8z3X1k
niPOsB2tmNjvaUKuM28pF0bTdNWBPr08Pu6y36BTxoX8vFB+bzWZBFPWGa+jlSFRxYRg28gV5KCq
Krrsd+4dNM3TysdSqJIxj9MorroMLXmac/cNz1OIWv9rOFO39YAlbwrttsTbQQboOrSj/oSm3Xh+
gwPET5J8+TsqeKHEA2qvq+gLb/Wut+6M1vslj+A7Z/GzAa9nDxb9uklBXAgOj9dplwMfZBv1bx4W
Z9t+lR5QF4IyX1RZqpz2dyEfDePBs7uLV+HGdmM2/bCKs8qPHJrabHDMWsIuorSbKsFWmT1oZfSF
Zmlcr30WcFsEsX4QtNqcrw3dlR8XH78d193gnti5YQp8o4sg45JkiJwQpSEE5C/gqAZ8jYZYfoe2
ak9tCU9qN1IThOrDAADj/t20POQPrvN/Y6cYXr9+ujDrsHgZGS1cjzc+MeOl7Xp0BxC50B+IcIGD
XatPFZ8kvnr1nif7rmLk9BO4gfYj5HrR7lMe5aKDRUBLiuUjIcJapFvl12RWrLNcr3vDiixOBkzC
nt6Os1dPKXGIStN7Xe1Pj0RQjSc2Jn68t4PwovvFj7ZTcxIEmu9KcIj1jgrhNOKVpnJln5uipycm
2n4Kt/KMqDkfviR+8q4X1QY6FrFNAUmzKnNbp0f2Dirl7ebwK1/Uix99XGpDVDApOmJmYh/Iu23n
1E9zmmpHwaCNqisOjdSijhvJZfdMmlhlopCdir0z7mFMee9y5aY0HbeGqjvUg2/+IvHdV8bNNKZf
J8nmyvyS8xX4ybdAu/zJYIxSCUurhf98I/UohzcRpmxmTrAWHAfK/HThKvWRR40jhoT5FiyfCopb
aizD7SwB/Q2PlLINB0psTaTWi1pdTfKNyoSdkJ+eGUZ6O/kUvLT1leGCqwncQQl6A1dRuQ/9FHyo
aO6Urjqp2Mz4GqG98Wr+qBrqjj8A/8EOCdg7eSDYxOtRUmPZMcWKy81eGAz+8KuNCSVQDnshnl2t
R9Z/FGFL+Yh5UgjkF9IidnHy+Lwe0wxHxGG/0fwuBrFwcbU19WcMCfuSdpCdfPwYO8R6IYmzZK3K
sRpmRgU816S5DH1ft01jded+hT0CXpBpFHeppCc3DWDHB39Oy1tSgY4MDB0Q6fTOV5k13wZdd1QH
zdmCtz4zYDdNFW/teTpPCsPdZHLhhqgUtpuCNA5DjSQnJDtZTyuHZTTTdrIMxqdgKdGTb0L5bBoN
Q547T19fbyI93RBB+MpG9TxT8S5vXkK1Diov7bzGuSvcwXU3ZdL2nYwe5LtT4Woka9Z2OhJyLIje
0lOcF8NhR4bMxTqJFn8IdY8ohkS08AvacqD4rDzm80RaBJox7Z2yRr2chwJp1bAsXjRB1Tyis+af
lWBTGMiRdazyYmmx8FFS3aPl+naX9StZz6Yd00/ubDlNT/K2GCBCKFMTK/a/Bk9gPVUDLIOjNK0r
fXiFVMgKgcYTZVgRcPcx2W3qO+hT6E4S/M2Y9VgUrwXL/FmIRMBH/M+mlH6vF2V1CyxBKfKAY1wr
eqYmis85ugwD/SHo13oXGQ3SD8OUdilR79hzqPSw/fAgBsZaIB9W5T75KB8xMk8QX22Z0Fe3ngS2
Q8gz+Bn1OfCR7nW1nc7S0KJYgacnPPUwoJWn3T9IM1X92Hlo8CWrIZviF1AGitSZzxuf/pbLSHAf
6FHmQoavUThpRcqOHuBM1NZEkP4ysjFZh+Hq7ALIBUVpHi25IBpTZX4mEYljX0+cVIZ8bqveIRjH
tKkahADtaeIB/zFtdWUP+F1AwYU5Dw/WCCYguCZzGkQUtFCDX2o6Fw2ZDwCUhJ8z6LCvVJU6uDiI
oDLK0wVsT9ksLq7v3oeD1Tv6tiMAvaJwsH8/fsrj+1SMpkVROLaRWMC8bjiY5yGSMrk7qEHYzfbf
cxEdpD+6eB/Kyk3IqykjA9df1mT+WyBriTad0T1365jLpBzJA44WbPJJiL5jSFNBCuMHNdGX9phf
ejHoSnB3HpLvQAb9SOD19i9JPDD5OoMfB9icx3Fbt8MIxr5dvVnZ057GbPvGFxcR8a8Ff0V1oT6M
nmmD6jdtvKyhT9SbC81Cptva1vF1DO9N5A8Jl68cEcfiYdXSg6+NRWvurST0+Z5FZbzbUi+2axkd
MgMZTEH49ncWhfZ8tfM/gw8xGNIGjcjnBmebfYlErl0HbXoeTBLdXBbO/qvTX2Fz2YDmpLzXveTh
Y9F9R6krawj3tHh8WVymf1q0Ub48hFFh9JljdooMM4wYZRNlLi4WfAcuu8swaLx8mXJe9183nwqk
+NAfLTuKDTKBVPh/NPvfppFXDf2vHaC5/F0FKZohgzzgNxFYq7TzXktJPfbeFb6tKuwtkuAxMyML
XcDHT1okFRFBjNFc7ActymqAcxyapKafp/tHqX4apUUm39rfv3ohUYwN1ogg04GkCPslWDezc0o1
NKEDhcXpyaa8VF3j1GgS8LEemHTQtSTUL/3A+cJzb+cIFuvZyW+P6Xzg/J5s08exJmCVxh8CWANC
c1T+l+pu57i0O+r2cXfNrIFjI7l4yvYxaOcHxEK9HQrKQad0DHbfx6rXMppGDzYgXwsInxXZADZm
Q9iX5gFSXCWFgkkaRyUL8YpDdAqFYMTygF/nUHzQpcc9FBbuIfSjBQZA+Vn3FefD71OGCc1xg5Zz
wEGS79eHewHjKzY7rs6WDikht5e7xSDFX2FlAWfOF5oXtdpbO9oQcgZaxSOHU0sJkbHv1spd901v
ppSIcbnGtckcZAPcduA4AsKIJ9j+dqaj0wzsjRuzEn1ByHfkuvBZ8nh9ZGCG+sofv+9luSBS77Wv
RSd/m6mFB1ZUzeFfBQxIS8nfqEg79UYIe4bVLeM/MDH9M8hZGdxa0GfOoKGqpbzZ0YQThpUsFKoJ
JXr2ZqSzlDt2khYw0nQoqG4llKYf0XlD3wB0f0MVvhC8eBzz36BY/dURPdRQAa8eSQiPL9DNkBG2
u5FuUZwFgKg7ktx2qUuU6ljRwsEpr2SkYOSAqsRsym8mHLcqR56h16xCiGzUpRyrdlW8XnpgUbl5
bCoIlq49XKZ/qh/DlbtrQW4gdq8FHDb0yDzp5Rb496Dm+q7YP219UwsbJiBMJyOM2ikH9QmavswL
sUO/TosMEY++vSZpAVkvTXGRZzxdedO7ZFmnKv6DoIZNI3+1LIW4DMVDM6oizl0Qfsk6nD/LKSAf
fR+Uf3wJf2Sbu+02+DCMSLwy3natrYFFfzWspwV0UqIY5EwD7+QLfzJgtWNBGwedOYacvNlAv4mW
CWCNl8/c0Rz27l4JF7XkbG02c3PNtJQkGrnTiswI56sbK/Ac24bh4qaCmIISSRqD1eyx9no2YHDF
6t3OeL0mfowUfgeMhImyy83g/IfUiVZjN0yDiNYQTfRoFXKvusNfPBwpsZaLElLZpOcRXpxa5w1k
0eoFTzWyC7w4+wegozJxQ2wUgGV0O4VWoCQsKIsfDoT0W/FwRO8vbDdBcHIh/ORcTYx2kqX16ide
kBTV499IfOwolC2cFoJpUc1R8iYIVi+9nuNGyCSKJsnkMefwwr1J0EZIt9ZlIdV8ExHm5velbYEE
Yq+7Pc77YyFCgambCcCXyHukSy726WL6NUeh2KHoCH9N8VR9Ij7CHCswLMAdf5jlUcY+W1LUGODi
PV/2eRo20bf7QWLOkGFSLkv4Errr75kFA/PjCSK4yjYYZ33KMjbZn17tjyjkTvDjiGIK9Z9j8W6O
06cdHSkQ6o/D+v0RZQawzcN5aRDmL4gQAyfTQqjudqw14Eq9TkiOPHu3KDbBxACJM5j32WVEx+jB
TuVNl3GB/LxRX4OcgpJA5JUNTyM720DrfUGluOCEMFm6YNr7+fWZExG58kbCJNdtPqLLizeutbh6
XPanhEmajLbt0AimP7fKZYPM0lhOnoM1IHE+n7OE3cTxhKnFrYtnvaXs/O3D13w8LhbSn2W08Mdh
sXEMFslQdX7GGW3z7IpBvvIDp0YTWNBcRxp9swT+WiDG2jOQ2eA5GGe3g1SeXNHiD03aVQ5E0dSv
Z7F2YrQSqXE4lFpMv4Xy/oZ2qzEK3VQETgnVB1Tg38POBYP/2F3vGlw4YtYA/UnnLI/V6G26ifK1
4+VtJIN1b9/yVi3eRYS1kpUaXLZS9Z3+DxsWfcAlF4B9w65KB7Bgx/l+K8G6QkRzfGWlJUVdJOxW
u/l4WHjK3FybqIU3DH9NR9c+xWEaygxJLiujivpNyn2yu59SV4xlFCv0nkkoyn70Jcm7wX/N/BeS
hNAGaGG1Nn/T4rX6XJF2zE1WpkXgZg+rlahe/xpdOKbKds3Dnfs6l/9oJ5tAcDWdKKnQiPFXa09O
pvfR/Zhr9hQGarZg6b+snJsckR/dCuWtAEu4DIhrCzZYRNvfXDS7QQ+ajhK2JWIehwXsazsFEQdp
zNAS9wZT9cay46BVkEHaUjxyjd29gwT4HqRDWRexsUBO9DyXd5VyNmea9vaJbCRpsreoUNTwxguY
3Fd/qwK1gAez91fWPOWq+7/4Zw6/LwLgFJY1Yi1NwLb9pYe4LAgX7N0ezGLTEAVPBvB6xPyBO4D2
MwAnmnYAygF9gZos6gzsziMIRYvxVUYYzlS1xQCCa7NjuYO8qRVnSLqyi0l7tfQ3u91xJD7XOmdQ
X17c8y69rj8AczS/CQwddjQaS+sV1V0JPvgG+604Mw2DioFw4Sw1EwCgrf12bAjRjdMi6HO54tjs
YpHSQrTh+NCuPWfClxvDUYdvmbCojgoefKwcGOkc/buvd/4oEQ2yItoeDCNEdVq/tSCWpI75/Woj
Y/xU9BKfgGxjXMfuiEVGU7T2v5XzCamnpWgD82Y2npSSdGrg5cC2kc8uXdQqAS1m7Zf3mw8hlGsT
ZlhGVbgKCXXWM7q148uTpxAOa0OaC1naRFUKGrWWtWA8AVc9dagUHAKltoqGMAq/ZfMQS0YTbabD
sa7JH9nYqd5njlbpGaEIkBMw1H18IyaFNQgvNDpRLqv7duDqn5MeVtYLqPUP3qrPkUrCHZcLXg0Z
z1VIuxvK8mHCXH4KC3WYTqgUdwi5YkTy1H2bUAY6ikeJnnGpvaDwlAK/LRRj/fd6TR0I5yiTva6I
Y75NDy64nhG/z/I5lG5KymEsu1DBpn5MVQOkOxI/f+7pFOYoNtLlwcP1Bu/Z0vyy21291BRHEOBa
VKZZp29MQpsyhNV1ps5PEA8xgvlK2O4X7xQOXQKQtVxjXxJzHL3DTEqaR5aYW45Ik3pgKVW5W7S8
UqMjoxt96llHhXN6FFw1+O6m95sIe9QcA+aPcAqniYa/Ce+yWLLNUPVfZHCiE45RfGpbQHOByr+J
I8pk9bz660pc8WB3ksLcWIKPct79u75LiKwGxos+k0xZcd0pw3pzyuTfX8mpksW4gC+14/uKRQQY
YP1YvQPh221sJ1IsL4KxPfAJcpFLdzFIhwaRdyhUklErnEWSC7ssAz/WlbIXV5A8k6CdXpx2tOL4
t9PEOqmX3Zt0XZpzlHFj818XvAFB2PBGjR7StJqg7RED3aDR4qJPzx0Lly9JI+Ob8mUGGotk2P3O
fYPvuSnx/dqTZeeGPAOrkRhRTF4DbtRsNdC2pPP5XGxHqfopul5DR/CbugkVR+yF1ptHQGY6w+KY
KHCW8qF2ORBW9xpta+rSVIVV4EsKq5OjFZK7gK6/Id0oiW3Lbo/qGYP7GevBkE7BBVYeMZWYDZe2
KnTR5ja3tMUhHTfyg4tB2AhuYKiehE2eBBCHXgKKIBMeauSV/pdhC4LLJdkvaf+AC3vz7UFKCg1z
jCnB93P0VqawgMfLFQ858Ut4MEP8x3JDnxr/+SETYxyUFht+4HKlJpWQy3s1mjX4oPZ4RsgjRrhG
r5ONRr6Wf2rRBzVLTUg646O+u+1g9u+/dJkBYPu3ZeXft6NW98SpH3ioaa6qFkuDX2wrO/l+zo5N
80CB18S0MFr7U+DzPj7yRlPNDtOQVCuhSQHVT0q1yupMFA/DRJrwBA2qBmMd0gZYaiJX3ocJ0UQb
L486cqdUuWpOsKeoH3ELUhB4PxaIRSfmoOiXw1y3AdMOCAXgY6Zv6sdHYZYBJ/7SNNbcvn86ppFs
cJ97NOXCD3qzNs/YiGyUFlTXCHAcl56gJwV7T6x+wdmPtXTbZQA/rAWpUGoVj4e8Nkajl3dwiww3
hWHgKjePqIbvNYnfVXTtRLOA1djLWInU8D9KO1TebjAAe3zFd+lNBm2rGIPZqlKc8g6xv0OBSINS
VE+4s1APeZ/JNdjLixbkL8+mK8t9R3vdWvgM05Ruqf+EuhFHGTCInwLlsT6cyIoS6xN+t9+nddAs
uQJnuDZPOKzOVbXDNgL8i3cW0h+/S7gzvnMCVFPAHG9DnHeXwqgulryIMQs6en6Dm3N8XpBKCbvl
uFnZ1rS5x2ySEVPnS4puH3y7iuopjL+Ib8rpjrb+g4IdcaUqBxjprZKVq+dAO14jaPR8FvaFfR1h
48eVqfF3Q+0tgGyifXC3rBQe+XjqZxdpdNZjCA637mMfMbhhT+xaqH1Ox0qR5z3CsurJXWP8kxYC
EZfLIoMz++e7F38NMoAA20uD96QJxQu1TRtbiIE9+rG4f0Rl7fhYZ7phuAJ860zG4Z2puyb7afU3
SPiBCBQFizfWzvTLrOeqkXhCI9wJJhnUYm1UKVo47ZQmmCsFbhn1Xuyibn+vMF+d9eGBvO1gY/oQ
xztX8amWPP6U0ozGWVCJ9XiXWWB5+cZCt1EOFvpupKcLkUyjMjV75+94Zf6VhvuAShXb7v4xe3NK
VnbAbe3uQAb9ED209fSCHqcJZ70S6/0ch7BMU5D8yHkiOAbCT3Wy0TU/UZZGRa25PvXxN+eYpMm1
rpeUBiMXODwBHrdtMcbPDG6k8DORcMRi3mBILGXSMD79nV1JEckGcUOIaR8sAEEWw8cb6j8YPYry
QiQAALD78d82pSkuK3iSXhNowyIaAvmmreCIbuo2vf7HZ7GKZiDgtEfyVa8S1+feRaq48Kl1hb7l
lFsZN1HzmbEKii6xokk0xBiAVIw9tXfjMaHC3BVWdu3R/wtR9BOzOURmRMqBUDlNjLEMdt0pV7fF
oE1Nj5scgO1o0i2cSFepn0At8ZCxLHbuZRzhOoy4iA6n84Zp2EkllQtAnCqhoErnB0lYGcFVBW9S
+v7sfdWrZQMdvrvaA71dge3/nEjkOJEU08iBxTPIYFYIZYyH91FWzF5e1iB9GmgtnRA4Q3j6RZ2F
jlck/Db9tOrjiwSuYKQ+To7S8OELgfF9xIAeGzKZ0Wr0VLUneNKIZ8MPXyTJxIr6zI8ynD0dYvbw
MULdA5/NNGg7BtpID7RchtOO0gqBs1lPIwNDNSfuWG8UngbNFdXrg1f7+37NlAhiufxCn1bhBdI2
9IWB8/Plf81QSyp4F2VV2Wqe7WfzZLbrGxdnCBTFUvC3CtkhfjFw9FW6whYugmrCu9G/uD/IsEhj
kP6hcceYvuI+w/CmZWiValOcjLsIbmIh4y2wfkDQZqf+u3yU2MRh8OAMEqURJLbneMr1NYJ+ryck
+X4Pl2N4giAhcuGSZjJ6P/qnFlYQw9J594Rnp2M/G9/iBQ97Dc2LSGrqfLZzDbBIPXQxpZhZmGKI
eV8dS1idwSIcI2jwd3gAo98laaYE/m5pHgFUoDdHMwVC9759JP9drh+P5SPiqea8xGtXy9U30U1G
8d3pGNMotG/BwL4FWkBacmi2U5pg5bgi1yRSXr1qPCP5gfCmmtdxeKX8Ibah8ZwpcKxgD2gk5T5U
H2lFwQkLSjktJcZPEFw9S/gK/8Ib7TM8ImRUgrqFd9PpYN23ccpt6YSL3BCE8GJlYaJz+w5jWr6j
eoJQNSasltVjy1rMJlIsMaWpDZTc5S27v532RTsogO3Z2f1ziZjZ9IqNNJ3fGasQI0DjT4bkuvIj
3MOI/+dMl8QmbBWA57JUHmsg+KNzDX86i7PtEdQXDUN3aUPYbVg30zqC/1vGTnfcepOI9hn/vCGQ
5Kj5uEwMU2Pjcs6LY6yMHz6lhbbyL36xpXVi0RL6eIA8XhvMyYCJ6iRYy0+QUfwqA5l08NH5Q4OR
sjFo/ylFJ/wkPuRGtQyVmJH+/cpThwIbsFCsgQD3UNJC3dML7rBjF1374C6z9gZGt4rloI/M8WnW
MLQbx3UX6/a1FjmJO96PJaqdR4G0R4ipHUti2iQv/7RcQIos+7kKYJsyraplA1phQuUrASzvS/aE
AAvTR4F8TDtQMpkwiwH/H5PN7xhwoiOnZ7s/F8tu9o8TnBt6/kPh8bdKnQg53awnORbPWBUKcoKt
W3vZxNMjuXRcasFTg9a8fO2xlx+ltr+OjDiXwZGTZez6WEEF0Uim2dngGF5sLQNzdZi6NHedB4V+
C8pboo2AAn+Qo+u7jmSlLm4r6S88zanCferYe/CxppUzNNgDOqyCgoO3WPDeyaa8ohrPfAKub0J3
fx0Z8COjhrC/EsI16p0qnBRZdXrWP7R9ISzQyq9yRIHJAdww7dA27HEanfS6wfYoDVGHcicDyDgh
oVF82cDyoX5yTxFdn00yPiDHIZW5o+DdCmlydbz37DihydjJkaNZu/5Fk76KnJj68zveb/OiR1ha
gNvdyuNI9AVsVdMuGrERLA63ASgLdjUE7EcNHqjqTs72j2iWDsT2APi/ua+LYzboEpB1VKvFlkW4
wYKm8RkHbnGZgAVOYOs+hrHOw5QIljHOdC2c5W8NgpslTQFAAUGeSjGgFbIU/Skntv4w3tZZurQ5
my7jdMKi55+FHHhyEWs9IAaEMC8aU3nSQKZPGZI55vf8pa44UxXdCgO7lLt+YCxE6U3VeU+MYsrD
HMQWcJ9DGiPS3TtzJavWlwj/ZDZKYSg1Q8ROj8AG+zoI8Q4cjnhllex7niuvsYV/8zrl993tjLvy
mysxwRo8XiuY8hKIYD3gJpoal3szzQTG1NVjd82HgkRUEepJC7T7oiO+toDaoZEUChANFLtrQK0c
+HuiwTxZ7iUcXlafXJt5W0pPVuY29x30gCj8iwRuK3SFgtGKhO+4diyOkf7qUEOYJWwpsEn6/vyr
W0GSl+ZRLJuXwVF9oS211p3Iqg6yzR3hEcBNHW6dyURP47Qs04iZ+m232kOUstNDLfwpxjaKg3ZQ
bS0ezbmI08+x11qEe0vp48FG8mRpSSbdJBe2oBSSAckfIEtVVpGN0QgxkX50SClNGjtyCVlUCVcw
Ay29HaK9Sw0MARqLiSVnBkUOoQPfwN4eIgkfJDQ2D4gNt6zq9kIh4YVjeJQuq3VoFyjWf+OOvchO
h+UGNyoYCXWGn8TT+5HIv5EoMgtkZA6oZxLgMDDKUgXy8AO1rOIRnC3eLDgkmMtQHVbOjQl/suOp
N0gHc4ctzB2iDNZC9VGl7X83CaAjbhbkwqYd4veMhm29qu6bmgPb46WZsKPlqTDo2xcTIuccE9JX
J8zdFR0rDZ9+DqmwwfG9EtZMoqmglF8Cm2oH+C80OJ51sPAmXIWvmTqt7KrG52/WEExaQq0fTu1r
nmdFqW7+TAHahL4GVouxzLOs6dYryQ27yw9JXQ0vhSHtErbwh0OpfZHLS1dMIp98LHmDRV0C9Zz5
EpwIG37BA0N8W1ekZV1ZvFoDsYwpzPtYyD8kGqR4Qz8CEV7ISa8Y9DQLoURrLCs9E0xOjGHUZo6b
bSmBegHrY4NOA2QPLaV6Wu90oR2Wsdot3W3ZOebMZTegwkPZl0wrHQxlbJJzqPMrewFm3DY0+o8U
kuq6GrxBaOE4okI0nEzqrVzdoZAUhtFFeMIwIzZuG+SFfda4tnwfQ/bowIZETNdKG4mcz4ERNB96
oIjh5tgA9OGFdEwivReHHVmBQjbzo67M33VZzZchPL5kLby9INXmE0uwAmmm2/YvaKKHhfE48xRL
+ORHkAUEh1Txf/M71EiJ1FHB/JMauwrqBxju91Ib+WTRxRjm47/1ZBCWpIqMjQd7WQd2o660xgNr
jYeEHbF9RcygCM9E8WQ/oFB3DS7vVp600S0CcUCVhCyG9+hnVCrg8cCjm1q+XhCq3Ma975bjp/eE
IaTxytSJpxSoe2tGMfR0Z5TQ4wnZuZBfe6N3mqNW06OMBtIcu31PRwBcL33Nzz2YLVdVswqVynX9
ULeFiky5y+fW1oorB6cELUTKA9UGFiOYo71GlmlRBNxobVkJ3GGrV386Sg8HNgczLvl977drk6Wk
dEJI1taL5CpodX8pEVum7cHUJaqOGJRXsPcyT299xIW1zBVHpYoS2h94AeJ36gwL58NxgdS1I3/g
F7COwRlQweAI38KY8kTr4AUWIHdtYGydb2n/wdj4EpGNQT9J6mA5chm6xtb1k1BT73CGPI8tdpHQ
mHwsIZJkkhJXmSoGNOiMcYb65RFqEUpEp0dUi6SGKUdP3Xk2//1QehNYGScP/Kgsj5LafyJZFEQ8
hB32Aux+YUQh9ruIKEoCiAD37On6fstcY0xXW5XeHwcBT0/Q7T0tKlGbGrw5Uz7fN9YUa3iBbuoB
Ir06B1mK78sb62aWyNgww+oue6jWJO/2Pf9rkrWxi7n7SwC+lGU0Zc9TW4V/QT8zqJLcbNso3OCu
BmIjEorrno0c7WHRxiQIBH7bSM2EIxxAx4tRGQCUMTYIHH/8aC/dbqosSq9qrlRRO2j/KjptMbbA
GZtcpM3FPGpMz0h4fZWQeZ7Tu7mpHLbm14XWEzwL1CfdMvw1Z9FyUOIrwxeXtFH5eAZgAd4v5OZ1
SD0/PnmCEUKjFnVRh2jDqStLDWY8fzwpwTDFoD6OGBXkSn/tALvjgQPAAugOqZVx7dnSor0vX5Ug
03tD0zNIPy9SgNdXF55HHny778MRGVXwsSYqtQP2EjrSQMPa4DqIHLfObyJ9WSK7d36SnKdtxmVn
bkXk/4D9rFm+5gqe2ieYPb8mieXmbuxCtJDXHtnn9QpGDU2xpRaeVI6ZGz844ehe4GdFmnUcjL0s
WUxUaxgpthx0/Ec8UyY9vufU9+q6/x7Q4IUqczIVX9zwJPCm+/GTqhTPLxiaQTlfd4DrdSnA1qb1
EQcpIkzp9ZUJTWzH/CLHq7ZePu9oxo1yu3Gx796exZsP7aOXJIJd0tG13IkIxPXMuC8lQRXREJZo
mDDr/8fB17ilaAW6Q5NbEze9hJuv6QQTy2JmzjLTBxyqzSeUiFx2cPNGKoykV1Mr0ObdzccTbLt+
EcGlEEMzMPW5d/xbmMMweBkLq8HrUmahvJiueVFXWkVdTaYE6V+z3GwIKqSngVEgGfjaQoof/EuO
vsrjUv9l1SxzxsvkCTVOVq5Lfkb2A6mS1OJio2bZjgXpehakIANH3IC5fWWmAZOqq7uDHRZf2Ljs
2IsP4qV7OWeeiZWqLB8mL0NKI+7GnB0zzOmCmSYTgyqKAC6m2g8ZkV1XhKLF6k8fXU5hhcsxfD8j
XxheilYaddyzRiItGxcWcc/20ptj7gW5736lTXJy2Su+Tfw6mx0+hrGTQ/MpXQ37YnfYhL/R58Hk
LBUKdOa9PlAr8bo9QV6EwJpvAFRrGhjm5kdiYWYfVGCy3u3SJbKWITw1VM7gzvFUdVTce7mjAQK5
qe/bYGoh8vAeqYzf1Jy4D4awlowik/JyxlCEwmhbmqxEgHxxSy5qRhyJuQR5s/wZt6V/eutxWgTa
vDt4H5VvbpO5VXOVndhLQztejo4WTnJkundRU74rRMPXCpoKPLLlzKQN8hhVzyb4aUj4xhDlDDK/
CjqiMu7Z9sBJijhkjw+ieWMReqoJ9nVZhtN6J1fYLRzqiK6fXBGO9XmsHNP5wSifEFPLBPYG5MpD
jjJy+E+TwMd9ni7IYsGC3M7N2MWN9s7v8Xi9o2yORw/AER5eGTn8ua3mXgqSirruhdq2Hhhi3XZ7
ZFe3A07zPQny+rkc96K4dyCkUVrd3iQu7Nd7nKlo/+gVpDpUZ7QCz8fwhFOJ35og5Dz+3CJBRzj1
KQyXK3/eY6AaSWS+zwG/qtzU+SuuuPdCk7E41hRMtWT/XayhG1WXUCzEX91EaJHZPvyKN9/CGfg7
AajGpxrvJy9yiVetdAFx3kvlgmvom2raCiTfthrvXb3o1+2uN52f7Zu72DgH2IA7YAr8SfsR/gj7
SpodcwdUgsRFaQjepQK1yfbFBjYPE3uNSF7SWN7sSwTrLcWyxpBz7KdV5cWDGeaHQKRhh+FBocK9
9VMW0K6AsXaVWiDp0GPznJKE+SnBn/2y6VCDzkPbG02NWOG6MyepE2phBMRiMf87x/O49YZFX1Ln
GIki4Ay7uaLeJozBGOs3qgdniZfHp2DcjYeMpbLVvGADZis0SnCnNksCLRJ36MyZrHr/1osjtqZj
gEdackAIPGg9TJxlJJQwUqLExRTTQ0jRo2VHUFj0OMt2Dawdq/ZsFEhjdVUYQnjhTKXsSRuzd9jM
Tx9KsLCNkZuQAiXi7xyfI7EmCDAMtERb5Z8jyS1uNONzkW4sv3cKY10HPFlwTdcJF1MQKUlccNWa
+/8ZYG19UX9z0CmSkJKcuSsHh1AVPVKWzcvPx8+Ek0Zf6Z2jvVm9vxmoV90yCOKUUOFBuoEMzMvD
9kNcpYYvNPWIW4odpDL1dF416oDASwxWFEP7hrEcX08fihQd27Sfg8HU4s8xHfTGG1zlHzorZL5K
FSaewtKiCoEn1t1q1AZJvKa4GS/myy/QR59imenTf8GQavuP3zyLPL5ZuNCtcI9D7vesOjoGdVPL
1OWduAm1FEK/z6wzixXSqyiP9087ZBUc3EFQGDLxONZNbjm8IUWw8l1CRiLiRv2G2RS0lPhZsjgY
wrnC/U8MD38BAQoY4D8nDak1aq4NbJ1J4lE3XTY0P2iKOGU9BgGFxxdCvDgxq+C37KqTQBggiFaS
6lvxPbkZwaOX2V6xlMs4zU+Cpe4GFPY3yf17vkZ3l+Nnwd6FwE0W7l9HfoSVEvT1BSyIhu/W98c8
ttw2jWvVtBiZ3OD1FckidYdnQ2wP5kRfprPyBoDgf2kJiTt+9Qx3wroeyr+51eip2HvlTpRTwA3a
AFjbj3t0yee1neYYsQ6paDB1EjDsge40WgUmv2zUEiLVN0704kx9Fz/ysC1WAIV4oJCGZhhsoZeF
iUbHmecHKBKJYHxY6HaJePHowKISuej9RnZ+NWALTxMXTvkmwN6kgGIUxokCqiX6vIE3q78eqSC8
XdcbBbG3TOle1dLxNvxLurZVfdbe6sWVa89rPZDHHQk/XykZ80fFOmh0nFa5+HdMbB5UZlra17Ok
Of1Foj+TFX4vfhsa+LhSNXjsyjOGfZVBCNvUVg6TdTreClanFB3e/pYYxvKy3DUc5FlN17GnKVrk
kzCugeKQ4DNG7xESCPG7hj/PtzgESCu51OKEMlYVjjWK+0ZsOF6GZypycErBoWISuuWjQkrdBD/V
Ze6pRgHoOlVovNykSm6Y9SOLoL4FOsbarHgtcTzYZfbxya2lFbfpxAYDa4qwx8hCClP1uSObQ2hf
xWB6t85HvjXSMnog+aNgmNioLFBDNC2kuX3PbM7DLn1sMdInc1X/OhFBai/ET6FmD+fUssikBQH1
y2ZDT+4weqTP9i7Hcp3pn37JZzeIFcUL1Hajt1k2NWwCqCm5nLRvhEeAx1BIImKRWagEQhCAHHtn
y2ljQXm2FXI2x+183ahZ8xDEj4RiW8N1AoO4RcNwcwuvW4+ET8lMtA2BIwJMxzGMIWZDsU0aW8GA
qmLbYpccGQEDkw3fGvYetfYHrI2mIZHZeaaTDtNE/EatLtHwkHI0QTS9jUKF25l2iak2ti5vpMrL
NAEbgig1B82qjPy0RGb2Z2K2df3j/JKN2+oe9uQCdq22oMBwJ8yy1qx1tLfTtNeD7E1eHyvEGOuN
6lgZ71KoX3QOELYVHXtIXxWQMa+yxO5VDDjepGJ1MdFHnaD9TmNYm3Vo40yvtnToeXBpDngLchuE
F35nqRJZPhcZ59kJ/bkfO48mDKKtIdL/upyMEt2y+t8KXhVefQySxiuKNlU0A7g2XR6RQrCxf05p
Ejs0KkHw7n3REb2ZS2W1X8w1fcgAg2JQ8EIGzVkRPKKVl0GRHYgrfYfbt32cfL051SaslwOgWbxL
8Ckri46ScAq3Lwl4qFV3olYAMGTlCPyiUoK2HOJt6O+kopeHtkgIJfCuzYoK+P6cVCA++ZSRzOpc
kk2ZfKxSyU3ByRahswL65t0qLeg1XpBL5e4ISVi1P02aZbh6LcL+Us7GgcXiy5P03jxj8soulQfr
x4eHFKSsTM2sOqwGzVQ3kH+YIfcUpWJIvJH44nxTplrF9xlGaEWaarNiPUTlVpBCfuZWOl+n2cCl
fKTkTpDBnH0dACxyLN8ZAbVuP4Q3z4UyGyBqu7cgxqWGV5kCXsTOmrbkemfLO5ix6dBTvkBQu2QX
URkVO/0yQGic8MoTj+rQAjtoCEzsruS2hxRttW9AZCgyj/5MNM7c7ocJFKA7CUxlgKsVVpAq6NmD
Z+3qi0twMdw9nQeam7B2PUjVrFOJdiskTAYA5sRuyoh0ojZih9ttLHip3Eo9DRN+qW6VywQJzmCc
/COp4qyZ4gOI9G5hpOIvALqMvKmmTsT82qe+Lz0mUov/sOo/EsXGgv61GB8sWSxcRxvMo4Nyk7GJ
CIHZ3WT0nsh6nsCewP54dQzfK416P+gTZUD25EKb7KxxUYhwkGEKdd+EQNZOjJl8FVF3SVKjeEFf
5ijxspvk+c0GTUvJ/YclFJZ/6HN1YcaphhhS7gs9RFYYrXy/SbsjFRUNHBJhwHX/dz3sj+32ONO5
Duk/VAJ47dhe+Gkm9chfQdtmynbjOjCWF1weonjwajnePIf9iTX8NWGmcT5k9ZjmTtfU54mf7x2J
u2IwN5dVvEeR4LUa/jep1bS6KWNLBb0YsGLXHyg5V7R8TbmElV4Y21yYQJWv7+R1PT8+Ky1ldl7y
oywPkRuRUq2QASdw3rVRNlX9FkjNk7nfZWIN4g6h/gPPg4QAiX2o+XwNp/iI4lhHZUI1C4B3m6ug
oPdTx6C469LXk76lQHYCtwPiBV3Sat0T/cfzOll2pzdkUfytWfEFyBrqSesYdvdpA94l3kNRgShD
HDF8AYjsYKM4AX8Z/YQotXn6I8eVCGVB1hCxPCN4I087sJb7Yj/ahSsEKfq/gPeWFRFtWAJqRdW0
olYYSNnml68/n0Cdbcq2rdgHQWLaVOfO6rNWFwB7qR70jZ2gJrAUVq2IXNixP7z0wgXA7vHI4vgq
nvxebhp2IETiDaxs7hpnOXGzBEFlV8E9QXmrUFw8XKywgzO6Sp/BcYERNGXq27ZHK+BpGba8ayR7
2KMHqY8yqxpzdnX3hQAZmKincblMe6FNBSuF2rxGcyh3lD5jXCwStbUepEDUbNt/QG64L1q+8eG/
OXWn3n5+PlLArQSKzUViiLNgh4FnRcyFv5e2Y3F2yPb24lQq+No61yhNRGIdZAsswpfnqdb1mC2l
6eujQSWUZkSLlm/z/evdOS2dnWAPqZl4aSw6RAdOHotssIItkYD7a/0EvM44Hbscza2S3i87hjcC
Gpw2c3Pyx7dN3tIKjg8Yw9O0y3rrKprZPed3qnJj2YwSsFXcscBn/3hDiUN7iKfo3IyPuSEVoUqJ
oYXFqfPZYivnQ7HTBM7bIKU7yTGFKtp9jrHgAb3VSGaGJdJwD2PfNoBjtnSa69tsqJz2VMAlYo+8
2jclgSuMy8p4TTbakQpz46uMxHqyh5eozdx/7gchQTTInB0jNpYOCdvCYwZzis02hEu+BheG6CTa
1tPMOyU/ih1UYEf/MpRwPnGakdkSzl6YSEGHMHeuHyka3cBaONt94aqTx1duyCe3Ja0RDJMUaJTI
NMY4UvKK/FpTvbH+0h7KWsgL7zldSGac0m+1cc5tSJcnpNDCLijaiYNH/of1iEsIkV4qB9FiJ8kn
H++tE9Uws2rjrgp0P8HJswytCBB5N0YU93GDwxKreFyR1ejyxFsuyVxfJtg5q2yGi4mT/AXhRw4Q
JdAeUCH+/d2uBizhovw/8C5WSq4oiZb54JxU+eSGJ6YDSQym12OXW31nQoFxYFT3Q1bsk4qQlEB6
ZlMGiiGC1mJpdFAkIUdBESpj814z7sVc3iGufM409p/SlUkZe9y7Onu7dmV2ZGzxeuheopUXTNXj
j6ruVNrBCJUNT/KRSbbI6hrT65HW1rmRZaHq2R9AtqWZSq0qbHIRF0GLswJndrFeQZBgPD1qQgpN
VJzDH7vFH+KD5MZx9Fd83O5JNDRl2K+zfA5IY6znhvXVyoSHp7AurmVJmfotuH6AzI+VZrs9T6Ab
WkbM1nDLUQu+n23pTa05zrtsbUbJMT+mWpKXpPBPrlMsohmBeoatv6WuWbXR/Uq7Ise7cydA7sF/
Pt/ooPSUccZWCDpX+yNkwQHqGgcMxZr+48YtFIgB9UNoNc8a2LetUTNuyjtsB3qwjLUcL5tpdO/5
8c/t0P3FDadg2U+mGR+BFhytQMbF5nFAvDt2oOKboT6CQKCbwsSWvlbP9ixdkNrf/MJBu+02C74w
VXV2obAAqGHWayZF5Ek8ZXQxjj9f9R6ZKbNc4ktFUGBoBeUPWRsvli8pGTHhj45yyvMbCZgILm9J
MHEmJWp+FF4f1kDBs1gJJ2HEbCwq0Z3hikx0dEAwFTJEvfUUOansAdJlT0UoOVm1HN4F+BV2AL0Q
uzyA8iyhCiV+H9hxkIXKe/wAm5sJHSvOvQhmkNYJ9axkQJN3OsR91YdIlGKFhqXo5UqWk42vweyW
fNm8g6kHnchd0udYrRpNYEVW1gSWEcx855FTGmz35hI+n/ve3cYXxTATmDaVYpQSmQasFyBtP0PX
U5jQMnxYSz2auvnxen/aj26jigngLcaxpJDorbNW2g1HXJBhLDlN7IFp4gKveYu5Dq6YSevDR0Pj
avv0y+OP6U9E9KIjJbOgcN9JrgoY9n6UxHatUrvOV4oVuZ0Wn60BABzktt8MjFm3iK2YWJ2PQyw4
E8ZuGZvi0CY5Dozh3KplJlCS9zYzg93hwKhlff2Bcs72Ccxk3D5OHobkNLo6QerdJbtQzSuPETE3
8IeiA0vF11XD3uBVCgrcIEaSBZQYGDXonrJRwWEnMAMbdmZHrqWJ1aAycVtVrVcM8KsSDMCna0AL
zQAoN0gEVDLaSDBjkJGy6m9NezXwpz/zBOLWSlk1nHsUPsBEgkNo/7pz8vijhDgk+b9w8RRFb466
z6gIC0voaa62j2R8/0+AdVG+eb5g5u8DJLsZee2DEBd2DZKz/NDipSzOwscK9VJTzUVp/gVSK7/a
ncSFRVB2dUOtVIYf7fI3sm/Syy9Alls1poJtzqWqhFCgHk5WzXnqbyU1ZTM7U2KjPDzyL6bPLnpf
F+9UV8pZkrF74seGh3lFxHrAhhkUEEz/+MXfesxFu4y04eTxWMaJiXlNFx5NPIxV13ptbOjKzy1w
Z2nHCl61BXUENTo0zSoSUVzD3r6cAlIpPSRH1YETmUkn3q1MHFr9KgU+Gy9Pdl+OV/+S0glDWpD6
LiMco04W3OLNtoo8AlIl8FjLZwa9GiXTmlu1Qumnec1OcQVrBLdzYWkz8luN9XWxA0+mHMEBljp0
WUsKHH97cc2v2ngan5/5EQykqpvh86p5pvaF6ae14ZPOlB9EcwwiXdhDV3NuERJO8rNhJptW5AJ+
JVjKjqGD8T13kmhQeGeEi5QhEjYctaPYbxowe0DY/aZRBKPri97sBRRlkMHiXkMdeTu1d/jjaDIJ
DVNskllrko7M8uyBglx0hCDcKjSRpqrPk9joYUChU5+4+PTNHQWUmtnmB/bruAdlaRb81RulvUT7
liRUJ1jwG54iGbljUB38S8IR8NBVzZkb4mCm9C+/0ob83vRGL1Jv4yGzvoYVfOw6tL7NdF//+8vn
+RwfomBH1qomjAyxpFIXtwqoFUPmqNESTEYLnWeQ+TGpgf6vOsJgIZzb20CVD1GpjMJmdo1UdPe0
VV+BST43yvcunYWsGbJXJMrNOlqTS50B0L85UP33XFX8st1tgJ1Wuyzoh4MGr+cP97IAq0e7c+nR
Mf4eeXUNJxdQzWi+aHfzAWWtMm1ZcEXutufscgW/6s/lquvaTggnWDKCdk1qlhjRaYwyu4Ij2t01
P26liLC99GRYvEauEjhQG4C2rSF4gy5iGW2N0fwj37Rfa16ctP7l3TPBvDgWU9DttnVHx8ifW+/V
U+PoM5VGs5Mbbiezka07fvXXteGAu0UzusVfhVUq6a1ghnkIZbdscLrBILZ0JuSoygU8toPXv56P
kilIudDr0YtNVY0XOuC7sC4+PY7UvW7yVx5DcYZREIkSLaLeHoXxkv/YhQpTMYmATvTRAvg3kB2Q
DcxJUOQtZT29hXksF/51vA9H/GUZXnfugEyiX31uKFkFscKei3PhYRDpqpvp1Aei74YIaGjWb2N3
NXwqAFg0haxtKQ9fINtBXCriT79sic0KHFP6g4eY724k27701S9gt14pXzlgMj4ZfCOcFinT6mKF
iOk64L7xnslLYRJhf0K3R3Rj0iH1LoPab6ZuenXf7xwLbe+63OPSpsG80SxTzq7ppCgTyQ9fNjeR
I4v/uh63zIyrZhBmrsCcbW4wjhygGu723Ohq4b3RxQwR1QVcNGmK1X665qePzsGR5gxxmYl6XsPI
lr8TGyTLBj9qu/S90pssHwd1dIS/Tjgs5ppqnd0G4qdfUQKY8b/hakhx2yQjwAK1/O0mQM6AhSr3
BlgVANjJQJ3eNu1JdBrfsnuYrDDt+XGMGrvLmbT8L4LTYlLvWt/HtyfjQHBPQZ/8S9KTlit/dO0C
0ZTo7LBYTfA+WoVkaeCiJXw2Ve0zbbgKdqi3vlLz7jFui8gEZyfD2ukLcETHmFZOpmdqR3sH7ids
8dH1rUpCgCUiu77kv/Tl7a8yth1Lw4Um+xdEAD005wN7xB20e2mi7qShODMgd0+u6XKqYyMP8Toq
SNpSQhIW/jRUEKRpgEUnx9tLH8lEktkI/tTOzTK3labbTv48zZ848OQ51Z0v2QyZan8uIoQCgzUu
9giqBN/F+s9q7VTwxyWATUtfFdJyqqWxX4IFTQy0KzuPJKb7+PY0sS7leadSKD62m3lC00BSYcBn
Wykwj6OAju2JA8MFR/q54CPObHtuq5Aupq8NunU6KUJFWUzfb7Vga77VHxyg8PtjNeR4E+Cw7jAp
YJFyG92Qmlh42OlwQv4YEYsIqAevIYzwYDL4jsq3JFv2ZTHA20/VQQd5by/aRn1kV/yyAgqNrqkV
b0s2IHZh7OOyZqDOovhEWX1v4yq8S37tfBwp1QSt6MNiDR1LRGHogoha3264BBn2Eo4gKQueDjOn
ksEhG6X4mXjdlcEffXBX0yFjp6YFXZmTpeme2C1SoCiuMmrwBLu7Mogr22/jAthEQO95WNxPG3Gc
APtfvhUsYoMTm/Mbb5P5oyKiVKUrMMn3R9pwJucQ2J4XQ3Qok3skZpg3MZIcPTNHEkgOqHMjQBdT
zkwrPNRJ4GEAfT3nFIvzUkpy1kEZUfa5439wnCmcx2IzeQ3HZxkQOO3wavl1Syi/6buu992qaffQ
r0hs9xZig3ULqB3gxPQ5r7+rXB3TTEOTLLojpPiKwKZH2WXauuiwxHxG/pBwQQd1EyKMrbcpzbJq
tWm0Zg1EZkqueXGRob2BcOafm/s9T984jOYtYko/Mp8FoFp3OFt8RoUYDQBCHMbhqhciWRRUKpeX
h/8/YdBKxUgjoFrtlgp411McVad0+jMneWF9T7o351NoX8uLf0jse9Xeg9IFRp5BU0AZI9dFugHp
Ix5XFixL43floxrKMh+iQkOlkqeEhZTVzwhgpCBGappIfkvqr1Ww0rlSapTLgw7C4EINJRKX1iGS
vE47LiPyrq2zygOnFRnk6DAbnG6KP2/NDLyV43+ELG7GgEdBVhbdn72x6qe7xpyLWNHOvP0shWtb
8gEDEZZp5KYQECmGLNP3VD6ruvw0dXGdKGD+XWG3Jh/rRx7rNF7H5159FQ6c5iC8w5ILxFgPRLs+
U/EM3aqB67AyJWP2uTcCzsU6qGhomJ1yjzMvfDAS+BldAD8ftJfTR7kei7ZT1DmfZmWgRD6eq6pG
YnsN+k/0vsS8237ZzMgUXyCdAbl773vTCUPjn7Q/pXWew+uypNqD+mhrfmLzHD7UAyDjgfDd2jaM
0TyVmWZP+Vaxko34BFnhzHQOD8jK4CTz0XzP52IV+x2q5Q4hhLTPt5LVJvRXE/1OixnT99RGFpnX
yct5SAj3Yq3eCZC/GHqbp0gvoPWDwldJuZbDg3SciexoMlMaoxptPasuc8CFJsX4ri5nbqHK4zlx
AOnOfzO/WZMFQHuVUrmzBqaMqKu2Au/6wVO/s+TLl89mDdhJfJOPcu3krFKAGM2zBd15rLgyCTl2
C3uAaakeHtBzv7l+wPEE4jFfFy4NfYT8KiQv+Xhg7IPo7rzZjcYlVroPeR8TkH3b6LvPbZFilnzo
fB+4gWkBkxWiNAwFGwO9gb6x56MuXXTtzV2c3gbPEghO/u4yqWSc9EtVKAFNXtwLRtRHn1b4Gc9a
5X6KOTuOHIL363YOE/j/e8WMzym0KvS3UAV4Zhw8uPap9RROh148va2BgxkScd+Zks/AbaHnckRq
86YwbknuZTvHzJaZ8O43NjhRuqXu2QMr5/0f7HWb649/rozA2l8HcTOfDj4rejYoFEv5M0oaPfBc
AZcKSOqos9rkmokUdkt7GyfUpx3orQhVd/mX89aPs2EDeUCaWnSPbnteErxSkR0By2vwja+SkBmn
oDDxheUkys5H7auGTsdtobVyQdvjnnLjr6Ohr8PoejNXreHsWW+fSvhxtI+aDiVoDsZzdBliEq+i
OEiApEnjjvIiMnQpUf4HDFzA4y6JIkJw1qPEV2KDffNamXYuCuUbVe+4wLy+Oky/dFB9m+8NeZgZ
XaIRBPj9n2cgr80bnS0kRUi3ScDGm8S3SZukIgLnXuzO0mod7qYq/0wzZrk9ddcQ0gFoUubVS89o
H8LCQkeeVyVXiRXuL+mduQMV2tnOIrtTd4dwMQhJ//xfwUXJKWP5Hk0YXtp3VTrhf/+zuFILFdPX
Muibmbo7BCEd+1Oy69XNRJyBBk4jwhDfFgtkM6sPbJONXaL3PbrX5a7zRYQdsk+IYVol6aX/IRwj
R4voYEmfuL8v5J1I1QEvmg3AdU+Mv9L4Ic9Ew70GHR/VpYdvx20u7lPUmlDhhcBjiQeB7zMZhqwC
RO1xWnKOugWvhlYtxo0VcJ/bxoajL81BN32wrGwH33joRwR8sdO4r3qnHk6PIsHOvOczWMEFBVm4
xI8K+dh8TzPEv979jIT3aCCRXdZuJXYgYEFE8FPlqdvbl6i9ekWY0/IMff+nDs45Xdr4iLU9EI87
ytxKVlJuGXFOAdHQfp2bdM80jxsCZzO2sVIFmCSemQWDVl2JxFZaATUsweKLTaY07eFjuDTQ7JRC
izSjYUsno5g/5TzWq4mv4cqHn1FS7Qd3Zg7oJ9U1u3VqpaREwe16q+JX1Z7hCq3QX1ciV985v0to
2kGzvqxmCnZi0yrXMaC+xE6RblY4z+8IV8Ui6Lk1ZEJ6Pv1VlSQxkmgI4l9pYHYFWyYQaAl6Lvu1
W8HkNJ5vGL/SJ50gWMd125ASIwfbhK+GWtngCnzo2p/q3u0gThbtY7l9n3btVNMdLjXpiqFj9Q/6
JUDJjF0mHcMf/U4R7W2wisHudoZCOJnq+qm664C1Y1xPfH7VDHZEDrKjLKELt8yQ+M+10jRG16u2
YKmirRRigopSB2zTzo9WUMVLE+FrY+gzuNGw2on/9HxFlv0jTmfLkKXmbap5sdzXGHfkw8x39qPC
+J3Tvgt713Xjmi0vpzXGmkN49IDCD8nSP6W1YZljBrzojDNGt2yusXBaME+Af8zjYkCaN1WgfEBA
HIZT8DSyBXR7GctIWd5dEKfNkGjAj39w9tBoL/sBqa+TfEZSEz/udzj1DQmwl5TZHj0jXPATl6sN
1a7yjKDhL1oEor0pihK1bWuj/JTAFsJtr5wBFocBwY70nnHrMgiT7FfwPs5dZ6WFZUL3N5n1d9Nn
8LmMms23H5BjKlmQfO12IZnowfI48rRqrZKU+8v4Jv127A4BydWX8NYS+feHTXGSLSh/BBhZYrjw
KHN7m9NWC81trhVDPhh59SpKxDyT8+7VO9CQfidPssDDOAWsqTHIJp6wM1WB73O4dITLsGd7iehs
vaZfTvG2so4S8n+fNL2hXIEG6ZQOFCZT42oiB6YsImQwTO0hZvfDdezPXoTP5YaCPqrfn50JNWVn
zHY1UGDamTO1NdasACpOh1HeMw8g0/qT3nwXrgEEeZj+iOLUjV0i0b+bJryTipNcvIYKGPkNtcoM
TLJJwKY9zDMA4PrMCXABeulWJrQh8GLjWWcWq6Fx2NGI3oTBG3ES/wlpiRRIMcRWB0rRqUiRRmtX
WdPqNbfHBAB7Ek4DDjGLpQWOak/JHFTdPmjBAF1rdtkYpQ8aZ0jZVxLhB7QJV9wOnwwDO0Rvs/pC
2o6p0nvcMTOYB3lRxjIisX8LOxCPijIPfmmX1zqTXxzD+rR0Y157+5DbXbJlw2O5PuhEiH+NaOtH
bs6qK70qVxFbUOfi+hpCs4YwmxtkfmlO4nijQUGPWh+BUF6A7xL2T5iFSGtBVjFpp0NTBFoEVi+T
MwD+awZ6BsMQud723fMNg1sS1QVngaDcSVLyLWjsTa64WQ6ALKDPpy50VvZegjaoYRzgyoLEUZE9
ddnZKHDqJcjDa3kCq3xQK4ouJb2VLJIJyxK856bsZp+eC3XRdGuXcuTyA/fEA08HvDh5GG0eJVJj
97ggX25YmCCyYRQ5Xx0PF3waLPe901RP1JffFE+qvz6eAF+T6wF7eN5Fom1tycIB5/WAjZCs2rOj
tNdE84sIHYMTabkTejgTdmxbJVimKxhU/452eTdY+Wp8nIGuVdSnuejL8pKNxBpiFgH80YiAcEb2
M2Hd1ZhAuT6yw2LdDxbMnOdt6xGffuBOw051LHxIA1XLwFDWi6C7oPIJB3cH+KZ2UpTaz/241zNj
vla+cph6Jj5cIAxWYSvl9ojmmlLdgQFzc7oNC0SVFTuSIcGCaNtaFYcNR6V5aj3r7XWLYb0sX19g
UFbKr7eAOiDCAX1sfD1dYeYKWZ8LcBiiPRhpmOjV4uC7JV3LZMmVLAc3nlOAHbyp/kZg2LzEwdDL
W+GeC1A7/xo21+DPCr9lkgsC8tiO1tEt6xA1Gdvr5VA/v6J3p6X644XA+GUcieE9yDQfFpD9ZF1G
jwJBiM3xt2Viv7rX7za916vZ7HjwDElxMgos1Ii6NsqPTYO8OdXcVwEI4R96LEDb5tXxSyB5dmbA
MhxhKwlR2Eu4tlLg5ODlXshumCiRDPGvjUcp3NG5d48ZpsnX4x0JC46VPxCzSeYVAEscP8MyA1Dx
FnnRczg/6L3qSudBujVIXtg75pXmQ34nZCvK0gpBuMOjuayD31LAsomWjqA5FdbdbS4AptDn2Mpn
9Dbu0RXkqrzfxRFseAoBpR+My70Psx5ogQokbfD/W9ptFREK0GJ4JD1WnDFqxMO2KH4RYxQ5gtqF
inP1zZs3qhW+5iQlRm5LFg8r2seRmLI7uZYpbhCalgQEvUcof2Zsczuczmn23hlyn0dVwA1pnINI
Qb3mAYu/3zMupuxMHcNkyNcNTWAVnbgOt53dhmEWW8ABP6YrUqFkX06CUdy0XgPoejfq+0QEEdpI
PBDGiJwZp0cpjzKYdMnKtePmD1eFHpZ0bkWYxMyHDwzc3MuYbPk0wraKmAEuT6hJPYyEKKJ1qQLp
n6Q/Ubfy7QlnU9M53yZSMyIbcWCy/fh4gYtVECHy1I9/Na0LAoxKpa7GjuNvQwmldfnA0AQ46iHb
TSJM5xHnR8vLcHp481ZVQ66zd2rsbhZt58QCUP84CAJ6psJeIi6fuJIGFnYuDVsEmFqX7+gbCGd1
mWjw6cjzLOXVv43gyND5bOQLSXfDjgowVoUrjx53cKTvk7U1p6aV2vMv5N/ah4Mp+SbBDqyKrdhl
JMuGXOKK0nTvd+rE3TB6+nVf/r9RRATc5+LjgJCvFCNJD90SOjiFjNohMjBGgREqXTtcPN0tu1KK
Cbdg70ipvBxJ2PHaqj8hGtWf4vvbHTpQvXz20x3ldXeDfJt0WUOnJWhkXSBP9k3y+Nxr0/tRYgB8
Q9Rn1l0Xf5p0JJkZyrQJJHF2+LzKe2JU4RbZvs+CFllJSmkOa1XeB8PbhBLEdMWJRjdYRm1nBEfU
pGA/COjoqf2BSuCNsj5TBp3HVvqVivyTq5ireBhnf0MufBWu4wnezjnFh2HtRFy9pC98qgkx3lg3
IGY8GlZkMybk61+vEfNpGAzVOTkF3MRXus+rxE2XZPneWY34Xzen9+j50W0E7UMoZt0cIon5ls4r
zuRdr1BbW8Nkq8r2tkhon4Ea9gN8D63Y/gE+7Lmdn9tv5f9uR1hoYpRLy0yGfR5sci2DTt2+prL5
EA0H/bYGPZZFQbFm+hArJKQBMwpM2ETwwiIS3zfAvNfeNPRjS/kymDX55TJqS99TTwQHSoJrkh0Z
Fwys1aRyomDkxUVv9nNNm4Iqe/fnO2RCDdyRw94Mn+Ot2EvFuwjCQS0Rzmrfku5Q05LGqy0FpuAb
G3luAVsfNrNbT1aMIdGnPGkR+F6UBi+rFRiTFhEKiKwAwqhM7IyFl27dQLIi+ZbA0gvx+RkW5Zoj
lmoxjrLw9ntRjlV2QJT+HAgYU9zNjjGevOT25eCD+QqsYLkEyI9tOXnbqCFfCqju0+gkc1HqtuVz
KtkFVtVQO85BxnkLBnRp4NM4wsh9M9W1DByUBb0dEQOG0evkhySblCvuiH5wDi3LacMUijEBR4AX
fd9QvDmGN85UrFAnEs99wkuvFXLC6+Rjhz0zyf5SXGGGzw4v4HfOucAyb6FfvrR4SbQ5rS77Z8+Q
XU6wrxsSZho8DynhmaVA3niUanUKC3HK0yrmTIFbAuVgn3NonAPgIlEQtV4T9xUXirQNMU08aKin
lz/hXQ0Qlv1yQZNHhBfPYtgyu1UoN8If/ejKXD2AlkVL8fBeJRN2fEcjh175SK+Xs+IcSszaaqoc
ip3mv4NWEsbOgkingdtDzL1Aut5mfhYyiGqKNG4K3MRcxoLQfWrmqPYHHYpAIuHOZLMs48KN6qMy
XHn/dRp2UwPG/0S4zezmZhtL04iJA9V3NYChYSxCfI+CPxwMvs/8PEXTrn1iTuFxPsd/RbEcclRO
1Hfjx9P3T69Vhoe5pOzwRunjYb6SdfsXcwejVzQRF0tBburCGtAE1iKX2kciQU2HQFkvNNywbqBI
21iUq/bA9lnIYE5B18o0Ta1B6Nm1D73P3HbfyGgD+NjhgULZuk1XY6Ze5nvjyrwNB3prYXQnKu/t
4aM5nCeQqhBBsOvbdp/PXF/zHtfks9Q9R+N9Pv3IHncdWwaM8YN/4p7Aqb311CawDQ7kuXKWgshe
h7g3CFwoKLIHaG/mEu5fSmDd8R0hRK9GbXX1Y8mCVhjWTA13QBVUm/Pahh5yYcvMr3lnVoHK1DI+
79sTSYfqd8JE7g8Mesx9KmDu/Yt/uH5doJCPdRvwTDh++M+D8fhQOzq2WykPgvKYntv9Su5fgvCZ
gm25C98cxQ0gsine9qQkVjxTZnSh9r80+VEYFgq6XY/zxKDLvC+d7TgLjdFPtju31E7sHhqiVzhy
PDX9hANe79I9l5lPkvJF5D7u5PQKRZ1a+P5+5tyLHd4bLVCOdLZQH/1rLV0ibXtuaDH8H/TpEjcq
5M4cXwtAcsKyDKXzkp0oizWziizomxH+6hRG97J7Zq4GQc9sKE4INc+QYfCkHulFl7XjUychtBQk
VixaXLWelwPn+YqoJGs5kdc/JnqkOeIF2HpNIgM8oVRggHlTUZLiAFomUMxVBgQXejdIGVS6izbX
hFrAj5yT0auxBt0LLdfmP/3A+QXW/0YtDaH7zm21+83uLzg2Ooi8EfAsaY+Fac4k8MMRRx+bF5Gp
9x/31aGCMkdmwYj8GtFVaXcYBAzLV6Bt3QXaRObnSaYhjgJvpaPvKAdSmCjYiRGFF0Se4Yt1b1fj
nAxREOFN1/3jgFifrErGy96Pls7uw7beKdwI2jglpGLwN6MS32BSM2VtkFZZlcAN6f2BSQAYZAMQ
EL30+m7MKgGV9p8BMZ/9rtvvZKgS5VIRBQMdty+OM0PskuhinCCLDA6QBqE1Y6kdPxUIgtVB4rgV
TLBLU5c/fjlS6BTSYxUr+IL99L0fYqOgnK1phmsp7uOqYj0O6fV9ISfsnrKkWdyIEqb2DeJ3I3Xa
NGIRjqou24sVXz8JQWVQzE0fiOLoUqf06ywTYIRe/5ScLpLYWPtKVN3UieVXIaveL5RThxPKiewu
maR1JzVBiBndf577RD2RTr9nWtOrvI/GabGp8jG8srfAVE1i4hOD9AcAwTY2KCmfTIubaTHIqDHE
hCem097quYcZyPfQLJI/wjAdUsUjVDIlghNh30m0fFaoMRPTOvf52PqUsI7/sj+8yVQ+eA3EzF7/
QxnouVYfisAhV0bIgQvvAgOt9d21jIl4+aHI0ofVm6Bl9vPXJaDjA5p0VWi/WkiMEQmEdiZq7bSK
Kj6hIcyk+QzpHkereJslb9j/jGnnIc0kD1ZYSkba2vYo8cbD4Ufk2XawSSM2OoQahLOWg0wfhb/8
bCY3NwGyiQKdWMQB9vBf1GfsZNBxyj39082ojPkyZZMmYVyLWF7MEnLZmTIcsyssMiJtiQtySuKx
1u8BCgfT/1BRevM8Ou/GeiHBubAn7zXyfky7kt00eRWYL0RZu98IDOMBnuoC3Qabhtqgdomi9b/6
bDZsvtNx/L2KzVWbZL08E9YPBFkKo1qI0pYLQ3OjGs9+UDDHVRGTMFL8MTKfEzsh5KRH9oAf35Hc
qahEEpHI4uMQrrokOhhkPxZcapaTuR3pXrnCBkepEy6V7UfIDGsqzz/FGpbEylbuZMjoJ37JP/YK
oG4/3ROuqfJeXwFXFArtIAspBDU1HFKct7r++TdYrY0Odt6eMzofpYaYJ8cNMCs8BGxq8BoMCR8/
KtdF8AzZb4qiMyUjAzE1g3ymBAOhAu0NZ996HTv70HuBCQyemNX7Hbmk6N2VqZTZ6yzL57yD2pwJ
b2CGDIz2GwDkmXhQ0YL2ZGY2tdJnjZR0PY3CquIls+e4+mK3maXF+SJfT1LCZEzuJyYyWa8JPyB+
rosYua3PETmKPX4nskFOSshsx4BXuPs516DfEBu2gs20DqU6Vtxm9MIkM+l0zcKAgIQNN3WamBdq
s5xjCgII2iO6WBspFXN8c/I71yjhHNJsPp+cXrflG/vZuBX6ShhBMt6z8iSfljV5AKSFYcgBdwgO
oegfde2JrOPXsb7DTwKEKIcOth5jWGLCeit/OMDg4fQpUm7tmHTQDsguoIqlFHctZ25XBBKtjebp
JZyhJ5afsuphX1dZSucZnB59Dq8Vb3whVtovF7Z6ie9oR4+clexgErmw95JHqo5v8i6LoJBwg7kD
/Yk2mioZrDs+l9Ogp9FQkeYfZQwWRIM+leqi8jJfHqjseThNr5hwceQfn8zpeLp1J0UjLarvXZva
Atyzys9tsmQBx5ASubWHh3ho0q5v5l6kge0k+UX1cpNykpXFgisiPio0vSXeszgUa5HX0dRQaaa7
xuMbAFO2dJZjbeneMFwHnsmyTcGi2PxBQTt40MHXvqpUOeuCep8HjJ1ysKY/fjSdmrUTkGOIS0uN
70vt96hVzoj2nOm/gC760ZQPmYoyRDGDIcj82Zm5swWj0hUSykkSPAubVK1uFlNHaqT3ikqY9CN6
U5HLTl+2njhV9EX7pF9bbh0iVxNRZMsJPDPMXoUyKjV7Kg+22kOPQVoF3cvrMdqV/zwiy5ya7naB
GpmMu4KuApEgjDKTN/uTFEUUq5evu+ry2p5ekO34CwxvopGUtNUfRkwFxbT8iRdz+I6uGIoWND0o
RcqJdNVJLzxVXBJHyFEmg0/9+27X5f9iUnEATPjdxsEL/7ErDsNJ1h3Jc/ydHqSlCFudzSIZAd7w
YNR9duL//mWkFDeZBDXTHr+wuAPOvrGVmvoyZRl9fNd/9ezlsRb2kUKKywjdqukh42YEtb5xtie4
WQ12YvVRXsRAFoiBQk6BouCEInCNtBD50C5cO9Fm8YERymYD0aRY/3vLSukTZJUBW7OOlHKxEE3g
BNtdhpB0OqUwOryzbIzFomSX/b2DwrlosHdlBbVuRd0eJO6U4hI6QHbAeFmR/CdJ9HvqdUc2BT2X
lS3AQAuCSg91Nxel1PkdLzBPaEd+V6/YIlO0+DN6Poh9Pvjt7TN8QTgsEeaPdAUqTFpZwvLaoroj
vjFTWSR3IRA0k/k++V8p0glOHlCfSO/RDy+X/sVW61X4O3wUlMlrPu1nsHLYs81skTdz/ziZ9iEO
Ij/1Xi3vEPNJ3YHc1UaKJkye7MDaQ9fdXaGBaPQxk9Y21z3DR6p9lK/37UxTeyDhEZV4TzDBA2KJ
KjY24T/tGpXYm1yZHh+k4SIe/M1lCQn2Ls0iHbUG4c9wzKJU9AKzQXyaQP5BAFelE8PxdDkUFs9E
1aTE3wJ2xH09hcZVw2NAlTOGNd/U27DlV0CGz9Y07VYG7ctnJAWlnLPhomI/M8OdLniIES48TKCl
U0f/6kyeHNLFIBTdR+0ec5X9S4UEVXxckAbGSazNjwiX2Adqi9tsv725WliKknn3ErSJgLMUHH0+
XaferYtRB1iwCZLn11X9y7EXeS504+b0goN5T/ZYH8RaqdNwRdLS0iB4Ia8QSDpmvmKVf5TN2+4k
YXUGBDA70z9rUQQUOeV/fReHKsfBAzIh6EPPewlAENJe9RMFdD3fj++n+U/E4IPBg/hd8bROiUIH
ekXGvR97+GmQ3CDs/+X/diBrLcAUgqSEcqMApnrIciLjH8VQ4N6BRZDeDJ/yNBd0r4zqPBN1N1Bz
GlouNZpy6Q3G+y9MtbrDqNcU2khG2XaGE1K8VhWBuhyJLxdPeaXwc1rot5QrxrP7GxjWw8t7fJjO
7ONnZbxRiWo9eif8IpaPPQKpR0+u7QT2CQ6b+5q8j6L2Ij5e6r4Elqclvw5FOd+GFk2wqO2Nvi1S
5tQwYWbSVXMXT17pyZWTHFXVyYcVsDduhmg8EbgJwECuvWM8MeM+aMUg2xZuyRN+K9rcjr0PFiiM
39oAk/k4B45eBN99wTIlfny3kefJWqMzdQs1WgaeSp/Tr4JmnWxGiJ9ti366hPbunXMgGwvEkffV
dSKZR1i9VhtSnQL1HYbUG3hlH/BzGkwaySgrsdQS48EXPOl7wRFFMVwdIetExBsBExtkqxJf/BZB
olJwKmU6aAiLXHRabSrZSxGcSQVeE0jADiwwqAPW3VrL17+wXUw1eKcQX+rN44kk2kxB6DyENnBt
yg0cx8C62fs3XWJ43VfNKmdHk/gCWLmITbBV/E96CzRIO/Inmda8GQOe80OG3rI0wusmeXNQfl35
cQkfT+EFs9WAOV7Ijqs2I262pGuaE/86dHasXB23bNZl3lrJ4c99s/Pe64V1iTic2mOCPlaFqGkl
AdvAYE/luXq6xhFjO74sQpVK/1R4+QYJcIUbmW7piGJH5oPsbmag4K4NennhBC1Jy/W43DYWIu5I
J2h2hscFcRYow2FqTybzysCl+8QUggreIiXPXaDwjZ07NVI/5aTK2p/owXfJs3LMTkJ4Dw2BmIQz
AjsHtB15DSClsBdmjBM5a+zdmcC9cqhz9IvzFT03y6c34VqEn/4R4XpUzx/JjoWYgBWRpcNvAmHh
caQNRwwkti2ZztnOImFI8PK9WYsehfbz16WjAMQpPXTx3vH7Pgxnuke9zqNnqLPoUG9h0xEuO2oR
g2y5ByQK8BGw26ycIhzm357mClOHg6vetx5M8wJR5GoaQLOn9Htv36TScTbFjGOlE4fJURs9CmHx
u76jHyRp8NewD67Eez+tiatknRyyakcGu7JijyQ4BZkciCVlnaNLoCL5SUAoOB5IlPjyVVMMKDzR
eI6VIIds40x4x9uqyxGFKJRMJ13YD7pOXbEwtUOyRDXTxLwBlD/Q6GEQIxr9Np2vZXoa9hjKriSy
gWwLPRklBW66a07meqqeVMn7s1I2jrAcA/Ho1Yi5eFO/vGgCypWUmmiNj6BdwN4RmqxdpU6+tgFY
GIP7MYly3JI6iPJlQfXp6cZ/McDg5KalUm4cEwPTfW0NT1WClNiRLwga8d1s8qYBSVR9InTbNPNP
Q0aSpvUiJve3VZEHvr9/twwfkeFBxWRSunmn0KttGrNAhyc+sVYSI8HIRIfNZLj/2kSjRKYd/vNS
nVKRUy2glolCM4XZK38yOV54gacfBvUvINI1dSDnydlH0DX4GUZGQLD4bH9EQI+WNhBYDXc9pKF5
kaPLCuayokRLtR6Ah9liuIex+LJKDl/jRmmb5v55JmnOJjOuK5qBMHzVAHk3F5sE4MsHczzKx4bA
TW8aIZ6AFc2cWN5z7W83MkAA/Y1hvQpDHliEd9VZZOTdy3Z6ak2DDWukNj1Hb64WpNgN+kXl09W4
1e83hVT/TLpkS2nN0/SFEZNEeeEaA21dffT+y2/aopWbhpBHTSTrYOH47eVOgBJ/SCjtVc28iEvS
jRBs+GQ4rqtdQjIL+ygmwwsJLwAxxtl5lO8og7X02rem3oStYO1o6clg67iWRqkMO86qkwbe2pMU
hkcJvAbt1pWyxs11EzjLDi5v9BVoH3Rvsk6DmRnzsRCtFCnjnJoIZbfEZNjssavW+69Una+9inOu
TkbPwAjz9O+T8zDOM2eXxARNWkEkI2poiz1l0n60dUVogbAdjDEkqZVqpViG9OPDalxmKa8yKRRE
5roL6CFIeeM8D3cmGfJddiTYFfzzKnYZCp7T9lm6deqaGha3DBQvpjhJRaep+0+Km2eF9LpT/Nmm
dN3HAJVAOuzSd2fj5uS2SitW0g4R1pZkak/xmlLibQuDUIey9a19sfEUR1KAfMFCcOCqTxUm3xXd
ZwE2RSs9gkBBG0jaiwbvDRbVlvYZECICKOwkgCAMpttw0kbTZuZVMzYx15vqp1mLvYbHveg/5g4Z
CvZJZsBGM+sXPpZve8/bkfUuAOhi3iLpWRScd6FFKe54ndSLqIpu7bq85W6N+mQvGYreSrHj5dau
CpZkd9hSwxVyYMNRfaZznU9cMMqwbTKRVEyF3OyiH8OGNHgzoEc+E9A5r/woLRvahWx8snznD8YC
4aCV1E5uBlzM89DHlOp02SoMosQdltUJb1gHlpbJRlt+nK7JMjjqOjSBahgaYZ8icRZHYTM2kqn/
6kVwZY+OuODCSSaew7GGnLR3oqDY5k4dJA/3tRzG4/RS3FE4JMfjGpaCQA045AYDNLhbnI/Ylm1x
2YiYT4I9oIJFw+qKiC30ZPQI+sigvuMaC++B+u4fBPmBR0F0vtBhP9tBS0SQU+2TOJdOMzQxnAsO
LAgCktebXBXc8C/cyRPP+ME8FA7jfS81K3VuwCcbSZnh4g5XdU4RMt4K1EqLO/vq3OLuaQqcPXvC
Ip/6A1eZryywUTvFIvo53w2vAB1IKZKlU1/Dg2tXE58ueGjw7Cf9v6RnCyGpqxeTflKkI4YMPQGD
xQQBlY0B1vmMuRCvOiQxQi3QeK6lpnWXA3XahtoV/pkkY0LXxEo0+sGPDXpEBgEOMdXi2m+GNEcY
xPzryS/J5CAgTmvGUk+rmHUZIBx67E85KoIIxuBppeWRcduvFYhVy6qgQQ698R4+xKFYLaSpiJD0
yaWux7G71kO4sZAAUHFLMkmJJ1ElmpvLZR8ZC/poCgvM1dh2X6aD51fOnJD1V6HBrVKGmsqqdjc1
oS9qjMPBrPjomkoSEok7w+JjKsDG/EMXBOVhE1yde+gTMnNPnqLWoWebJlL746aWprPQdQVw06zj
D8McocRXTayL5MaGd+C4sfqu10jf8H38j+15rk2Wj6Nb4SmtJnifyNoJdUC3OhmodUP5g72gpTmk
wrUtCcRlPiFJXCvP5ZE9cyIh9LKcH/g12eNCY56Qg6plZHQHrRVHY+In7Chk1eq8i99GHE2y9RxC
aX8WMEDtpd/0TAkfuyuyGc8BykWIo/6i1ks3MHFKcWLt+PecfdTua8KsZXQuPrnDENco6oa3rbkn
RSuvMnsJyyr74U9gTzfjlaf79Mo9eNsT8z/9VhT1/lTXj+y/6eu0bMwYjENDoEAOc+5GhhwiyegP
3L0s1mopEIciF5ZwE64QbrAcBaMWM9hOlBaRcqEGGrd6QZK7Dp59E0nAd24hIUMeXiElsPw7GhkR
Ir689BOmmRWiYg7EGRHAPGmU61O8tw6TAvlcl7zxjlm5okOgkBfasgo1CRcmIpMDy0Zn4OGicdYx
IpoAlJHuDA4K2cmI28aG6pBqkc2TBDIlJjuSobfFoqwMlDqKn+iRsdZtL4KyhykhwJzWwXi2jV5Q
tisIt9XDPEv2Q40U34aTBE+d/dRb67hL5LNVFTKy+3Ds2iIEpSXoczoPIMSCsTwKTVTqXpSmic5F
k/MaxT/T2wWUpVxJEpDZOpQyOC4Kj1DrTJ9Xul0B06vR8nbcCIYXvNHbt0HmoNcfyoTNgi31MM3f
XE9q00JQplc7afRcSKajRSXo5nhuiQIgdSnhmQei2ys3ZOb8anwtaohOz9BmP43fDrz0J8izqMBJ
oJdYpsKrsddryUBq7unY08dWitCfaX45u64bXovSZfcEHkBIzYFQf5FVqc4GdbLIJWecduIsZ8c1
2zoTKbb2Tzc/HKtc7uaVTaZxmYFrg7TFDBPInnABkfw2AFlU4a1kU61BJh9Ewz45qsDYQkI7WRN9
vuYEyVNudfhGikIs6gNaL5/Ktg+vULDFnHWl5Ayk7nGh7CBgJnSQHgT5pIGoEIyTGWWxIalmqGKV
3/mDQ+S01gj6KM2pd1DWz8I6aH6SGJal8Ne/ep4vvvQfWnN+TuS8vJb3hLBH010vjyOg1tudSLg1
Qk3ZSL+c3Wwr1+KUsFy5Ia+kKE/6ehapaeTTTjQ+ABNhLyE+QHtvUv4Uy8z6iPV0DL6b5ch2X+C4
pfWN/PyTXaFGXt1Pc5esgrDFFm/DhdCJeTZmQFT89mYqvLEVW1KZsdPf0PLXa0LE+bBvXF+CmY25
2x0mbO+tGBlAvvJdQHUyPlrVeI5YnUBcN3BRkHDOfhmhp2Hn5ciVagqxGq5Cv/NX1jc8rMwvd0Wd
0y9dL6O/LVIS/+MiACyW6AkFMxfz8fwTw4XXl+OPI37za6LuXWd4O7SZtsPZ/n81FFI0CWM3XYRY
Ww7CtHbw3P37udD/WTWCQ414yLMrlGmFnM/39OGYfW6dUi2UCyyF4ubr0uqwc9qbgfxAv/Sd3f2N
Az26a32s8mYiIeksKNYkhEsn34B14hyGiO5BWDb8FmYgj6ygx51TpI5aHQiaqsbmVZdcDvnNYw44
rTkxEQKWtgm1IFuKa67OVLPV2j1w6AML0bTWBrQ3gvJebq2+pRE6NhTfPlPdY/eCTrE8G8CDOQBc
GORxu4a6H4+xlO+Il/5X96MsCMZ/c5ClmkIZ6BHbTtVh4SGNU2zqI4aHYnIn1unZ67ay1PWAlLgG
2+fQTk7m+6GFYcFnsitzpBAw162c0zLbBuHm3JbuifWKupVFEj/HdoXQ4mXGu4bBpm/uDNalRxJ0
pcvfTxaZDo8UI6J2CcsnYTdvPm/jPgLDYmrLw/KN5s6VB02dBfEtGKjKIOD2+67gYCUcj9eLV3AX
x1eQx2L7N0UpTo1FzBMRPUZa8EcXbT04CmM6ghOQp35hOxKjVs0MlijO7pdQSp6mAIFPhuqctqSf
EfKmDIvSQMnb5mBra4fM0cZBbFuAcji9OLv2xQpzPOZq8QSrbshr82g5nZ+5apxvE01h+EMLQuJ+
R4f84dgz40OisD2ObKa2XyI3N0nrto9n3eyQdlylqAjGCSCOdWLryKhO9IiB40Bnmds2yJBqRE1J
RrJKve5vy7ChsI4GDoyMLRxahj8FHT7cPcXSsoAaTudzbckEV4wGEBJTbyw+K3QRAscJp6VnXmXM
qkiGfosJkhihyK7XqRAKg6UDEyCSW0hwsW3cMx39rCSn7Usd0k+jRNxDpqdnm07AFqcm0KTz/bF8
gdR8Rk48D/MqTq9FWeN3kf8piYjD73zPNsoDH8WU9MlmlkFYbtBKCAD00WuE/K52EdBQfidgzYJE
gdx8bd50TNgC7zVvwRSTs107nXPMZ5TP3u4OkxDks8bpmopoXp7CwUsIghzZ0wnE38qWR39yOR3+
NZkpyc3YGdNRqQSDW8gUxwj3DNXGOKBbImeMM/66d5L4RkCaGTIvRH7r3gKEJN0UrIUD1WxMS9+L
HOvNL7XHc5W1Gx5RlOjQbQ+fLdoJNoxZVkglhls1+kCGZMsxrk78iqfIBDk/vtXqBSxjPQD/Kpin
kO/+toSfhZUob/sHhXM7gJYKxr8u7m+96HdZ/qvw+cqzU5pjJDagWM/cRmcEjSb41YqVecVCXMKT
dfQ13aHaC5DiABcDJENgRLlJ06GZBZ6q6o1w1yn3td2ont/bZDqYoHllQ2dQoK+WqFZRWsjNnqfl
8d4IK7pkETQRuXea6WqpTlTZ9BuxwCeCRpkicNpfO6tnBI6ZxY0ayhQxpGr1p33at1biFfC2Cqlp
QhV2vEDbHGeS1f+ZkjdZaEi3B0Df6WrK2xe6JcSU4kZRBF+7JNmA73Bpzfvhyc4AUACDOuXInFXu
d833+RakKGy0BHTLOPp6X9ykSgtKvPAgwKSkGktMfWkekHfRpAR79z5F5RuiTQjAkgKF8wKUHIJI
SQxu769BJPo1D8tSQflyTOjWF4UvMwRWl7wTBnOuW8c+v758hwoIeit+jhUYhLUZfFJsulwtNL4E
caF50PnGxpvWseESBKDv5/mrc/WjtyHojT/3MpAWT4XEOcbOqOh+GcqHx3Wl+d+gultwVY9me6v7
m1JAM2P7aygS9aT9J/S2wZ4d+WKChNx5pENKQStVRIL7Fc7cHW64ti2KiYiDmTKgOU5OVetQoTm3
PSdPk/sye3xPyhbiE2Nk7KwNCSwnQd669gY9S3Fiiy1i+hhcRXK9Uylpq4YPrcvjfBuMj4jZvaab
LnXZD6DfAlG+zx7wBy/lbHB/RxDW0zGoypIGjnDDK2/mHSd1g8947VJLoY/+YCfxL1jUTknW8jfF
r3IBVIeZalOLocWq/YTR6Re1tpCQVO3ermUafGiCW59Ltcz+FLBSIvPuuUsdB2MoAtshaqlJ9soM
2Pm2yGVAXzP5ZcKcPZ6gNP8CZnSrHLVSE/Xoj4CxMZd2ltvrIDnMKa8FDW0uK8g3eExiBKLFdSim
U1psK77hU6buC6rDYYunqkHztHwFI8aSX7Q+bMvY7JuKy/QRDE3AbfJyR9ecyPC4RQdSMjtvXw19
iLUGFic3gD4gu2NoydUevJ8eAkkFfvV5Qrf5Ma660j4b1hJaHFbmeOHQBeItO0mrQyt9fIEjqwm7
MSYCD0riFHzmKH3QlBgbuLeNO/XEHMZ3lwwopo0Vtic5CNVmcYpFXmRd/Wim5N7kL10IE4JV0wgm
rj2oqT20w6hncxDERDx6AY2lFChZQkKvzF3AAIsgALtfLdxLyHb8hKl/0AnIfFnThq6DzQGZp5iy
R9kH6unt81fIvWZStiy1haAQ3gW1EG1OjVsJbMQd+xckytSpejTpzwrQGCnYPhGUdFMVlVUT9+Ud
NA1mvHOrh/n4qtR4V6YsiL1OgIMC/uxi9HlVRvBIyYoDazo1kLzpMb8+rtrLoIC4Y2/LVNGOsZS/
GnX3uB5cptfiamw4JmPwXIDrbEdl1ZX2sikHcK+CzRKXi1rlwUq6AmTotXA6VFy3oTCqTraxm8dC
8P76C8T8UKncuoytDigVhnf1tB+QF2q7Y0zFN1jKNZ2hIPtFLtZLqR2lyqRoiT7uU9TL7pdBd+mk
vqpu5cUNc85dL7GlvoAlOV8dYdyqqflw6pU6LOP/IjmzGNlswU//NwAwq4hOxzSIab8hL7++6INT
A0MyRdQ+xLNacgZTq1jegpWtIepdBRrRwOe5IdXKNNJ+h4OLWQO4iSw6tR2RBhPcLvtYe81oN2fC
g3X1qbFdrsxQ0GgKKHwvMsbLpfeLCC5vYeWtom3AFw36U4PVwQAHbbjzmLbdpLbDNCndb64Eor6a
kKShKPcEVRfRyZGVf7wSHq8iQIlYEiDOVdBUbb6dXPux+TXRzCCnrnSPg4Mid1GSDY+PnopUHuhI
9SNK8R/gfpaiwyt50O81TKh/h8bYUKsF5wtjqIvXOjR1xO1MBQYIW5fkRMJla5+yjnPLxs+upXif
wgeMTNSq4c+/JC833rb/sE38cflrbaRmtRCawMQBrbkYC6UIT74UG7Smc+BkketSk6ctouyK3HX9
QNawcxquHN6sEjK0L+Kh0JhXERfRZb9HS0/VNVdTH5lh6XVzD1ebonhLS8bOefEGO1ikF/PxUMgk
/Wzi0UuoQGtXGpt0YelGSY072sJsxg+tLZ4BPtpsE6WdpQjQAtQZGQVxtGTJuXgoEuGtY456ecy+
uOqHo7MD9IcZr/kcOAHDGfq8kzEj5HF8Zccvvbjxbikln2Yc9ieFuKJ1ooIoXxzkZEB3bWr3gopQ
HralCk0zyvg3hIHJ3moUpcgSBLObc/z7Z89a/OInDpPRVnxIempHwipvKPHBfKih8aDl532vtruz
BzBmuHvxg31OKe3cMTWgV2Uon9a9Z7YO1MLEJ3hfKJiZ2P1qIOwHGqmC15EiaP2nElIW1GSmV1fu
iE27ua6N9tSSOtkoPhP9suKAZLAJHD/PXDrJLrJECCXM44LWhp79aqnIcWfaHG6uJFecaftmCqK5
N70y2fnvez+qlhwJLXdXtVKmn2Jks1qngvXcck3wjvQfmbln53u2XwxULPcaQqJ+D/jxdczVtB0V
ZEm0DmHqhjTc5VuTqLMY5UHKEIKx8ivUrTsXVT68Kn5LuNJ3SZtyOvw/d59F0gw9IXscGg9Arl29
UCbcNk9h5POiydJ6YHsy9/SOjd5si31j7Cfa5OhAmVbRQOzL15Vn1KSXOn5bPzmWay2M33bNQgZ9
g+SMRKHQt5DbhWImnkgxgyHhuRl+HPiVlXe5QqTP4E3A+mYoqdr4HaL9Dra8b6jm9tu3zBzWHhiN
mT9BbJSU5W3q6yrsWTId78J2KW9VduJZTVVSnbpVqnqmiPAyoE4cyq8+awfwD4OaTzLfMY9+nbIT
YmkoC7NuapGKNXk3QqbNdeFB48iNfTsiUNDxeOCLHDchrGKC/ZZ8ucqWRng6STQmf/cuykV5mEJD
x1Vb3wYOeAZmK9Yrh6nWxpyWkF+k3leFHE5N8vAFbJ3xT4N32ZhhLDCmnMWWIRDli2TG5vLDWRnT
40m0j/28t2cAlf8srhHIqiGmaQj1Smcko2PmISXKOQifTwPn0FQ9ZmcExJ+XrNhwIJexB7jR5soj
3TkkbMe6vIX7Yom+dXSGXyzUghV0R/67ma7gC1iPPxMC8iLYXn5Ln1tVFeoJFAEunmvdd0kRffOb
YlMZ2AxhI2FU5LSjYk6jQF+LoRRyYj8M2876ykNbscf8ZOkMN73ku7iHT72JDGBQdJLDS80QKv+Q
tG91APtnRZgeXkHVfvh3sAZL2rAkaBzcFRiiTUxhecBdFs7fxUmSX8Z26oFJ8B92gwDrSoKM47yH
17o74ew/150Uz8wLjD+bU4tRZHtR2SpiME4rKs3s+YF4CKAwWox5TjGSzS8WGWBFUhEF4Ngp8tWZ
ZoRP1t+V6vozbDyIhMmDC3LBiaJ8YwX/pBhT8sWnWS9hjkOfFQcNZ6syjJ+BaMLxPKE9xeToYlzQ
NUFY+dlL/KHeGQJ1/PERilV6IBuaIOJGioHpjexr5NU5D/ZwbBygqbK7p5ldbHpZwcuGbslShUZh
kAJlF16aoag67kI0BKbzFAAdkV4EBwNkUoOwuLOMNxgSRd0kD0jA935l/cS3C4zk6mGd0C+hEc9/
nRvTiOr6Yz401xFfKHh49mRG+tCGSD3inMwFGv30WbuGX6v3zE+vGuifvd7ds4Bla1XO9pLxeJ1W
ovy4lRFr6+U99f0l895L1tRcdUD57h9XCUKegSUuYCut8irXrJYVG+2P7+A/WRrXzZTekMoS92j0
HNoXDzZ16BYVKm0bM5MiNFK2xIas8ofJV/yFQG9+AbUSlX6kkStp/yu049du3u9OwzQQSLT8NLGl
W8A8yyvm0Kbly+924qO9ltgfdLr2mXMhcyYNUk6HOwt3LUOPhDkd+HBiD2Vx650FqKJiN3iML7mS
Of/jBdzk0hOQkjl0nwQn4NfsEoWvf209gSM3CLM4oqQPevt7+jL2mYPwXjMKM0YmPMnR1q+6kK+s
v7AmdMZb7IRv5jAsyjmNWBzv/g+Wrd7fwT+R1zGPXFtG3ffAlI2/13Fo6JFl8zHdYGgw8E3hiCP+
SMDl21AT0nb0YVIcaejExry+wAd5yetu0gHJ+141tTQXfodQyzrWgf1OlTA4bjJCP+ceLl2BqsJm
EfIN/4L8S2nH+vJKL3v1BuvJOn38YtbEtHSj4fbSvUS4qXhzhpY8bc5p9sm9wf51AWqDVzOsLikS
H3fD6PHlyck4IjkzpBOVg4yvicef7lRdXdJv9JnH2XPNK6inuOd4QMg24WjURRzliizmE7JmMVJX
kFxR6Z7YbsaYOrQCrC00VqBuHdOFMkYfC+Sp7MdmISJ3ohseGlQZH9FN825LZMa1oh0u8jjta5ix
CT12D6k9T+1RMS++uLnab4NLH/YBq8nDXa6znmw1ctCvIUn8aWFtB7UKRQyovGYaebsg8FkvJ/G5
eNdfl4ekj1fOy+YRengh+cI7mu3w9ZBQ/CY6Oh3qVri2v60cuRE35b0WyJBN3y8IJrbMEYYfN64t
AHJqo8OmGg5hcWHQivPWoMHx85nN7dlRv4+TROogW4LX1bVS3hqnsfX1Lknu4YiTiQ4aNLOTKZAg
p5/v9stDkV12C21m9EMa+swtlIbL+OZV5N26JlnXd601sD80/cikmhjE8FVyHiZa5WGaJCh+bIaC
KVT5QJgXPwWIPk5giCF+ppBbTPOZj5E0Mt2kpFkLICGWzEB4p+4lN2MbNd6noPtv035jHKw0hrfc
WT7uUyt2uX8eucFJPI33e1AFGtaniBA/B1fxyvroGFCw1EfZtwPSEKo6+zxLpsGfIJQgqCGpBnk2
yqOfy6XVnYG0cv0+4dIPzS3/5cyHrgE4PUiQqRGVsRL9vYhnO8g9wYW+wXn8/aCcffBRGG4iDGKa
FhAmbtC5s1OgPWh1CQweoPHjQ9S3zS83v5F9jWrgQXrrGlesgPmQrFiVdI6ArMvVr771JIbEDllT
uf/NVXTqbdQqinoJ2Huq1Kuvf51m9NPbE/3zuwtjYg9M+veTaIjjCpmPGOYehhkeXz/PNef6Ri8x
Y4hEv9Bho9igWU4vLKs1JHJnKkX+ZV0locSkBrI4WBZLPl+zXqtJgVQh6BTg46H8aulhcybnApCp
8eMIv6pgd42vXjidAhf1uF8YycEpiQSElVeskBSgBtftvCrEJ8fBA9OIH77gIzEPMejUXlQIgdg5
0em+800G8wZ+OQSPoiWpUSEZKmofoDd2dYJkhAIFQshgv24eAn71H1QxvxoFgKSN01DZvc1x6Yv2
Yk4fMI86E5dpx7hMC2KmW47HjACgF2gXVFCOGIMniWajD61/04Y7+qRtqmdHb1e2Brz39s1MZEcB
Q53gZTKtp6LdvRZk7VY0UAqjV1otgtIvwLWFC5mXynILg3SdPGtgiwpR3QrdnlyyEfnhVFWNdCpn
V8mN15/b6mf6ZBjJ8kY43h7vPKjE3RrQmO3dvzWfyR3z2iPA1sIhXVNRadd5pmgDrA1n5tHhBZsH
gnZmgDb+4yzHFvSn2FDyoUhID0r7F7Nuq4ZIQC/s1gASn2CqE1tB8t3utuL/jUu6UFpoLKQ0I7W9
8dASMX0WvOMQvXlQtQkunH65m/cg8vi7/AAQtHaAB4daulT7tNmr53pm7JEQhnpfBINAi33pSKUq
PJcSVNgy47wnugShRpHhQJXVEI5V/dHiyKqjv9itdl3T6G7xFtEt0DFjWrT5z7I6J9sIjXluB6l6
jKvv71wc9oSv7S94Qol3tleF2mfLBS9WxlC1HX9KzsiBm+XRDDeJkxYstGqFuoHTvTxju3QaVMvp
CWXCS8Hrpzvuy+8qzuHS48JwdWr2hiEVAvgoDypqMxlixDGjdESzIO6RFvMJCtpNH0BZI5Ykuo2Z
ub40Orkurg4cjJevnmksA7oxpMndGwp4b6sqYesMDb7JUcV2jjVDIdQQEupfq5C3rkKqmbeKNf+5
KBuJ1swL675lVgHoEGYYpm4afprobChnBw/le2qbF9JgECAG0c6f0QPB5fLvK66u/4sPEQJ6B+xc
W4ck3Wjt298mXJ+KZwVmM/PGkqmXm2fGHPnh0uJ2+7urPqmjKwjKqZZ9CKeze/Zldw5OAqzd8l1h
LNpqtoCBuXGznsXty1NWEUKo523dsKrKGNrhgx/gmlC0dQ3eUwhC4MTTM/Hju/7uIHDzpkTiunAo
ff58VOOnB05ECfDAdTnLIVqFBTPQTSGpLkKsEkuh8TdgySQJRkWa9cHMePxk9lFa8t1jwOetKZ3j
dL7mcG6Lr/0coFGK/9XkrQI1u3z2nWrwPWNejFVblIX1T9gHnD/xKK3cuxDIFLAV2AeoybAuMLH5
B4xr3uzEjEWxPfdeIrVkp+/y6+/C7TeSMCIstqO4Yy66eSvPIe/8hReew64J47awbLaGpS/XkwQ2
0TAnUhmIs010QLnk/ikoLE0l5JWXjk35ZFRkUv7JTVI1bwceYT3sVoLTiYN+UrUV2lEl2xQLIKXO
so8dsHZARJToKT6FUbGfudTy1O+CxPiQFY42h3wQurowgG1S2GhSQxd+L8wNYToLF+POmCqrjM2Y
T9qskidCKhU6LhWzWL6uXb3gyY8mORSB+e+ioTcxXilxWCIh1VKHS7281n8p6nBx0ZIPa+OPlwDS
zEUhIS5VqIUyfxjgLMs+tTo3odJ1DYwL66a0cUnI2vTnP8F6jUzI7sDvdKJuzA1QiDH3Tk//h/X1
5nqq2Bv3TQc8ENsIV8pONqyA1tHiZ1rm6W+KK/yPOaDS6WUHKumpCHZFIQSj6SHPn5Dimx3kgK1U
IrRHwGSxrvj9LvEqbdyXJ+r6YTXp/R9M4LZQjZ10jaedcwEM2Xcy73C7dQOS3OE2Pp7EkjhWHv8z
+acwed0B/ZqbLf3zp4CVYUVYd9KamW4bqpgQ6xSAaPoba1G4ma79pziRrMyAHbuxDE6wjzYcDmvB
bUpG2Mu6+QzuetZjCKFRBpU0yIdVCZTaSM5SqeIdpJDd/Lm8lAwGRPWF+Vwk95YkfXMubtysV3rM
0ft2QMmopty2QctFL8hM8/iQz78XtIhr3RueBXiezpcbpUp4Q4VBSbfRRj1489yCCh5+lZNN66XC
D5a9ZeYiMbnf/rDa0I9RD4Fq4+KD8NSRIYaS/y5QNI/XccdVN3y/klAD6jW72DWGvNMye4+XGBgM
C3EqZg6GEtRBJ2+jsCwsGFSWGOFbe1TdMSFfRCgS+uiAq0hX+baaPtuAPtBpJGMJyh6SWHoYzbOz
EX9MKZzEX4S365ZkDAmsxe5Cao3MXgEsDuBNgA+fnxqINOmhj8AhP7BPn2kWI92ssd56IY51m7PB
cVemb9QWzmhL9bLmLMAXfz33xT9qEDcB1/QWnXBI3uYqS1IRuT3LxszmtMMEF+bVf+5rSNnXWb37
996ld8G5EzzpawgyGnkSplK3YBWpKPGAjcDJ/tY61cTQhyBkBOOFHde0PXbB969pcN7QdyCxAMdr
9rM2SGtXJo69txJSo7fTbbyQMGAR2lPX5CfjoQ/RWX5BlZX5xdJkn34nwdYGA3rTd/62tiZPsGxG
a7TA2sexNac9WwTmpSWuU9kHO19L/hp9Rbi+TYdJ7V0J12AznBpJwHH/J2LiDHwbRwfdYSXitBxq
8Srcb+Yu6UE/+BSbzC9SpS9imY04NfhXv1NJ6cO0oUo5akaZDMm/E4A9qZSDj3F2Y8iC4BqtlL11
oCCqU/g/90o2uYyExaSkHpvrxHlhmULg+gbIqRAwePCWL09dM7FK64eaTgjgdl7dlzBlofL5rlNH
3N+9KYOsdYTF6/pJc89S/y9cApJoquD3VK8kOy7hM0iwT3gGqAtop/dpjQgp1EnEiZgTHGS/aNZ1
g5IaAHiQOlqk7L7+l3oLFfg+TsLDAdiMCRa1tTd042BIY5ZND32df9g4XDFJyihAYeFejz9HfNWG
IZxc8ILEdM3fXiD4zyviN1ouEGFOCVA37WXhmxM8NPoGQdeZVVkOmbZulbGjyYY5bPeH4Ua5tGYN
k/KF+oKc9w77EG4yAAAjXTbdsNRCYDtvbK1xjZgX2/NlGISF/iVdmzVhXP+M5Xvk233/fKlVm4uX
G8E2gphM7CqZN/gkaTFID4DjoKq/zseAlpMIU+nHvkyuanU3Vq2k/vBZKLXDgWvSyB8HxRtNWlVT
ml+PMkYnKD/yOVRCQgmIZe+RHPqFEPQN9R1UixQlCy8NMDJMw4YKc3RReBjfSJBfKqEJXLfFgguW
BsdenOZrOIyan4MXU7Wazxw3UirbQft4xEikuWpkAqAuR8sLfIZtGbx0AGIG8o3ddyZFWr//wg8B
T6wlpK1rxrBMuXyOPOYHT9W8YlJpZURaOML7nv4Lyq/NJIgEuj8XBIvRmvHFTtsbDFYyvaFd/NOK
IDCxIAQSaxtmPraUnAbfuO82L+f6ckfcsZJ2fFZZ37ucfwc1R5nE3ZbXMQVadaA5fQxXsGgS8Ea1
4OOv+gtaWj3RtYbWd7T9RJOYvheOo1Ge3PuskKg/R12voUtuWeFKCnJg/IE/Dh8+LnaWmGAAgwQj
JzDOw/ZcdwNdnOAyyJQJ/uG+LpHl4DmANrZOUD4Ma0OZUsrBInGat9eq2NCYrOvZoYCOpfCMptHh
TKpN/s6EiEsJpfF59Pf7cTDAj6QUxve+ru2dytxq3jMj8hSkddk6ZR/RRgs9lZ4FBEe3rvVEymT3
ABChHJOMk7Tl6aIlRLIbTY0op24AmJyhTTrq4kTpJeSwfYgmh2bgi0NTjqQJPB6C8/Mwreb+Sql4
F4nCV+VQWzN6emIprCNASNiea1Q302oSVklQluLrIQl/kZT8BBhf1SrzJx4taoXUHB71TcGh98Em
OaYjlMzUoIQfbxELMkgRz+XDa54JT2NJV1ODKpwwASCsjKIvAMznmMBKLlQxHFBX8vCK4vLxHRNL
ojmR2AECVqIyI5WmjYG0ElosdsK6UoZGwDjrywq8SgeJGBoF+VIG93xDHDoe9I1VvGVXzh3KpAGW
ZGBh2jKXRRaew6d7zybVL4hc7PEuHzBdQKunn1P2zwrO3tZUz6Wo+Fm1Es18KF52+MLck6x/87OV
dMwX1OMxc3OwE+6PX4WqdDDYtgoAL1Yf1CsdN19+Pt1kPfey1kom0pHWe3mnQ5Y7TSW6nZI3rTjb
BgWxIvOdCgWjHn97SodavFalCamFEKb81XBeRCYMrv1n2YrGSPmDn8O/vclVm0cIa7JeTRSXrPma
Zjj4sbnflvLYF/YLm9GeDYKbO3f9sNY0yn2VDECIjruu1T2af6bhEBhyRSmyIymYJLNzoiayZQ/w
MkElQAWc4jt2WEfDzYTcXNY65tAJaeGHOtjarDlcb7ij4QFNoeBTcieohb/BaweomP+XPdxyUhe+
TIm2b90Be/Ignviei57AImtqslgljWqZ0UnnaB/Y8F3bJPJdjqoLlqaksY0kKW0t63fFYbdLc/Mu
cw9Fs4MUFYlWJPyAB+xwkbfpr+juKsfv1sQyPy1sW9meyQpZTaTX03HLnMYFUgzwsvhhZNVkY6nt
akgWBN/YHUgIlwiTEdTz/IMLeyKZgKcjx5yd/rYcneIG9SVPeJ/5sf9GMSckygsDw4yJESoQF/pP
2LboIkP7TjD4mU1Sn/gPTWYIMepo8gcne5qvNrwxV4C290HFnpzbaUxHcK4ladGhcaNkuo9bm+TU
pUEG3y8MWCAUttAftaI1d65ak2lonLOjC1qLnj7KukW20Y7hqXz+jwPeuLAa48YgA5cAmoc0Kr4O
lomQM1c3dkI2jfYOmOjg3qKQr09Y/g0Xyt15sZnJfrpbGpfN2Q9HfRbGgVBoUuFfBZIbR1/5Yeg4
tVc9YhccEpSkdNkYxLUpKdiECa6fkhWuuC1SxwAKTuEFBO24cw2dHbvDVD86Cc8iEwo1Gdr0ckOF
VcNd4wEfHNoG9FO1O57cdqNJT7v6DXhYj4OtVdlCpadIFhdTWTeJtuJLYOtjcyfmC5qw8BPivjz2
UEiTQSL93J6fzWA7G8ET0EAQUXvfViG5hKt/BRgohe4IDDsF5g+zA3O5DRwyiK/OPtNemOBK2Pfa
I5OgmcoKYViG4fdtuG8noRnVRSO4MGN7p1H4g0VsipdkSRZS8IGxuyuGRECZJiarWIJPNMaEjFEn
8TSreAESAqKrH3PIfwF6aGIfYrVRnCimbKliD5sS7HuM0GWhhYwmuaYUXXgMxw1s0cZcLS4oSEXa
b+5nSOtpicVJr250nzscvAUHtUQ0B1St3ir1HdNl1lG9mizDmg6Clusl3UwzBDkdwnDeGfTK9HW+
lA0NMCejXK/QzLiKqAp/k/41h9mfXFzcFqSrjhawkW90meVc7CkWLuCWCJXKzXBHY3JiL9z0OHFk
+I8rwYoW9t2+zuFCcsy/NnjusdW9YBb1+fviU+Udxn3YROaW+AQMiwuwe3Dg/pq/wOGBUyVsDTWO
srfGVWIN15y7Z2CaJe9mebQKzNKzSgKEaonHLqQRTgHvVD7KTR3s0NgPC5iBNhCJg/Ovs4ap3xNR
QmG1QwTLrj4WVSzWqUbS//XjXZwXt2QR9NDpnPcMnKyNTPZYKzhs3uuFjZRvqKIywlGxxO5kzozL
YBubMEszM1klm/fPTGVEwwyqtnDSh96FK0W+Xnh/Q8DZPR2P87jO8cDqsagYtMc+77/ZHH2QJBje
5NnSgpE2xjLPAPSvzsl44PDwzrKFBj44uLu+bUVADOEPUUGY83y0PWX+wdTpGdh9ydPmFSk7v3Ek
o1Jvd+ROzLutt1iOpWbsFihaJAR78Ng3MpeyVTeVYlQuGODFgIIUcGG3mhyMO669adYcjpxvGb7+
CmJUOY9+FNtajCgcIk6Gbun4zehhUeb45OUHk3tW0XMHJOV/Sq9m9LRbdgLF2QaaKPdAGHGlvKcB
6pGOxiZk/4oWrKtfZCKz72+buKPsNBHC7fjAkiMvkJvjXZII0N2jJnf072aenU+Bua1kaGE5aDFv
5/KM/4D5SY+tVGLAlGfpIOYmOLr/cQoe/7nMv5fkRzPyJxJxqXmgTV9punBcyrgiHK6A4qG4IvNZ
5mhODm0qEbfbd6yNv6B0A8OqQg2pQmkD1VFIIACKIY5JlgqJPqcgJ1MgANldrxXSMJoCQVXijENU
0GENb5pjVCJUWUgZEr2ryv16S51s9fhmzyZJBh97Kiowffr00WPAtM8yh6ga8a4bXZhG/9JyW29v
9WxKcF6EBUWKhEDlaMEg2fEq0QAHozXPYbq7K3wk+63NsA9DS83wjSmI5zJ+/NXFqLNPytPoik+P
Vh2EhFd/4S/00Oarh5aQ6E+WzvwXEvdaGTxXezRf6v6KAVhMiBwncy5jKtHcdo9/zJj6JqCnsrXj
gZiIMkxcWwYDRtRPUCLB7k+lPEude+SkScQf0988Zg4sDE2LnG2a1LlmWRhhkN33WHvD+qxZYuBv
JjjqH36K2APPryB54NNrlA3KRzvxXJnFxmrNrw4bwI1MYZ7RZxsOXx3gEpXMi5GqMnAd4m1WqE8d
7qZ0Fspio/2bAh5R5lPZs/RsnigruQD/OEPhZgw0KCLCD/PoeCMHc4ULDOAOTpv4BgmCu+Ka245+
rsc9+vRFy3ptm5a4BE4jCWbURzUdTZ31Yu7Zr7z/Dtt8exllXnlr6JB5tmNVYQAYGuD/hTmSJOo9
yfYtTUTEJYD+61MiGyTuxfbRmHaU+y8i0A7faN7sd7tLzEaKG079ERm5FV8Oq0XoQ4+PQjyNhWqC
AR4bEutJDv2vdTcIFF3dwjNMM0umEqQzcbbvvKDjI4rmX/SyyX62A73zbIB/acPl5dMc4eP7ytjJ
P+TwcacrUn996aVnxX7y4JSu0KOimeAFJREKvoV9j4a+ZAqNWtJregkfbj+q+vZrOa7cefnGTjU1
lj94pA66Hr+AG2KggpYJXKzdLTQqbq1QibvAIuIN4nzLDn6dyjnyb4zyhTgVUtmcMD3bEPXCn/hY
8m1eY+EkOTauUBGytTPRP31xdhOq1XvSnlXw6vTWzGvIH2ZlzoBJ8mFaiJKElFALJe5mDqT5e31S
AQruoDM1IqQ3S94VdefZB4JFkw9kz+5ZvnZTGqOZ8Xjx08PEyHygP86wEft1Rt5OVBaoChpm/nHR
joL2pAUlXNphj3dOsH0Z/ESTZ5iBZJ7pnUbDzslD4SjhRKp3sIklgiqiRfx4PtSncZZE9oSQcUd0
4G0b7cuXwNlmmo2E+DQ22RB7mUrGJW/tpQgnn122Dht2pL6DzzKuW56Fd+XnDWF7grhKpyeMnijR
3EY/vK2yYvoypbS5W7dfoiWLQLdDrc7GUV88s9JenPUZtHPy+W/B6NylHybAJ7MK4Gmbu7X5m+lZ
oc8bAMWiE8Kfb6prOfqVEqSFamBapRa3sZWYQCJrcLmXSZS+Z2k3r3cLeVBJUHyqgdZ54VgKU7Sa
C80qQ+fIoe1AKWeGVAv4MWibKlPbJJOhyOOf1LUhUC9asXTdpyA6rx7IHy5BVYA/QnhMWBr13o80
0wB1uAQOSa5PpCjP1eIwjwXS30fd5mmDlHSpyrkkEvSaDVOVdBMNv2aN0EItfFEV/pGinFrVh+xT
GhWRbsEZLBVkmlDehai1NbDgoW9tvyN4xljBJz4zRm3V9uzqIlWVW8Fpz2+QhBVaTHOX9yNffW0e
SazaPGASXE9HLlNASwXafxnbqIFV1T2ARVWGfe3g2byn/gwip5poVliqFs0DnCNT/MKOqgigzfcn
Hj8HDrHkmS6n14OoN5q879YXR8YNOvYVsZ6B63oQ9OpZjoFC5nibTndrpyqvhVmmh0RS6GUeEKAV
CwJ8G2XGGYicxGKWLC2+vIDt9IY9IZffZj8R4BufMhUZosVauibNiUZc2GyTTl7Ec2gB8lFM8mvg
mhiKGChXA5enBIAqE2t5f/BNhFpRw5kIs3IDK7JWM1bzX/iik6MdBn4KWl1Or8Nwq4kIrp1Ls/Mt
/XrHvKGJpGDw+9z1rt2hyEQoBBvFNm9UJsOtKW9H3ZG6txzzlGsmsiIJPZMAVbrRCn6hzCoxPRXR
lqJ+JGQivpNMsnXI0RQEXgHHGPjFbeRA4ndWtEVVi3fFodi1qMig/gXofZPX5hQU/CnCXtDAl7xC
cBtMQNQv6Oq5f9/2v1/2aoGBKIrvxAKFjKajun5NF/plUtjAZz61b2v3L1F2vB+ohb3BiybxuK5+
q2FvAJ0DR4B4vXwRQJi91cPIqX2iTwKIm+9imKewx/3UysSHx90HV5a6UQGipnaxJaCbvOL03MwC
X4fu9Qj3E2efLSQMqwC2CH1sAGNe2a2p5CLC6mgPFZCCBGnOasLXORaVHZvaVXntBMhkqs4mJyyK
ddx0ZebWzfKUVnCGP2T2GsQk/RQNM84HkuL6iiAzuzrGHGOvwq4guKWsOhUYyu5tnuvJoCV1YItR
UAFoAe/jF75SKMIdXteT+kUMgbEf3elbQ5750fMS+PrxD82imRDRp5EfRVPn8AfzZeJ8YCmmZb+B
rMZ0N8FLIAhPkCnrqGhca5W8+H1giP5HBRdI8aV17MOom/lDvRXIQtntXkRnJOExbiTW2Ekwc+YJ
QyRbcMNPiaFva1/Vh2GIqk1eAtWxaZGFvljsItSrdJGHdOPlyVmuEQRtlCfXmEZfZVXnGGcmowKe
m+dtHKMRF2PYvmfVFKcGQHLHbm8ylvbKo+kFosT6MaIp3dBIVbcWj/nt4dPlHk5QwtFCV0xJ8Lei
s6355ZVJdCV4r1vE2JBFpsrPoqKVJLwKV2bKMU0d9vocSb3UienPNoSBRyYt5+/ljBSBdHoat3JL
xXzn8iC9Z4C/ffzyRa4Ip2K3Gk7eGC8ErMuHmfPGKx4yg2r56330+3sPw9Q0jyN0rEq02i2iq0vy
N2lnKSRHHBi3okYqiEVAg7ArPwmu+WnWDHi+zdmY9PVPH7JJ1f6CHAx0I1oQWRY/lgNHr/4v/bht
JRre8wJhUgS/nxkVbqf2c/87+uL4/ewP7om9btdqUc56udQa/m11+BIcagcSPUTSiBN2IjxTVN7y
75Dbwjx1ybdSNOa+y2jZvVG85jm1tBKTB4LASMlLaaHtozRA89dRiYfEYQj5x/6KE3ihmESA96Cd
SL1bdOCbx5sqJZmw+doljnUnufXN9NrbrcHe97FEKqiid6RbSqC1p7Afa0VOJzBLRgzJcXJ0VHfm
ShY/tHnAqxliGkUy/Gipe34fdTdPgjxrq70ZLF7uU+TwzmFDzyFahT4iZrs7HSub39E0wF6a1Mi0
xoua05m3YgQF+USCeZWOciz42H6AiXcySm23cedKLoP/2CJD3P5jXtQzqx/wBryOkYTQY3d1YxU1
zihZ25QN3iKa1lsI4QZNslwKdaX59SKVYjO/8cFRqxAesuWYTgwPBjN+orFPzV3r+KCuZqFP/uHE
9K3exsqRyL/Fm8D6NPZLxkcqZCh12WDtcdr2qxuyO8mTcXxGAO+5t+nGJKTrweGjRlvP2EdWbySy
cUMZbIPQOm5euGF/ANF8zv0hleqx+E+SAEEeWV9s4ltrx1om4VTylwqwNe8b5AYrNIENyDLWgqHB
qbC8NSQtwGqpBIfINBlR3sZ1JujW6XMFo4VxgQM8mbws4pduqU5ZieYH27bIidzgWhNXNhw5/FEv
bQs15NGGuVQChJIVl1RUzJcxzdd8Vp7F1iq3M4wMu7fERZ8qUPJ+q7O4/jewY2+ZJpgThMKf5DcE
GY1ixJQ8xmqVy5kwNo97uQUW49ehcOkiJqf11STIIkIyDIBuOXFDy6gvLOBXAsxsW5a5OMyMfOj0
dGChf9eWucWLQeMWC4qHJKuGgtkJpvbzQPkhrElffu+Y8jKSQjCwJMuOIb/qlCKCBIt13Te3ZPbO
dfYzZqbIRbI3TpDgdH51/AsyG/74kQjT9boJqLZEq5uUAE4mT5ESnF3loniWojQicMb9WXvYL7ev
rK5BemJoGzjS49+c75Tn/wcSd2Gw+Cvz0xVqAmmxK24BCP5KwxPFlEcUaSdy/P4fkWQtsn+pSxi6
csmGF26ivusu7Ahh+W74BQcoF26f2ncxoD/prkCPVI1pyGni98Onr6F8vbQNRX3UZ9j7PIG4o4kt
9WZGNVOaT0aVsbYKKtFGAS2j3NSg2/O2PcMolZyoVtuL0AVRhf9a9zk2bRHqQmobovcyFW9VFrnW
amRrP2qASYYvPWwcP+SJQ94K4vxW6HTvXKepT7SVulNwm+SYgZxoS5UTo97wNvdH7J//Th74HMQ5
ihtNkWuqQyR71sPY2Is5rPuJRvZrBZexaa79ZUCzwZs/9WDeF57UMTn5oEV/wutKVeQTNNlmHgmh
97yS6nVmTV5stiISycLIPx13EYWiyeBRHtxA62mOb1fjeOUD5tw7XMQ5v6mBb8xpclvipgXsBcnX
Kqd4Wvc39PEBnpSG71R9V1kGzwsHgh1nHNbgLP0uOrdUivKoTRtDYgTbG7kDMC5496+hepGqmG8W
FKE2RJdYdoyqlL6SoJ5FxKjrKl9wTp4UQYFb2t6LuheoLlQmGBYL9ys0lX9XHpKXgYHPpmO/0fz7
dRDvsgIWqJIfQz6ksFWkH0e8rY+Jg6lZgafdO3vUMiRW6qf8fJJQRlty/3htC+YiXN5K5OxjejxK
mnJpu1J7hvBHy/NXCDO6plt+6nHMgHl24En8ruwuLslLvwAdUzNjOSaA+P3xKfHFGtgLfvd9K8H+
VqqADfyG5dpEgMGrkUPstZjerJKsqQUC9h0HmnGOzt/wL3CTVaRc4G8dG6tOBupy/YOHvjtKI2Da
Px4wHnxQyShom03b8j0txq+DGIz+MyqW8CAbLApY6MZVAMySReViuvQpw3PInZqgIcptUNPrk3Gm
kLRTNYYhttRF4pHHzWLUuRy16zmaBee2vuot1DnSDmQhrbUvy7ZBE8a1tWvDLUWf0nE1OyEzfCRl
esUsj+EZpp8URh8E+nM2WT20jFDf/c8vECraPbYD3NOyKLNnMGNRLSVjlCmtAM2ap+ZyMT3FEUBR
+u8hpUzhFNYvDpBaM4PGKFJDjQBa5YghHC+p00y59JxtaSTfUziZdTopSObLMdobzcYiHrC2hgBM
lPlCe1xFoon5koi5PGWosBf+Wj3U84X/A2m3LKCd/4fSinGeOxT0pDTEOeHryonQYg7xRL6NAGX+
g81M/FD3MjmNHJ7JgskyvZFQ3TgYZnQrmtxQivxmb7GtT1d+LOIdGhmNqT5z8YDmxPZgLRn/vYKF
xIdByuCUxPftXsTw1q4DBkq9TFH0P87XaK3lnGd2XzoYKCQotvFUfzOal67CsdgJPiTTFZ2bAr7L
731AxkSBiywMQwEQBq4syz5baTjpsjK6Ied+qf6EDJDAC/V2kz5LA468J1dZRPARsVJBWYFxmSy/
nXVv437JddwKrwX1dMvLktB//5lpegenACd6mWAPgkHRLIdHJSewyC271AacJLkfCU96wI99JZvN
/L6ZzCNjO+RlzTijXAvrmhHieIWtCurBMXIhLHOuMEH/txLbYRP6GX6O8NMx5GErlDUCGIvEEhOK
c/y7NhYKFKdfpca9MhVKHS7BANhYchq1+TfCmIdrMyIneoIScmhAfyA11tQg0x1hT22U7W+zMbfR
AqtNpqUXPFjaWN7owHuwh8xEQq98dpPy5TexTWf6GNnLFXlRrQB/JnyCK9GiYygC0cvv2yixuUOv
vVSYrI/oB7uv5VJ9gz4FK+FaqhCbG9q3mBHy/ZErFtQCfT90cWSgmAEBgP86oNXIvZONeOu0/IRv
UVcsaDDfHkrrDBFKLjMc2i/XUjBGDSwcerrWmn0UgBL0/VIxiYVynGmMo5RyI9jmBagU8zaVeBjO
YltS2B6PiZYIx2HAGx6xgpPdSaYQ9L1I3sJLI8JActJlD0ROQNe7rLuL8W0rf5ZlSOWuITLoH8h8
5mOlMMuzzzr1pk8ClETqDHAAVbDf+efpUQBUv9NWxhB4GJkXzfb4t/jWa0dCCdL7EbDyACV1x2b8
bYC4/tuewDV6CbgIGpxSu9A62Bl4+3Ez3yjQzWKaXh1GASC7ji7xTfodqDKWX7Nnw93UKb5ph5+s
+dizt6Jh6VYm2quMSDHPp4uV6kTge/IjN0z9G/vwXP+RWTt/dnSuSqA+FNxtVvWPZtzpF80vrlNo
Y557z1TaTMbZsRC4gCHKHHRUExI8h7o6vNtLQ95k1KER8SbVRwFBNIO87IpV7+bFBaidM1dahYiL
0WB79GEybIC5Ga/S5Ma3tbp95ZvBb9Xi4hh/1Sp2F/kLoDc/gAgpaWmfFU5y9xnLaVdE/goUyiHs
7ReKuPIAhqW+AYcYydXYcjyR0LOOuIoA7TR8zhoQrqjg/HuRkHgkADIcHzSGABsDzUD5xTHN0gUg
cV94SWPWzLI/Ds3HjXD9scuLUsefUdMkCylmpD5CKlE5jAIQhdva6VB/PQGKbEoIgWvrrH6p1QVh
QaAM+rhbbBGRg0HogOzpboqw6ykFVfpc+/r+5m6q00vq5EIcMUeiRjBcWaJBDEnfOc7hmJVNhiSH
nI6ErOZizTbbs0RBJo91/4zHRpXuWNWAP+Yp1zN7J0hmiYn9nR/u2VX8z2xWmT5jruU3PU+QUTZn
flnDvjd0NvRovQClGbdWzdeSINlgnxs0z4aGpr8az1x0lxFQNv8L+lIIwAegl2W0CE4i9oM8AcEX
EE3FoZVXrUW5N7KdNZpQdBWpXIWfeSE2XpMpitGZ4t96ULXdfFLgekuYgwXvZtq3rw8xqLCCW5Y5
IuzjN1tkWJ7oF7U/LfUeHvjAA72Yywx0KOEXrid6cVofpE/q11w90RvP+Ap3axJ1kRMwmD2/qZZS
/djoZnwXkDVLxuqFYnFiQA2YnlSWORFNvazOBXLQIZRRkR5vZFwuto7fnQiTM9qcEeCw1+2c+/Ve
UN76UwtfYPlBWPrRgOom5rM8vD39tetWm+o2IQA7Jbg29MEJ3TSx53yDcAQLYy7Cog9mkp9dgBaa
Ar/lAzBczLz3UnUNxP8qysDEFTmExRMJ6DcnV042e16ZEyLB1Rmjwyr4C9ctYPW/50XPfxUijr5T
Q4Ql1z2zPEFIFw4u3kQhaT7HXljOC6wx02SQWQazlgeMlPFdtQ/P7jeIbXgZ945XM2MfsYXB1noS
VFW4dd+UXAwSEu8vOhg8t5TdKTGiVKlAuEpmKLY0yYW0atxDXmxs8BWUAgbYwISN9no/qGcOndja
5ZPzX543nRe8L7iq7GjhnNpGaxMR69ZQNDCh5R8mygQgKmGMHVkED/3J5/zSGIK1c7fdd43x08yI
TUpE/2oSvzj5uBLXjvvCZN9SpNCvV/cO/G/fW95UjSsS/hBCFFZYIsICZw4p3KpqvaLtiTD2kvmQ
Ba8BFqvMIhOyTeBAZMaJbSUj1+qmH4Q+PmVMz8FgZjHig5HSYFZrVbXX53IC90ZpsPdbqF0zXZhf
Qz0Y0+1LXPMAXY2YQTnz4g913BCeLHw/iBEibzCoDD4VPiFDhOQmayn2NAf7UhsyvkXoBmJ+/NAa
M8HvgBKQf2TWeKkGTDg5r9Fi4PLKplTyC0RW1YRHMFQy41CCri4V+zHU2fri6Ex7u9lai2rt7MFC
5pe0xO08PDzggjUpNm+QdTUoXYnqEL087hi7DpF3icViU4Ltn42Hzbzi/IJlaOlQBBpCKGhzMDMD
HxH53a32KzIgNv/xxTlHMh/f/qHVvidZRoJg/fZfjfk8eYXEjw0b9Q2vCQQi7/W5OOOYKpGfeh1g
vFas/HJ+vKS7Gnm5rQad2OmzI58L41eI0J8D8WRBQsCUPU8bTcTToB4oTf6z9kCAnpHFeVlrBkqj
s/Y7rP8jtRKksJDp/2Ut2ySps3+rzEQ3cxlpPdqIdVPVM/0eIplZTJ2nMgZNwKkQBxlUnUrT6jnU
m/y24ID2wozvWgEoPaJRKsp1MDIBd0zFN4bebLKlkR5YXui3YyGhaLyfFnwj4tFWQMwM5CVuM3O6
0T9p0pihy9/6YMhDKmjkJtzWVaMhT4pAbOHUWdwqRtkRiyksmOIDNpI8xiNdkBqwNOI56+cFWKwS
WOx5r/gHec2sRYPzksN1xu9RCMjj2wiWJUakB1/mFaqvv9dod+TQ4VOBPxcmGDN9UMqAhdRcJhdZ
h0MMCbzUBa4BUNX03sBq6U4iMBQH0+Ofnf2HbZjuo9JeqKDm3NGF0rW5heR9SFcKKsBOWKuh0ZRW
PjSX88XD+imBzMKoM1hVRWBYvdnoidIrD+OncWZDvcvmbUZgJkUoVHV91oKW35qZj6PvT4dfEJtg
0z0ccVYc33KnetfSWNz9MHZsAwM45p+hvmgkgmdRbcPZsRhc67LsgwHlfNZu/J5Qlx48VSKIZbvI
ZSoa3vFOVynY9gqp2geOQ4fgqGNlOomfzsg95S6GpmGwKPI42vMt3cbq7zyK1GYSjcqwFpUlcl3E
wWdhKi1Do4JynRWyfanipqA7s8NI0saznaQNKoRiT0BfZxMa7YUdyiXVF8gYolG5/CARyH+n4UZI
pKpNJGIf4tY0N69kp5CC7QTirLlhaJ4qddbq5O6K3kkPcDHqfHPyqNDU8r/a/0/TQchpBT7NLkzV
DAyicmF2IPtSs/HwdwZpOZblXzCsTts9TOSL6fEoLJD/BwIBi4Ok33+HLMsAP6DZfAauDYoAb029
Ph6wLrCp/af/TgFm2j6wvQ8jmcvpJJ524mTWIeq99OMeqfadhJFgOI3jhc71+qc/DiK0RF0rmDpJ
MCDcDOX2pCSarLVPDZ64yDjPOcWbG8vMhck6HZNZmvVGGzzECnkHBUEwRWioK+SfdlNp/mlswflZ
CX8UJGPAMEn3p0M3dq4Dw7NAIlk73cRPD+TpqEbtvU8grwhR1C5xqg+d8tzVTc0BwynVYPiQaacx
fTZHIun89SZg6UFGNhVzlfqRAfZeyQju+ypcORXq5JGCC7zKyGLrkz5fqE6Tn3yykykPwsO+si7K
hPI+qQjd3g5YZyLNbxmHkTubPdwA6LI9ISuBODmA7237ciO04U7irOMH1e2p0gKf/2YDvMDsrcGC
neZLF1Z51RqezAb7a4FGj5fHcerKlNUdX0tdbLw9ug3uUw6HLlYH76SKC90BTJfjs4Xld7XGwfD3
761cpLXE8XV00PzModuD7CE98jp+uaiweOneCaXoLppZtg+Lwfz9sCvsywuwiQMrpVbidumYr6vO
soUxo9/37YpL0k6ffsWlkDFUc7f5u2iYJmN8JH5ZnIPAVIB9d+1pqG0pBcdmYqtaK3X5nALpWB6S
hTO3+Rvtzs4L/F0YTRWCqAzAFxjBp1gxUs7P3YbD/pJMqpIjzfodzp8MFl0kiXaVTUXpBZ+5mxGk
8YIMVmzGG3WQygWfhGCOvO2XksBBEY21YR/Re23BQnE6CFonNuMYVqJVxAQmQH2wM2E2MP1rpH48
lNfDFCSnmZiUsBK9lrZtIHYubj3/hA70gPLU0txfvmirslNk2imhO+dIX3874oZbfD661HojO1wv
+yhw2E+KARRrjAii+9WPhbwADFnq3pw0gT1tE0PttFusHMgLV8qbiOH0I5tocxPPYFOYJ4yqa+61
2BMh1MP2yTd0XaclLYX+exi6lrWnxLvI04BsU0beMRM7aop/IOgN7Ijx+Lhe6UCplnbDxqXWqOVn
pXTgd0/2ylZS69AIyx1l/eZpdjg2GyOElfY5Yh6YOPB/d5Oyqq+NPNPXyBB0Poq+vnVC8F7GpeM0
WeFg5P5WT6mQPBCk/UxcH0IDVezcqeKKbcyySUkpWMVuv7Ah391wn1WPADXY7/sVK+h37CFru2kK
6xN1ZOVlbQZ1RcuHD65xCvkMVtejcb4+CjINY+LZcWi23ZeFRcRb//IY2yUiYLzv4KnH8ci+n8KW
OBYzxikNYG9wf6BMfVns4Ee/e2/PWKEpu4QMlBn4cgooGVits20q8P40dqEUYea3ukt+SePnuOgd
kC0FN5/A0DsOSlLzjId7gvop52BPR0vh0D2b0Cfg4suMP2XjGHO+FYWH3eHiW//zCivf0P48OLv0
2Ewg1Gategv3ybxlr4Pa436AiNgSnGn3JiaK63zFCaP6V0PxyaG/U1BEChmcC9dsBSjy5IcHOelP
Lj0aPQjNkQZSOCL78b+P1iKcUGdGXdVfGiQrX3eMd6Dm3GA6Ubqb9f9ruGGMtgJCBorKoqydH5Dx
W8F+vgJ7KoVjEhupVlSUMOg1HYqAJp9h90fOj3nWGeDMVOW/cnd/4+Nfkxq7/TL/427kTS7QIqFo
MoJhSvxtmq5ZmS0ZWOO2Do1h5//87FDs8MUmpySPQkeI6GN55p3exFvxOrK87tDsJfApy+jxBCfM
9fIZ0nslHKxSroFK8jX+w9xYjw32VeNAXnUnpH3lLIK8/WQzAO14oKG/BEW2rnvdPvmNW4qKbbmQ
fd9z5fzeZeISFVj3SipUE8XQIt/HkiS0UwJG4KhAawfQMbMz0f/Bw7v/rPD/5pkQ3Cu6FwR+wls8
rATO8i3TJxMr8j6yvND7IOIQPkmZbUOTlRzUZYSJZcYdcuMiFJhXKg/0ckbnOXoLb68SQJXAGb0D
39tC+ILty1JSFSqOxeZbD+Ou0IxUtQ1roc/lZMxva+rS+qt1rJ8KR03dN2/F31sdKtuj2XunS/op
7YVH9mHWMn3j8bZ3Lx08ak24M+EFqPTfUZfI5I0lfxYsiQ138AMtVq6oLYfHEqRuSmyjTiIsspDI
pI7h1lOO+oHvFs45dtMP3T3OA54RSPvIG3dJnOg1OLDlgqmHcxBJDY2rLNs31m9pcANBTPqNccUx
yVz8ZpnsZd3tDiPZqa9XiCn+8RUIBC4qTUxFTshBumyFagfv6Hz2TifeSwm9b6qrLGUUoYdumK0q
LfxF85GV1/IURZIv0u/8rrl6XGEMYgnrAsykGZH3oFMrkwbKqsWN+ck1JyTo/ncaYE3DNMjgev0K
ElK/SbgXMFYPTyT83h4Kh/1RBnknBRBOrbD1szdG7PM7Jx+Mh4hEzili/NZoO2WCsPIahMLxl/VQ
MrRfxQFgUuky8mEnUfpXFG45FlgVQmXs3+HCgffN1mGvDdOe2v65iozegTABE8rC9WK8q8xma5TZ
KLUsBnaTQQ6qg4YUvA0nHvhUWCNv+NZSxNXaMjWeYenKGiJmTkYNRb0IzUmwjm1kidq9BH/bc5b3
jNaRAOyfJA6ZGwz7Z+6epDswGAE657kx4RCIcjH0M3zqQuzQHonKFb9qZP89TKxya4PmQ2wIao4b
xoALdEcMZGZpdQobFYfwSgo8cgikA5xizzR2unBhs616tungB1Q5Z24QRdEIzyipAST5ORh01JCI
RJpgSWWgzPQ82Y3ltZMV9Lf+qt9WQj6r7erF4QvybzaWbBS7VzRgDYTj0UJVdhN6svKXMfMmiRFZ
EOMtIfGOsMmaHRf6bsmzY3puZnm4bcPXj2XvJulFgzVh6QcAxlURTejUZVKox3N1ZLhdmEuKVHnQ
t/0UqLIpgOBDLXiqhjOGuZqfQ4Jhi0PVcZSMvm6SJnPvHTJMvmbMIYgk1kyNelsSfVvbBAwQFBSi
bO+8Q5AR286mRPQwnzj3z27+mznTbiK97C2nzc8pSvuZy6OtP2KhgwSxIQqqqFw3q5gQrah8VfVR
b/9nF25TXbjd1J/f4vC0L0NXiYCEjEDVzTV22ymOulOGJGp3/ETomjNp0YAIERN1R6j+rX1hU2Sm
7lXg6GzyCzkCS56sSImct/5h1DuaIgeLRNXEMdSo/eFQa7HPjmPZovcWSnqLirkBISyMmLQVYV9y
xluXQwCSCKekcl7gSyGkOG9utwDvQsAogtA5iG3PnRge0i7zmirMf7aJHSvaXOXEtK2LxongOCCG
n0dYClpCUH+K1eA8l1IWHWGHMxaSPJO/kTZGfuMQXnRIVkvSV3COw/sv20MHdIdyBJl449IL1pQy
omxtiQUb2ygtWOYu8T3xbZr2xN/i7cEHiL1qlo8Dm65LniNbTbKjSqP+UuT8cmR8pPpYDx2H3k48
vZ6B2XkwHTnyNR7ihDBC8MXan1fyCJr0Ir9zN7SRVUes5pzsNupEaRzYMGa4VRk4wmfSF+QgubYu
dQjlKnbIsyPOQRcA2GHhiqXWqxOWTg6kNCufR969QtZAYhf7Vw5OXGLWLcooC9m52IrP4Ltys+ou
ghwee3j89dq8kZrskvb6ug/k7rH10ubl4G9+Mn+ydI2WU9yDThxbo00avJkSUbQ1xuV2QNOlRnms
zpV/bp2vRWx3bo1dMBYdoWArwki+VH0FS0tb2epCs7evYdKZGwSH/+IlGeNjlO6vxGZN6GmgI7+i
kKCsVcG8ck59+y89RstMu4esfXE9yUS6V/HwigMaI43gssFqPurg0tjwAsFieL+CItMsqvRFn9/A
1gW/NaYL7hEgbAoqNn9TOAS5EmGpp8Vb26q7auiBWBO2BBy9ePwPZQt02BS2kkDI4r6qiF44EpUp
UzgosRki2VyjjkPUxvRqPJjSLzKWmmUeA6v7WqiOSvFNggakyG0ra+b05ra9VQQrpBcVo/nDz5jx
7WPsWx9793WKibbs02im70TfSYvWa+IdG7Vl1lrBSus8xIh4YvCGi4OglWPufh6uJ1RiimkmmdwF
5P02B8VjNBjyjpBj/mJk13D53MCPXnWHgzb4PqZ9Cd8Z/7nexXlRsF7mI2YTAP6CmCyUA56JeL1w
LlMTj/DRQhwmSK6/NitGTZNwryQyOTnFXwE3P9wJzg4GFstrsmNKX62MF6ql35TdfSyFjwk7nk4x
HBQ8atsRoa1d4Gbp9f36foYd1Jf/7w5Ve9Tu34RvezefF6qvljfMvp5oIGrkQQCDej22hblOWKPK
cluTvCUfGksECDF30pY5fZ4PvIMJgbCoNnnG0FCxrWZJ23y8PXw53UiGhayKEMHJiMKTAqEi9QmV
NIYtCsfqu8cyVrVAJ+ake0nNV+Zj3hsRgI79E8I8KM/gHzD9FSZvzCwbkhG7O55PPcxABsPGKLVX
v96j67qsGKvZQm9aw4Rf/Uwq8xf2kkEGpRrNA/ZxXhcTwpvRPBwjZYyf+BBls3sBfyvbk45wrAlb
bH+fRawwK6LvCv4MHxticGOnUFgUahOKy3oWte2bLAaIFu+ftIlb0PTw3MiG3Xve7IGRObqhQW2R
3k/U/v3CDQiUEA7PNfzL9pNzFMR5Yarw7SckoHb2oOkKH58GMeas8GVgoFcEHdBuc81hsUPp9yz3
Su78AZ+zzaNT57pp16GMzdvBEhx6YEa3lTdENBnvOlcIaX9gB6qBLhW+ci/tc7ejAsGg7i2aj2Bd
L0wLXR1a9rRFNyosKJkw4ZDkilcDovxU259JtO7NSdKCHAeMczQkHlJ5JY+MjsFu6pLuT9j0T8sA
x4fHCB5r43StlNon2vcL8IqqGAvlkAbhR8WPywR8QdyPzxDogRm4BFi+HaDYNzF5iFQi+rhWYojy
sLA09cpyBjqyjOryeC1Zdz4zF/JLD2VlcBnqqH7jQOBP0GvaWtNiC5JcnIIzyY+pdPUvkq5x0KFo
KR1fo05foUD5ERFe/EWY/oaID6I4l9WUzKKAIwQo5XgrJQuuSbthmawJjsvsUvDk+1JXtIglliEE
a+MJ+knYsLUzsG5YNtUTa2YoUdDPNnnRtpyuQAQb1kAmgVWkMjoCTYUVqooqsW4xZkkgU+A1J/1V
NMQR1f2qYkXKSmfHFLzgTVdCPFXcjIcTZg2iKCfv1MOSaZH28ydiCck3OG+HNnM0o06kFLvUQOb4
B5r00RlWLB/sK8GMk9xMMslhfw5d2vM+gjNxOu4GLNOJj3vxHFyDbJJdfPgZ/DP1DI2tXM0un62L
VgghDrW9j2o/zN0NMmOPy+gTX7XlrWRbGwpEVZLxenbKTutcoHwAqcBeMwhxcvpE+Whbwy1SWi4I
yYzRAJtgLKJSQpoxl1P0FRQOUmnN8W0Y/Ak+FR1492BrG7Gd6o3qyNOV0bPuJ3FGk4aswS8YpBRW
Ycc7e9L1qZecXPB/d/MINCa1stqvgnFjNIySk2L0neMmxIGeTDC4nkv/Oj5jhVGb8D1DNxZk3cJ8
NWN2FiFIiXknMS5nZ9F4iDFI46JWvtSxYwul4AkKjFDWTbjiOQaBX2G2g7ww4OH4idkDloJbrvg3
Agfg7TP7kZyFFkFpInUEp9uYuBMkWllQblzmEDMXWBDgeO3L955zzdPrVeVKmja8zrwFmmXbdUvB
iey+XQ9gEZGXmPclqrWKrs9huEfN0dQxlFctC1zlGNT2fbImpZBeVrH7Og5ypMAc0czl0k8dEbMG
CulM5ja5TC9AVgn+vNFp1izdSA7Rc/GAc7kQaynp8LzOkHCxT9nCfNbmZSnYiJVgiKlrV7ExcmZU
vzuQopoomRiorYKiweL+IQe3fEpeuXw1e+yBjEdaMI4yx4x1TdpGm8gkpEOSdO5j5gwQLVjexoId
LU0GXdra6jC5IIdz46nk0JUyr4lTnjxFcwDzfL9ztSU78DCj1Tei/jBfJBjNPqN7f5zYeK4TyFqx
yCN1MmqrKCVMPfterH4tyUtQ7NaBTfHtu2HMhe6GRsGpEK+bTceFxa6hGEm4wEcL9E16j7s4YfcP
I35cke0DV2DDlILBp+eNTRoZkKCvXetuUudIilJ7nrKbghtfbDb1w3VdbxcW7MlG/2mMvCZsue/I
k03XENQK0kSAScWWcvjJkvuacKeWcjl/pz2wpt4osStw2f+mdudOrFDXYQOLeIFHoNOkBze+TaFZ
ZW+jih0nM9bonerVY9qMPVzSPK0OEdTRy9NtsUJQdn+ZFhJSeuE5G69xmt8UVMrkFw2sBlXLKyvb
fBYWO39P0HQEVgd23WVUhjd9oorvZmz/8SzLHR4EO0rSGSMyG9IjMhm7bhc7GBtLF/Lw5TA5tp5S
TycLAWUcRUR66GFMhZwxOwUQ6Q7RybND0S8DrxDBi8grS3K9TlAI5c10I6WGY1NVY+BE82TIuKd2
p6Ezyckv2WWrD7PM/VLIWXrUuhIF23VqwGP0fdyApgh84tRUqA6NyhaC1PnjJoaw9xxBR+VWY/Us
RHAQ2nkB8UWk9IRpSuf4s1qdO1qKVqxAaMl8NS9YaP0LUG8cz3k+QLJ0J3dYF/DGbB/KDMnpYICi
kJJiQPMsRlKN6YZy1idK8qSMbI43YzSioqbY63tVPU7MvNb7xDhI1TTOam47IorSwVe7QltPYNjo
3n62So1gCJ5tEZJoiyU2SGY8O6NlGeAc3qKrWK+hJcYkECL/fVQ4EGW/dSbocwn7ITKiqFOPdOM2
+Fhs0RlJdizz104BrjlQRMWeb+8qxfjO33bXFcxWDpfUuSdM++CrHYP3lTDGAgpmt85tBqBJHMIn
TnC7CMz6cQXSitqZxGadi0n+vCmJFcCEjjrZHYUxKcPQkKZ5wC+JKylbv7r0O6HFOVXI77jxnnAk
mxtTQQa32B+AVXoAVd4UiLyzeT8hwWNcxQL/LEX8J2rAhJmR8ZVlGjai7SJvhnMNgqH3vu8Li3vr
niAeSLVl/Aqgz9hZT9vobtk/1Km6LPRrxgdPrmL90UdbmasU8SCri+SDEl5Y1VQGJl/lJj6cai4j
Ry96WEFQgug5v36qGfs4VkU3wF/Y8nRRnsqfQp5mmiV/ZgfSJdq83+f8/oDX/F/b2ntlcCVfQoA8
I/mrY1qOhOsfr527Q8Sch+cERO3Zt+6cO9Qvu6cO15KQxWa59s/OMm/u+J3PbyV9aq3gyYxzIk3j
944oQaArhOYx9i5HyCaM/z5VT2VIPg4EMObWDCeSrQro848mwnUaUdTP7TFPqA6zB0NmvFyabX7C
bCBaLBq4w5cQKAV5FIVJXz9D1dMrgq7Ex5WO/jC+F5jP8Al0nHb7P3hHN7x8+XRm2bA57Y8evtpC
GDtDLbcUeTajQb2ylhbXGb6cEVDKmTc2lJi0p1Kda0uWKX78+ZrxUdk1r1oyARTEnpUfZ0w6BDth
8ij6MPzmhquFOBWRac7ZXkKylhMArtHobQ+hmm6OPBEiVOHd4S7hXvAsEYNFMHVVmML9PO8ODrQQ
E1AppY8GL6Ed8AwIMJtUfLD2Ex4n1PWWtukg0TFTfpNTia7bfwujt9XTodI3O85uae96PfNxcKnF
JZWsLtNpB5pMQxpWlEast1dQyF4teXb3gXBNm7yX9sbd4i0wys1fBITcR1aQnhiAzVH34odrpWih
y48XIyjW99ZQ2rimDZCsyoqWF5WnyjMrmLLBbOu0k+yzYyskVHy23UtmgMPTjlLPj6P1PNJoTQtf
ujkbzcokzqpldzTezDLvF96vtIMBKbejuSpDWYalXbdM0+ussRO/ZjcaNV/KQDxHHwmc44yR6Ilx
VwGWrRx8c4gsp0NKKu8ypAkULwGWyBanLgkzgYVku2dj16Q1DZ5cyhzgqaiVuW90GIj/wVsoAKqv
4cChR4mT6Vbh1wkAZXoBc0SOgUNf8QB765g2LRKiMUbPb6uup9xEK4I4XSBToOh0QPnO1yWbVyNa
at4xJSkwMp/hGnelJA6POMmQ/jHBsPzlr2t96ql8jq/lz10b7EIbbvgnl1NvVWMCwPw66YruYagy
p+O3auotiKGOYRhJLeu4zc3VfKARfFhMnS5kMjPgEKeAX9Cu4tvJ/oL8RmLihpuajjqMRa+mApBi
XxHG8rYUOs3rOBA0NFUM7V2QdRudQygtdMN0QyCMT7OkMAIrVcOg/fa4Ho2me1xPXJjMX1I1s575
xO57uCZvdZEJHevUS50jYP9FBsUqeEioTRc9U6mISn0o3cF7EUdlUJPEMBK40mJad0XjCKq8Ys40
xkG4LF68NvwsJi+t++8khPf0wEYjydbfyPAO8Qdr38PFUfjQzEraToTlJbisu1fgRzy+ge/Kag0U
ZhCmZrw6aqoBlylBUu1TdR8777KZW5lKubxCtL4247P67xtXVBMM+0wQx4H4oYK3/eWslzM5Hyij
pjPT5ot3Oj4WUcsuzrrB6NYIpKK2aPCRXTwP0V5+fIpQq61hwsN6Otgco80dMTJTyqB47HP+6Uy+
VoOGuRgdYuMQhY4+OGQTQ/D2Ok9YFHakzxEC06HFKROwL9y7SgureIPPdT7dEueAwWg/WOdfctBR
eNmf/JhaEuH0k3jn1NtSY21t6QB5CqssMVy8oiM8rMYnHGEmGuJ/qby05+Acgt1OIDX9yV1AEp16
dzr6fUKFBbOQnkSSTU6KlYXGxxYoKywGCI0SDdyR4O8l4HJ2ekVH37F+f5W+iHGQXNE13sv6V1db
BCgucOKZ4pWVuPnVVc5uCCHV4jHV4GCs1/4+j1D0TpTFN4ZW6sQh2jmL8i0QOVf+Jbw8/W3g+yMM
bFmHdlAQieHIYBu0ThY6Toavr35z5/ZkM5nHRFw3Ulw3u7uLeap2CIRRyo/4MhWr7E5GOTTwIdLD
eTsY9DDTyKxl3DHM8LOWw8QTD86vQsJnfOnOhBuCM0JAbpDJPQNLYrhv8ClKyTq+mh3SKVnQyhPw
aWQ50S9/zw+Vdoqz3q/DmoQ+WNkHghnKOgDupM2sbqBVcEJzC0mzwwuodMxJNrgGiZOv+uUyXpFB
zILap7mqq74VIQq8RUqwLfkByiz0uFUoxoD/AxjJk4Bz74IaB3qQ9O4Mo9BC4C1LbeC4K2cY8KI5
mDXmCppnXauThyKCq8DwN8yaJjsmy+lefimAw/X56Po8USXTxGv/T5fb9wg8/Ujat4tCJajMoYvb
PgxmVBClUtWvMr/h60+92+wJaS3czjNpMFSsElktG5x5ixKooOOtLJ13y9B9lFhoehgOyOCL064j
BSPGBvTvLqC3mtgWL3AzRT+UBr0yrCCcVmmrPO1V0YaFmJODOXeU5YHVvY2cKgdKiZtCQ7Ap88bK
7yIFx1P90YiJedQeop/cGvYQKyy9I7mCWIthRTAmGLw52tIHwiTu1WbVqairaI15SGslt5I3jM2z
+vMHi96VQfdT+ixI9bW1bV0Mu31tIyGkq5kivpk3fLCMrzt+rUGvfGMEVV+k6k6JiYy5GimPx62t
cBcKJHrTfBF14+CGXEMFG1oRP01VZyRu6CgK3jtPPEkldN9SHXWmWE4iqv8Y1gCDkfCNx7BZbQo/
XFFi2KTkUgXekPLrikDY5GCxZMr3Z81Rx4LB6AlWrklxIJ3lrSRw2uNVPQmn2G85xgo5COL25KyP
Bdlijsh0UH+xN58+me45oNKFuiq2tAQZ/fcTMSs+j3Oh6kpCsnyMgOKzLuH3GHomRjhCxNTfw8yd
15Cxj4NcbnO/F/+d9jdmhZzhzbvlde99EAmct+M95ToAVakzo6n3/1DIBBgAN+9/ZQEXMEHACc3D
BpWJt22HN0vTObSpwPxVf6UEUsIfJvf7cNfQ9dtPzBLwe+HhUikKb55p2i5eSprQY0lF3rtSHyAl
oyXn6n2E7SlumZnkh67YuEXaC5T36hH2SbQZNmX2tt94hbyj/U4NZMzxf00X3rBc4bcASywCb3Lf
lD+9if9NwXA7ND2StpV5Vv9xYzyYGCK+FfeHIjtfXgZsz6MVHPm2/oO3NgzFE+vhZHM9UeYQNd16
jwi9ppIuQzFAmcvJknmaQOc8dZKu+grpv8HthOChKYT8ez/t6NFRmsJIgtvZgWk0P21u9WMxdo/D
vtjN+4dST86fCoAT4CfKv8RwGJXWc9lrxWGmbmLUq2S4AgiczxaxKd7e4icXB2A3Z5YoNYEtt+nz
H6mh3Z478xszS9Jx+Hatrzde1+BjjzajOPs/xbkVy34CZTm7xNpxl2XO8HfxITa2tX1KytxRj5q/
0Fi14TL2o4mn24+BOpDEPISjE/74+260OU11W/r/rTEIMRmj47R5gE8sE9QaFZErhvjhODMMuTox
wmHNmMT9kSt8gNnfQcauzSL63P++HhIDkZv2e07eaMX4B6aaOjSBBWYK2zgDbmTFaYswOPth7QV/
x+YBDlKUS2QMO3KS99jgJFfNVxX4ktMm+yM9ORZuRnGBPRtp9LJ5jSH9TYBiUd7jLrJBdFjgfnFa
oP/8dKjT38JftSmw7RvQf21l7JdO0+h3yUQUKmdOrMpKs4SgO332kWxiZbr7G4HaAPYH/LYyvFty
hFTloUOnHwd4rQ3EY9oP4DlvPuqCdrSV4ScsjTi7PcYvKRTWjQPzsz8pPJN1NFQj04fB0zB4VnGp
pglNHW+KQ0oNQ40JYtrgwh3imIgGwS34KbfO+VONZbf1DVNbHRgOMv1RmPIBUONiqOvrx6dQ/O67
8Qm9fFmNXd4QuT5+JZbsKWLTS9ljL/YOOr4nVL28iRSieTIsLL5JK2HjsUPDR6+qObD4BKHKBBzm
U3dMYCUO6PXxFyluPfSRQxGXNj2h0OKlPAYZWf5Nbe//QhGZHZ6X1O1NMWuT9htSM1JaMDgg0uNQ
VAZjK8pnBPJt98l+0C7BenOJjj1JWTSeY0abZxTZuVvVunyLQMWuA3OT4DxqYPyCrhsFx2LpLJK7
dcMiVQM5Nxo2lTlRKS29fhJtab+vCEnJ9DoEP8qa+OsFjCctGLOc30fTGtAxOBWH6tyPZNUhuYzF
qKTkIzGEQp/qagnrCsASCrqdf5Z5nNG7fGl7Z6rFrx3oxVnh3MwTtvnyjnJZNg8UeUGsmptH9p3a
RPc79ZVKd0AQ1NplERM7jIrSZef8OGh/GXhi4gGkeL3+mVXcktbI1tmMXl5QPcCv7bHHUiUEw+qa
1CzoHltLNTIMPco9gzNbFaz+JHk/uU+6IA/jnSdG5hdLsNNbS3zged0mZeQoOpi0rNz/XOX7ASvo
Qfg6LF6rwrpCMLXQTNW2iM9LBm0CxNC5xX6ZavjagPd+lIc1jdbvwqw6razBzhD2uVPQXbAWUhtz
+XxVOXYAFPayzscSdHXHrb3f2prLCN3WTffv+9Egyo2ichucEznGqEqFByJnE671x/qA3l/l5kak
0eoypCiHm/pQk9I6QOgS8PwWC2FtjN3Gr66qsBococNB8ilWRBk7ic9gypG2oyz2Ewy/DNjZ/SZA
o8ycxfQX5HT0mSDClkvZpkNgVAfCJii8/3K1Sk4n+DoSqfE6YQcMMbEp2t5xohQwm6gz5LJVdRf0
DaBc7gTTiBr7dSvbhCMc3wQZnfBFfOHxTime0OARPO4d51GMTqUJF6yDNTni5yZFnocqsS9Id9DM
GhsnxmJat3gLXJsbnemqfF3DIaF7RwTLT4yXtItwcq9iKT4UktYnArDKhVK5BJbOWsclKxZrEDKo
wafOQslqyUZEgsKh30araWSLPh14JysI2V/o7LIJoTvmnRRycgSaNvS2R3sr1WT4hr7XgbLEJXKL
R6rl69dlG79lmghY2Zxk075nGAEyY+WV8ijDm+QkFO1whSBLmyZWFFpQuc+8oHws6Hk7JRaDv0y6
+buDiDUTx9sBWcPGEnqHoVo1lzG4/90mBuzcq9EoVy5Z6UerCY5KjgkZsH43nBgUFzGwOgtRAyQN
iCdTb311JwftHayjZBJccRdnbndLEX0b6CypY1WmW1RV03uE6ggQZvCaxhXyRvxotGQzllAxZVfZ
e060JDuWVimkIo0jv2z2Pa2p4lDAfU7nI7RwkNaA4qsq6+vYuGfsBRf995OWB3BYQO1r86cNBqeo
xVsREttsL8CjbaI77Zs2CnORMH0Og8TLC2xp6FIKTkbkJ0bRyQ2cAx2JrzRHArwuFMqixOqxf4s7
WJ30rJDrwubtRQBPvCFFcNTlwbvgjGRQyE/J9auqqjZOT0VMVUZSCaPgha3jWYtbB3Ygy5Ni1byG
u03BfFv1FlGee1uozqcCczucNec4O5C1Nx5FLs2KZQKAxphCbAdx+zo4GmmjlwJ8jDQCWL/hwWUG
BUv8017mCN7g2qZpVbizYU8OpCoagXHzkh0f7fOq40Og0T61lDctEQrdeGH30RWWSQGjWXl6tkfH
fZO2RS9ObBR3e0dL24g3ZLVlSA6hy3Fdtm8ll+QImEluGEwJ8utT9Ph27COKWuithN0UX4XaPpZx
aCOEsxJ6RPNZXCHR5Xt5yoqc5fIFQoxBLRWdtCpoV+/xa03GVp/aGUXT9cC5P5+DKpk6pvY6ysmX
TXAzCYbHRLNd9qxvK6rAzMo5Qn/5qqp3R2YH+dggnmGpnop7nNTZqJ/5pNxnQKijE/IGunaC0esh
MM7tvQ9dZ2iRvpOZWB4MVRUm+HpGH2Ci7FeOzEKS97t+MM0SDMF37TVAM+G43y1BHEVMH/UOIB8P
Tt7UunQdTWEuZfksIS+l7IiEssTVqs4USCkX9FDsvv9ItPJpUk+wkda3Q/XUoGD0bd9VKGrIPV9Y
SCz8rzK9dOKOZbZ4nl9j8ZJqvzsY0MWSbT17GhYyFhIZSN1yTVOaLgwKDFeoNBptpP7nTGAvnK8l
rTgixZUKuglmEhvKRbuZYjcCNpPIe/Wv8jneZAIV3YRQnTgflQAteJuQWr1MMkk+74TZi9IJOz05
qUtUJMjadvEYmb2JpLhgfTHsLsl4evUxjlWdgVOvvqeKrQZS+A6G/NHvQtEONmzugLgemRzMDboJ
NSZ5KtB1xTCXQdZzGVGWf8SqH09fH/xSojeq0nPoki++i9kf10UQshGJ60wJgxWABBJk+NxZ1HbI
P8K8ZtWF9Qvqtewilro/BBrVrJ37PhhcwaHOyQQ1G158w6xua8xD9hxTAJ2fIBEBh38NsgqweXXe
ITyDGONyUL9Vj9hKjGwBUEwFQ5nKTyysFbp4JvI68O4CmmTN393gsqW+Z0gTqrNBSlE6F6uuM8Kq
jVSvvybVD58aDk4CeiAedYvbEzwv2cXRDVq2yTInmjzP1/zLITD6A2lHC06yCFCBtjfrrLweWOX2
Ze1qhkHRJUQDbRP4ahRaCqIvxqHTqTbbev3xcfaE13+OgPM6AUTSdYwjRHdf414kaF0KvPFaLu7G
UiDjRHMxzw/EWZHqG0R+1tkSRQNOQ4bQZI+W9jBXcMml//bMVhi2f/jLm6egAGyGIIGZZZte5UlT
RFQFC8pm3ExgGJoFCwFm5XA+y/GuYQfxV7RB0WYJJDOqvxTbhTi98jUOtTeXfmesLVven+fvIT6m
o8moOkRn18AsCtbUFuduRKdtOzMETmvbAjYzX0dMytIkTGdpLGaKKbCYNGFXjt9iW39a/Oshkz8i
4EsRRm8eonkSuQOfZ2OdkYDiTtXgFn8C6Riuu858RWwbZpTk7zhift6BKBbDpqbVBrgM3GbYDfJO
RhAsaHlf90BXTXuwHyH4qyh0bLEFTI+uKTzVKJuj6Y4UKB3b3U8Wl7Apn6vnQDvIG5pamHTWzmPO
RGfdVBxGtzDlIep9zMKjajJqKSroadCNDa6w7eYa2xI5ZwXtNbeBf5h7zv25pFlNCttJuk8p0XtE
ObHOYxmaC+4d4tLBYM4Q52FpTqSikA2cPWFcVget0Osu6I2GVUfqogpx5uutE3ptsnuaGB9f/zK3
xBveHCwY0jMtJwlegdZuSLLLg+LwtZ3RGCtmHJGBd5/+fvLhl5QAVKuanzhV7+tEx34sZTgy3i6X
15Sxlo2QzifknaqiS+cUp7SY1P1a/o/yG0u/nG9Zp06ssa8OfICePwhcq3uvPSHPI4aykOioya8E
j03dseULq0++pHgKJfiBE9VQFoGebbRAvLowuKEkYVNBmrCMmiHTai8COP3Tn+k6HYI/6/WTKqrA
wtkr7D2GMZ46z3Y+EvMtsaVDVggSH+QjCqcF1pwmtPh4QMeCJdh6Fvbq7ArEMWpGjZM5+JkzHnTA
uNVlVFpnt5DeevbSI8bwPwU9jk1ZpVqSncUIoWfcsUxL2KpZkZOiCiiETG9G4YnbYdLbcbGDMChr
BIJXTxzWoG/4ET0gW1M5WspdUw5Zmf0PkTfI5Js0KUjhM6KWjC9bAt6hydz41lp8ztigNqu8SEO2
lpLiPBeqJP3+EtI/W63qDB+hUporm9Gt77ZumPLZTG7liguewYw8rmhcoQvWJBMbAd+DGlAQtZxZ
7E872F7NwsC6YcmUAwUbCwYUwaKF7cD1VHWqxyhQNsTTWMudm3CP6Lsqqmp/wBOa9dtqySVYA35+
nrV0wm9kN9hXZKOUfR7U427zitmhA5bqHkUfOm22BJaYgf/FQRvQHkwELxh4H1ccBtf0GL6+gVj7
rv8ASJ7A/UG3h2sgAhLO2/YISbHBSQR1Ncxp/F4bq3LAstsAV6GX3vLpUXWVwqjCs0vklb0JffuX
sfV05Ejtv7u2wYPfZLVCw+IHaUHQgH830R+PWHSRfhBsWKfyZV/DnDQYWgDeksaImPPDkzsjdrQo
VGTeJcmMz2p/s9Q79r3wnw+DNm/2f3nqSvqIpjQ03xblAQIJWPnocxzzNQ88hDwY+gfjFBYDDaXk
4z1GFfE+DlnqYKPyHbzP9OcSNWAj9NAkiPdU4f5pCcWRFPt+zYvUx5YM4p1DZVgyib9yNNN2uWww
86yCh3J3Gs88aCE86h+hEJJ//QihxTTjeV1S4ykxsgUpt/0YYxAzYg63ZjWWirEpe41TriefoCEP
0OCgPgm7en9uubrRdPwNy83/KSAONSZuz1plq8Vr6IpHGqDUlVyieYZPAUofnSTH9xA5CxTzLHI8
RtvQDoRGp6WKzjQg4pVvPnB5TU2tDOLI8hPkjOfhrgcZqM7yy37N75EWoUw7GKz1alPtcxHIHYfS
GX1Gk1UmWD+OrgQXJMOuhSC+1O84IlKILhA2zYzU0GwV+OsVgDHWgYfPZkI8AKtNwzE39mB/dcwf
qFqYxtT6ALfEmFtq0GNeWPRlrDk6TU6d2OtLZbWqpA2puU1Tl1S+/q66N4vA8iWP4ldjkLkyUp79
3V8Gn+P25EmRyCGoyPHbK/adQaeEO/l8s0B5ORUV9EZD9ChZKc8qg0/rp9DRTd7NvK8Gz8sBipHR
aUHRu66f3GjLjVPifb+kG6P3x7LfE5KYv4TWtEpsdNtTG5lJ5huTj+CZiXN9TSa/lmYA3051LBZh
VB/ytKgSOkAbGcIXIRdDiqMR5yOVkMftup6QWJSbRLC29y93nMZtq8/LP4sGNJl1U9dvvdNC3ubg
TyqLFaOlT3UfTrI/9OrZADfVM8hIKGzgovseOgS+140687k05igPwNx9DUuh3esCmOy8Hfy6PSHZ
iGyteKK5QSd4iBnkAsnGeAOeK6Vvgu4d8Q0GJbLoPIEsrsrdT2NKsC8TiYv00uis0cRCTsl2paW1
H9ie5KAUJ6igByPXQD3UdAMegfHhjnktIoxj9z7nk/iZQwlnUI6KONqtCdaQmeehf40T+AEIhP8m
22+pMaoTzgTJHeZVTubw08+/rvoAOy0TrU51E47XNAB4n2mGd81+1lwtS0lhQwWr3Zfa1BAnItJk
RZaA4Ufnh4xLfgn0qqivxWf+rVCJJc1n3wZ+An2966hOU4Vd78Wf+pYcJEaOf9J0GXMbESUCA3Wj
BFi/KflR2K8Hp+sdyD3mz+/amLbD9soHHPHchXRMK9xRE1Z5mrH+rKG44OxWyj37zqkA3WmaEO5R
dCxpf0qlEyUsqoaV1X5gR1DUPeiUwM1umcZKLhsFKxbJ7+iaJFWDGi0IgKmfduGiAyunc139Xjqp
vyXYefdWfrK150nw67LrU7Jq9gFn1YV/nzrdLHG4Z3bCD5bGkfn0CDI5rDnhr2BWbgPIQ1dev1GI
9+MGuXX/aMetUHOAS4ry2wzGSyki5IgvgsfkuK7XDaZLVWG9eiGnzm6KOTKga0dB0z356x5RHb0l
Kv1YCenjO9f7SnYlWT4MlGFky4DutotF3TFleiPv9ANjt3YpzZFHYoqf7LC27l1QMmA8t9KhP3ZN
kqYGUiME/WmW1p+XQPkMBZ3t9y+v+eF5phjOrqiHhZnNG52Gxr1DNaS7/GJUxG+oRRN3d144h82a
jK580CkV+E6s5u/FxbwuLzyVTPgquzAB+E0esZxZZtQIpASs4+v4r6VygWAymfXHWzg9xtYPJKmP
oG49tMylhVt6NF2hW+i0IAWkG1+C0w4VcZF3903sstlP8DUmDz9SD9LiCYkVWNpJ5aXKztxM2dQD
5X7S6fwEg6/xrt9+PRuNCRrAvhXTgFQ8qrdJhUdmOOud/kxw+28LwmAlPOFnJ5zqh18NL+hbTfRP
cdSKjR49LV2WlZAMJ5V0wbPFa+uC215jgMfj+ZyVpfxrRDI1Q3t9c9gi2qTRH8nPFkOtdDelUmpy
qu11/fZvYjYfPy70QBgP3Af78l6wfH52s8DXfVyVjGI5AMBeTxNorGDr+fsy4gE0/+qWRO+LHVoW
f8F3CVJDKQKIdwdUrU78SgHRSk2c/GbfNKnB6uz+YGCX2zYxulEXQix3j3U9ca8+7GorCBMivt9j
vZPLhU8z9asC1pA2DeLbQjVnhLGj7ocYMTLxk144XYUZduTxCqZRpM5qSGQSqTS7PGDXtNR1qZ9a
XWd39i/HAI3iPhTdZaURGRAJxxIuu37ZG6ZcijJg/3C6RD5SLsvmlXqIEjOG6w0eLQ9UJ42438Gm
Sq8OBMnlFRXurn7PhGAb5dNf5XxT8IkbzVW9iXy0xBhskdimUhNifCTYGekyF62iojf1jKJnkmz2
0q7TEYaGyr9UoIX3o8PFq1tDxvsefijZdpDqxI4DDbkwMP1sc0lE7BOnikkW2nfkzJueYWFJTKma
piXxA8djrFNpB947XSH3mNqk134pNbe2KJLUu9cAC2pAsdHTYwaaehQ3PYbWiXFJ8BnO309Sn5YJ
H2q7TUX/DTCRQj0gKjWfKP58TntgZZUw1xsPGzxcybCjTHeeDIt1HgkFw3SmQ3UrTD3pAdS+rY5E
kFtdwweAZqduo4uvj5iY6f1RXFca7aEpw01QTCHtlhtF/chEzCSBd83Zdn1CvCv3qeieptK6P8wy
5/6p8N4NMxDC/ui3FUlUgrxDqIGUXm2K4p3pSOxK0vxHI9rmOToxPTe2bvaBugo6LojIWmLF/JkY
+KYoAkANED8bAhm9rRcuNcdcFi8sCpovJ60IwnVQ9Ie88uJX6ZZ2OBPetdVqjcFY4wSp8n+vNM13
0dN+qd5QHupv2P5sq2uNRgIZJ41KEks4ftpF8WfJtpx5ui4YKWiaW27PJA67c/dIWQWal2KieX6D
utIvi0U56NKu22vSd3FqX/iPpZNKe8q1R4qf1itswBO1TC9H9X4329OAfAPHWkmefEgBXAkFAX6K
3AFNeSMDWDjCpopdEsEyGrFMcxbZjxS6WobNxKLg5yRtylMStX5voMwjmrnQ4168i+LLg+ovV5lG
KePl5tpzmzbCUZWcQX8TzQt4PXKncj+xQo+kjgd9hunpTl4+uhu/23q/++BZ8DF2jpyueWeA5aiS
ula/h+7QzFubAequLjp+1SokT7cgd/H6PGRh++5NTn7MvguWKfoqFAIc6q5tjgMF4z4t21tyi2j8
kpAX1IkUYYhfg5Vf5QxOE8jdy5JrRdiVO+NiwJtxA8VTmw0AOW5VMF1wVOsUGqXIAb0tq+PVLcrl
5Z/uev0wqGqZ4YnUQTyY+/xRw9SyvEdN/IWd7sijcJafxFf7fOe7nmKfQ3tINmytzzRTcRm70GY5
vKE2a6Qjyu1hhqXmfqg/Rcb6e0gbdF2GOJos4wYP3//puL2rf/olPuYVfXZddcHYZVaSc7IzFLQC
If3zXJDI4xIRGLayKUuLkGRyq5Kr9VfgkzsBUH2QmbXvkVZ7It7X3XcXMwOpDTz+62Ze7pugP37G
tswPsmocx87CpwyPNzhOBs5JVv+jKDp2+VqaYxaikwoEqNRXB6I2/JgJw862svYUSV1YCnvyzr0b
luqYI/Fy/NuYqAM84E2cxBoCi3/bd7bP5Wr1iTgXNf6YdeDW6y8PvcOALBHBRa0ILa5t8XkaRkeO
6q3u2aahvkWKTP+CeFsEhebqgLibSXj4/KB8jXpCij4jYwxFfKf9/yT5H8phVBpU3AEohsrzUmls
eUFzKXRE2qTELyI3tEAYZM99j8AT2O054emoaHgUKKdcih6pY4YcBi0es6OqMv3nCC3WHcHNu+RR
eQ1E41SaweMP4PndY+4V+C1Z+nlYVYySisAeiXWRMZc2nGXDXMn6+qTu+v0h0CcohX36kcEkAVC9
0xqgKvnVAEqnD16PM92HOosIUCKZuPl+lj/rIaMWZ9rnmHCZfjeoIoSXi54vGwg1bD3elmvSzYyi
CyLmtDs8S/B6v1riyB+Ykk5taJ9evEYDNyepcOQkwJwlDXfz6OKqrZW7GtwPkf/iXiYxg3nwvA2t
ZyA6Ld+rbzMlfZSIhQQ+OZnmzmTIT17LL/yDvMZhG3lxLp8ewlB07KwgebgbrCu4kM0sIei9szmO
nJPvBwzJtm5QYXZBNe9yBCyB7tkE45WT59tZAhnU4fjstoT4zHMvtDo2WVgZjZ96u/S6N/wfa5HK
2eSrUGB4wpsdsC/w7m4BdxOxdTvsyrTjpY3tPZPTHpT6Iop+FOH1mcJLonSQBmjlb+4Zd6ECe32l
Dt6mSPiySfgkPcoVWwNLopzbP/zZ+EjPy17dJcWN3FJ3cOZGfi3P9Z2R2iqZEnkrfY4tkRYRQPFi
HCAbpcJiXwxND+gsY7rCySLeSVlH9vKIRgie60bwwKDg6DY9bWNGKtloy5VCqHLhjXVqYcr5nm5k
jO05HNTts0n/mtg6fp20MKhLOLI8+1jDY7vFK+tyuF/KNqINnScOGJlqTxh4A8p2kAfoGPHLW503
YzKm5DaIRsZFh2YLfsUSAdc+wjJEfw0j2TNWp/iWPjdGolodNFNCCg9PuPQ+RDDS562labdUV+5t
jsWsYj9axxAIOQJmSFxuA0FuUMjJRigOpqlJEKTSYxelCX9rTf05AhmvrMkXoi6QVcdL1WIYfC5v
u7ZC+XILK4h6D5dg/gK/bPZLLqyoeQCRiHaTPtfb2T/hYWKyUyoPPfBgcI3TT+ADOx6XuQeCEu80
IAgfON0loH550+pCHqmtP2+dcpI7lArULZUAtkSZ0SoVD9EWNqPtb0M6wNFQLjT9ANErE3Ipq79K
u22N8wag8rdsiPqzQfHcTvXwRUt9J2ZJ0FWrA1FsqNw+YQD+em7XMwbDXKwx2JzZDJtjSEO7hy2+
1Vg/PM2q8IBkZk5y3ypwrE3hCTyM7SvORCkwVBMC9+Qwg8gK0lVqM3asOvN9lODPbnUxhQmUbeS5
WxYJUPwlw6sRlqvwB7impZJvw9fKLC9jIGLsHpcxTgInsOpKhJza65lpl0dR27HwwjfwBSNxH7Rh
TsqQsHMivYobjuddo0ojGPAdHDEPATWuPbUEVI9rGs7mwUe5AqSME1mgcx6V0BYasfUzo7LI1ySB
CcoPvF4QA2cn4bCKZhc3s29MuiwnZYagVtPsWeX8Zlm/npYLtQSLNO2xjg47ER53Rn/aekWecg9K
y4ZESNAsRmlgwo6Ot3wy98/b9l+64cGtmrkLAjXxGPloMmjfyTahWCdpjR2j90i/18R1F/5hW9Ho
q+ERk/6gwOTodQxxWjHfRPRP4602TcMzXD3llx7VjBAWpOuFZuxgIbfFsawzmPnJoKqmSOFVoG91
fdKt+ny0GDyI0a0bPEqFF5IslO0Nb1Sc3bDfxZl3CNh2DZ1NWOLjjxk/dGQsEUNz6sRvdWMq7duH
Klq5M9l6vRRRlerl7IFawGTeq1dVs4IZJViprhb4QDd8kEKrEPlHx+8KGThOJsuMWyWiJzLk7uK8
X2xmDw5nIL8s2jsIdjs8uV8TKP3+L99SygrvX/U2r93VnP0OhT2l5joBFM/fDAmO8M/gmbrK3N3D
eCoqT+5vhYfBalMCOrzeugy2PUPWnZLqKaXJBT/hQLBrmecLy6srbnVprcfHFm+lA59tyd3ID9Gp
miINU7vCoTg4ZJt4iALYS7VJchAo6aNkz7jxwjR/PdIL442QOzeQMDo6whONCTMyYQ2TD3sZmMlC
SuTDXMOgsDdSBDmLbxwOQ3jtFmrlWCTPASTcWL3TI1cm1jcx0wCqrAx2xu9be0CKtrSbKr1ahiR1
RxycAjLU7srHd2FWlXAXEFHxNReElhEgFwX7dVReTqSmizvgrpLjg5pU6JB3J+4BThNXULBC0ouT
JLvn4/G3aFADFwbwZNdTAgbdKbuON1hFuDOjufiV/qW6Y3Q2WSewuyzZgE1IbGh7/7MMj1CsEDte
cOe32Lw4OZ8r2B7dG6RJKkQ9DbTZBTsP7UC0qHEX+tVu65ZXNtqFTzZ4V7448RTP4AtdatYO4TtM
EeXgJ2WRy9ctYq1Tr3G29h6fZcdbaBaXrWJ+BRhAJDyfEPyGGPLKlaVcaE2YgUuuf0oZaVHLYDPB
JNuyhb9TMa6NZIVJ01Krq1wo5eMBH+nvGATR7BeTNJumQkE/AlLMcScYk0jqR0P33iwaPqOM1gu0
CuZkfX1kGr6KWch4JIcssPkenfiOf2K6sydtLrkn3UDbzJsKdIp/zgLnkqwxALK4T+XgyLqxzHb6
Bt37A3t31gD30C0wrsUOXQ3i96RCwlGlUWgRxmgiBoDeOKg63cNjhoY5rQCmtUoQmxAjxx+1P8qd
8b1M6651qQRcBSdi4yvIY3qRS0572FxqmNveDg0olzUd/ImRZL94GzzlQqdZIAkSnOWlHtXXiGZR
KIv9IwOk8A6o12XaRoQKahg6/zIUJPm/jvOWwjF7/RT7VpHOPvuAU0C6SIEPUwY2WLJBNhee5KlK
31IyvwZg3fLmDk1DGytE5U4o3l5TRZFC2WeuNv5iyrRKTln/6y4z38gldAR8lnKuxNa53iFV6XZu
MZOaQqvmf6QqRSrlHPSOlp7Clx6J+93y3rc95/eoqPsIjJQHGXieBFSbJhcqa2ypycbaipih0ZTn
Mg5eWDl8PxwxakSqvUAwcHSWcGRqDc+8Clthkl47DYqNfkSZRd8xki8NxO8Cy9hqG5HEsedpL4Pb
VE5+F0cyTIeEUv9ynAaCPuKuNIREA0iNg1QsCia68m0FTzW3jwjv1DkuIT02Fj7Xa8w1pJxuA2wK
8Hu3BcLgeL9y/zojNYBG0nRpCIVOAW11fr6C7yNysqGfEMd8TJ8auFgmOBNWQkJ7tMP34WmurpBs
Qe+xxdVNRiytcNfKPLhMqPYqX3DxxxuW6BMnDwwFiRhHkJAavewLBUQOPwhu5Ss72gDbiLsqhCOH
HVlt45UwB/Ed6cedA2TzB4Ht0B1rhawPlkgHeKM8VvtBGeZPw6a8IOgHDKLhavl3fk+LIXeRhu0A
/mG/lt4n0MfuuYryZeY9HbemIR1FHONHinX3kGapkDqmcsF6VxQr2jsQSK1SURQLBMCnJsTEvNg4
ZtwoSR8tbQS3tGJPcXIvwCN7O0RfqgpBp3Y7nJOWZmghpc0KEdclWhA7r/Ry4oE3y4gqd1FEgpVU
H50XEYCg2KQ9RaGsxkpi9RSm/1Li7FQaa5h1smTPx9lVgoQKoEknUk6WbmFmeDFmFPMMsmC4eqxA
1k1eMQfWxoQI/BMiMY5NhRTFwJSG7rbtiHHF9+CSoyOC8XYyzZlKDE8sPGpDgIzAvCei1DeH2L8U
xrzudMN+MY+PXNXghljQRk3oGRNoAtsz8Qp006zbqwxX1owCLn3+V4sWvCfr6T4JeY9clX9dnmb/
L9dVlOdHY+12Zrdk6YxwIiTBKDAKdems2r7EELbpyJ920X+n1kh6yGQgdFnhd90dl5YFGiuQfQGt
mI5FDKWaQu+kcYAXz9RbyEkzT8LnCwSzUEIexqhZW0B+i/PXoiGL95PdMusY/A+DV3b5TAhigOHz
pzMIWsq546IvD4G3HCbqtI7C9ZluSCwBrjvPvf09Q70N3rBzQJhUXVsDMtS0DZUOctd7ChUw9j2f
2856pH/8UR9QXWo4CJpoKiId/csjMyGcPRQ+7OpxSj/uTiys5XWh9N/Dr0Up7I4Q47es8sTL1MZB
bqeEnrHmAiKCluskHvkdraG7Ep0SXddC5qUx2UQXoAUhsOoawaG0LR+CGLMvQZBFYIu7abWqoAXm
LnLYcF0QHFPT9+xUqZrrDMls4jWSVl9mks/wikmkodTZ0Lzh7IyTvgDsreuXIQyu/AJhS3Aj/1Yg
aavYBhu6AJjtRuifujnmvEX0OnbUiymh5a0JTcIU7sWJzsP3yLt96q0IPtLtGo3iNxysGxRWjsdc
pTV+cz2mfFtN9hbQ3NjvAmM5sGmimshplf+eEEU9kiLxb9EXf+7+vWtApqyar8idfauoO2sUtD3p
9PfjFeLD2gFdqNc0+DXJE2r4ghY/r9rpdnVSKtLEXOlylK3gbJDGXfE18pNu/zVMCkkKKhI/DiAj
dZH/jzvnGXMHbtfsCrvWGl2Si7mRj5SCW5dmyT2rb7pMPhPg0pEWkXKBTUJR5OJXfHlGwLa6hEyK
HtP6sVqdCLYruxi8QQkT8M62qQGeXNYpT8V30Oro/F6Gk4MFbewCYNp0MUnPBxzaWeIAxyZRnAFk
RVAbcTEb0VAKrjzWWy76Y2zYJFMWl5uS8zfiq1vE49wQD5le1ofQVRg1y2GYhDIhniMOIm62Y/TU
+foLwY/bkchj8vP7rI3kz2GTZFxKkjBsSEicf8P++A/2F2rozodW2BqOF0FeHXyd3kQjdqdJ+hUx
uor2I1bJ7AzgEFArCDW9kVUYfXFhInTUbppU7fPf+v0DNhMiiqXVb3//EvfDE5+Ay2Qbx/wJxKiG
wp0wnWNEinNuMa+//Y4vq41v9inEjLpnGWcf6EQnCzQglr6TuKfoI3owofTtQL3+OOibbzs122jb
YpOlEmfkMp2O/NPPJ5x6rH9FkHZ03pH/JVLhM3T5eheuytV9/ZzacdyQmOiEIylgN5V+/Wf76Lf0
/oohAxjhwfGmvXntvobAaCJHcXs6NOw5inpi0k+IacV2GGBUxjmwnF2a/OUUvP2erkVKIxrQZeIA
6t4miMQZBl8CLNP3CLa/6HinM0NgkOoPZ6ja0cZCEbfs+D1z20w7wMUV0L7A2//Lrw8hjgRqMNm0
deXdBxxkKY8Lzdp1JPL3GrqD0hafrev/vCui3jyFkcTfHdB4MslqhNaTj61cpwkDYLV7QcHLU0Eo
kurx40hbpdmxgQEvFUPQ5pA/uivP9CQj5WOfocvNV0MQG3PhSSIZwqCdsF4zmyfNLJEZxpi/h3rW
zLX/gydm0dZ7Vvw/5kTtVwcNzR0ao7/e/DBhYrj3/C+qOLhEosO65KINabcEVDfsYAbKOuOcVDNk
Y9felhHt6wrebtCWrWThNGytUfjrITqa0ju6ghl77kKLWHey98NeYJYxlcUxwTUJpWZJvBC7hLj+
/7sdqA7L+LaO73WAHRKY76qR7V7qLSvXiAZRUSfjJxXNG/ZhRG/HwTKbilJ2Mc8RNCBqD11rMn0b
JbsTfkzKqmjfIKzW8a3/lv9/yHaleoU7XqLiA3QMuUqMHVLX5y324VDq+30PX4fgOBV+ZnJz9Xi1
piKATr82cLZdsPM1Y28SXtJIUUKZg2K3yHxVr/8TUncVVc4WSmXTxntI/I9UA0E9pRMNPqnprfWm
TbGSidKOL5LkmGCpqN/w0+K9gq8jcFBD7p/bt1eZkvXfc/OUsZkbS6ICYhWc5jc3HGCPCEWsWP98
wgfhzOQQH4xFznDF9SdKzfdc3bPAFfPxkdoG5Q08TVtMpBB/uSI2rijBhNf6zYJEPGtja8TrF4hU
bTJSfoBZzKSmFUgXwwihySnD/gFyhVPVubnsOnhotF+rj4Y2wDy02SFq2Or7dwV9Arnkt+Z7giQS
JG3syv2ntgft7AbGCzNLBPaaYEAhLEvnT//ha4ioQJxTGzZydvEsirJHz5zMrhKwY4EYtaFnGRYg
GyhBkm+Zx69Qgtn4uPC4bVimjlFS8VLFitpojaw3WwYdwmdw96bPEDaznPpp5Tun/tvZkLStcj78
Ms6jo2nLTSdMFxLp5rzErO2j5adPZ+pbvmd606CWGG79OXAYY8tHNu2gpYeDtfdustAohqC5o+HJ
pdEYlQUdvwu3olIUd9y4J5Z33cOT3ID1oXFl4KWCnLiUQEICPG4LU+i0b+1u4lhsBmpP0Oekvls2
+1t5okaMjvSeoxlnzp9HpmNnLr0n73zctnhbxRM1cgnkbC3Uzw2W7Hw5iH9w528i4LBBWjpK0Yyh
y28838IRZq4jm8uLVrGG09jH/PmbDVZ+8/qETP+RiN2Z8wPTq/KuiT5MVmNvL9yjjXHevMl8G4G1
6gr4ziqPIs8JFLMULGyWqAjuNgA3M7KksrnJyz/wFbs1+lw6fUdfZLPs02kIGRB5dfmZlOjKx++H
Sc9gQU0YJfVxTVzog3VmVfiN5QPN1SKTuocMMXkhq6rkQdlN9zb7uxPE4ldlaxb0wrEAUXxiMc9G
9jz9xwfwT0WJn0HlHHnPbw598KePtoM8KROa8ZVKcV0j2RVp9XJCSP/D0lKWSCjilKWLhkmVMzxB
T9bbut6TInDOrDTAeHDapqbLwN7x+YDsPHr9xZYY+vaOL4ZMem6PWrrmhxfaHDG5ZikIomjfItno
KK9Owe7XFs3+nt523kUa/M8+rg5lcF+0wyWvLStgzUEIWehQemDhH7s8dEFdcy6VtJrLs9qeOxix
A8IEoVvR6sJt8R7hYS9ufo4XT6XXZ+S8ztwdGsymk1/D2L+8ByIsIdWUyWq6dlcW31aGckd9WUqK
/Hy6OF/46QkVl1Veq5cM9+HW5h82Z+JxZqtEgxDF2Nz1SmVQXuKKIv9HSLPG1g/UA+4Ozd1lzb9E
qmME2BuKJXXrpOb1BhWlw8+pqUnZ50GKFq4W3wzkGXUcj8VGCSNthu8L+lWUJjPQB+8agImdHvrm
aOXVOIuY/pXcYsM64D6PgROAHzAkxQcneNX1PzOOyg4IG5NHjza/EbSpGFIsT9RXWKWR3qtKcdu+
8L2wAfXXCddSoCIfap9Pnd7uCv4H8j3dqrUYtX1Yn5GxOe2fJwbh8NB8BUv74cF9hF8Za150z8bD
TM5XXINnjKdULkk11tSqH3m7gMmolCDPNfIJz9OTsOi3RgfWvE59BgX170PHmKZMlW0vSsKl7p+g
jqFOroe0dbo117P7xNX6m9bCNPRxct3+aqjSDwSmUY/CK5l0mzE0kxOUx5Of6Z1Awd984g/rcbZi
XeaIIw1WZli94gZQ/Oxn8uXYRN2fZ05uGR+M80pdXh700Z8D8cU3/Qu5jR4qgqkGwg7zvlY4cklr
Ya4p54LKBjAkXmDc3RMh0l1DgNNpV47IUG3hAkQqT2V/PqaCtePDUXC4QYsP/2Xa525ycAiv/nSb
hubx+dFJFbbpXghNxiawGa5SYrj62Ul43vnGmxlFdAsYmZ0g2Job3lI0lVSeFyg6JKlEKyMf2yyV
cDho7c839mn4vGCjC4Aldt/Yve3U3UmJ+LMhkyMLXMbmy357K4riEIewApFObBPzJ3y4/zdMsctk
T7PmrXfRhPu2UaOQ301eS2m/sNX2cfZq1sLvVb+Uo23IPUikeU/5ZA/F3UGyOeDWjLUm2Y+Xu94x
q7bUgaLjaIwRyo4XEO3NILCjoFTOeFGk1x2u0kFnx3ty+5TByr0E092q4qrhabUeaiyV5Hp+f+03
v5bKfZJI4y7W87QKgXJ9eLf5vGQ/wYZAxowRkovADbho1VeykJL4AF85eibUj4NJjYRClQXX6g0C
QSW/XpUgLwtUeHhdvzZk+R0/Fisc6Q2AQTujuIkLQaf6oAarL1cP3XKzJeAzop/j8ogq0DKaJ/bo
tsZW9wEYwIi86s4GcACD5G0mbGa7f77Euec2xGEVXaQPh4sgalt8qKS5f5/WTLMYkrEun0tK6LvA
rk553dhYAFLqQ7ZbCvX2odX52gXBsHBipnaPpPJ3MHneYzCTBT7TttGYqC+09LEGvRfnVZeGpZv7
SGQy+V0mOLZ3s8vE92sHltfeoF5T8DDXzEXbsERtmw+FU3+dM/GXzobTIQrl1lEiGqbGvpbB7zFd
e4YWge1O0QUqCDa9z7hyZs6ehEAw7z+aeYoBOEBz3V5wRcV7cZi2Qv/Ns6f998nio4q1wv+BItU8
G+pRLZphrsnOrrFN0VKaBi3S5hcUx+86uqK9WgcQV+P8kJyXPxTiPnw+9clRHQsQXZ9HEgWmWmhM
OozMo+w+lEEo8gv+rjjGyvh3dh+ks1A8TP94VUHJK7s5PhCamQXFnza0Piu4V/rEwSSrmoo7l23g
zjRMjZnn1hzY0bV++hDK6YW1kWgPoS1os46bwKalm4QfineY5CkzI9avV+Mw90pg6mwR217VTFUe
cEALdC/e/S0Jd1ayEdfeE5suR+bx2U7+LkQ9E4kSPvldmb5tL/h70ozzl7MqDzImtCQK/w2ZttWX
u4uZ8IN8IxUcbfRwR70qyWENleW1KteevCHay0bRBzvBzi4vj6rdIH55oM5D52aCiDd+ya3HQ2SW
7uWhDmQDlD9I4WiyX9zwSemHuxmUgDu5lFehKZV/8uou7kRsTBDlfLblrE2Ln94QD7WS8jzLP5op
QnaSp5o6pZiY+LFi9gRPXPTC6pqynABfP7Pqe/sYgW051xw8oHOeMACD1dHFwZ+mF//yVGmhdO2a
pQlfPgPzyZWwvpJOaewzMR7ERqc3v769oII/0y3FGVdBUtyNTUmo1t2Oecpz5TgteD4qXg/nqK5S
tTE0fjrB9pTrOvPgSzRSAjfbtD9V0oTniS4lWauoIFn/hGJP4IgkgqRdV7ED77PLYe70U9dvWd3i
1n7cecTG+4FAhxWKNqq38bsQKjSlNmPKdF9BR/xehPlG1ecp9yq+hiiZNpc+S3vMLEz3qBXTsAUs
M73Wew0a7wU0YOqhWDEzr7EObeELztIlO8TvuzhjtSWepLOp59zj5FEqqxZLrHETLUbiY6CkesZP
wDjkRmeZ3O3VJ4Vp7FqUF8yu3jAxgZewclN02uWQS3FvO5R8ckrCmQ881AIhDa1CUQeRgU8LLYZ+
zCBNsOsajsmzyNnFQ/LAg8i3DC0EdYqW5WxcfkUYzTjEVDxoWTIjL1XTYGUMscLJIXX67I/D18bl
DvC2m1Kfcp3falTkUo2PZFlOoYh9dlqyth6R4dNqhh8G+hfhXhykV8XmUWSrbtdoAJfYIq0JhO1H
cwKq9qfTSYMnAueLsI570tOxrzFjzcqv7YEKaAJDMecT1e+JtjJC6rD5Aeo15lhF9kvWji1uoepM
tCZxT8b2jQ/UQuLvDMlfWHPHtbehFbPu92ZlMF7VK/zYNcqt36u8mrvJB18mphyBZcPDLfCuQOP6
1Gua+D4AgiXFYuoVcAP28jfdJ4kSfVmPq6XalAXSMZEDPzsLRKdbjrtlC7ec+RARzYKZJs/yCI7m
LmcrJ5wPGoFhy7eboDdTcFVTlRaA+Ud9mS0FSM+L4Y9PNPNPeNZ9NS+xbWY0DTqQAFoSn0KbyaWt
8CbDcBXsSM48hcKCkineGscmJmV+Xq709VK4be2rug0bZUjQgZ8sacXi4Fdk9ULAWvOkMfcHztxr
uayefJRJlBnQLO+PNwnYCNUnPnQ0WTjgG6KV+B8LL86bd2CpnM3LrLsii7SGhRf5wd/1UqIbIb6r
XhXPs8eMtbM57C9fwCebN/N1KCUT04TnX/jqG0gLKypWhcUaZqp9e2ortJDuFmR6qFEZZe1wg08q
DvNzFpheAcwsJnFzTtjTIOYi9faSIE2K/MdQT98PS+uKYopclmm+n+1shshPgm075LEsQQX/N06q
xpvunbma+Kr/aKsscns85OPbCYDsnQl0xdsKL7osaQ9geSaWNnBW0votub2N3GNPDGxlzzBkJqqV
TJypyQSV45eq6yxBizzDhcTevTahz7ytT6sSWgjqIXkB7zADgUQk/w7fngtt6IAdELPqmHpo4n8Q
zsdHbjjBuAAsvlgsXPQC1z4Io69QRqHdmNPxPNm6OXP04UjKXsFbk0lGSE6oLyrT2xl+HlLz8v7K
WFsL3Uk9peG2uN0TfQBcQ5YbASP/W4LmSUgl1kwtXD8pfDMtv4fB/y9mpYtQcw/mKZYLSmuo05ee
LBL6pecrFxzSD4WgHYlio4+Bf7H/MlUlX07fBxk2CB6qwFGnjYnkfObpT/rHnqdEx8BAIJy9qzxm
UaQCyEIVh5SIOdx31gsCo1ELmssB7FNAVI5PTKEag/0FVrT73pM36kUBMgNMYtnkoVwVEdleGW/8
4QVJr0RMT9ofF53ngmuD7cxleABMNe6jyxdk1M0WKJoFsmp9HXmpNrks3XWSHhzj0Voe86kjNLeR
2UkJBLulKQmOa8xtv15jxbuYMpZLc41Dct7YSC8sN+7GgHMinli7XncgBFKcFesJAQHXbCqcQ+Al
CgQa3BcPgLPCRVR8e/5azSiHUjtJ8nprknBraEt95fK9e9jImnM+iz+YoiZqkWyFZUi6qTQwPQU4
pdOqMSUClAUlWS+5jeqo3PvpFJ/gX0jTUSFkt2cPeNgE6sCBjg/gLQshLrmU2LJOBOoShHZN6WsV
TRiHSnevcoR3afIpU3UFD216ORjNpHkCOpiqjbnMbudzzowbYrOhaL/wrE7gl+sjtpQdRFovrXMl
ddF6gDOI+45+Ltnim9YIurNBT5hcZ4atohjSEw5evGv7WvuazhvfZOGEb83gizc7Apq8gqILjdQ6
D5k7mfKq+yjCKBp4CHp0JfkEXumHxYZMIgatRT4fM+B7ZUqkrGXmq/pKB1WajIZROyrHeuUAks//
n2z19Bla69LQvE4ai7faNIhX1nD/hLqMsWYU72BFripBc2sV8dBCNgMLkpYjsQtdu9imRAfZOz6s
1RHJu2ZnlFzXyyt3gMOYxjffoWDfgi2LjOTLusGzU10Tz4CyWn+Y8OXmHeLkB88RpsbM2hp6mM5B
Kpgg3oPsL7UfrBJfVrRxJcspglI+MfSeHTNHK97JQ/uTe5EK9QSWooyvWZESwXMHbB3W4dbyTo1W
8f/vkRfvdKo0wPGLu01AMKcNAniK5jZy3fHGKUL+dSA7VtHQJvjeh8Ax5Co4NK3yNz0nqH9VPrkO
zD9Wdc3N91GblBBEmCJthyzdY/nnJe0xeRIet1iX4WXP+ZI8epWwVQNQJiJr0fOd3Q2Zor5yUgF2
HRtqV57t5cOwrSgltz/NMzuPRTVW1uYRB7vfB7pNrn0y/D90+zENUEC6i2IXDTDs9u2HAwqJPNcf
+Q+fx0apvlfb0mCu0C/t9+G8jeGKKJi2k+YmQ+kAulirz9d8zWJ03L1weS9jJcxyZ976UpLBOjAM
3uMLQ3ptlhOUYiG9Kck5go9esW1d15SvofhPcCsJAMnyblOCYynWTuduBb614Go6Kv3a5DcdkoH4
b7jUIaYEYTx14mezi8ix+xHzruiVmB/QTYhPCrg3mWghQlfge/RK4J38Mi/91cZ4+XO94cPM4VQ9
P7CUgbVIcV2UjmLk7VAezAy8XSImgN4Ki3WvxknqnFGkcFbgR1+iXGlJzK+0OVn1OvXqaCxzKCnS
+c7AeHRkqvLRnGrp8hr0/8wmrFaU9YBgl/t/EGg3LcZxSz8733+A9zgNpenVugDTOAkHiNfe40ZM
s/ktqM+QxJnRt1B5gv/QRPhthRxk6ANvTmg2DB6R/KRE9ieruU6d2TjoUEZcqnghz+2EjSB6TXmy
IkZSYe/m4hDw2e3bjj6CH2KtVTgtA8Zd4c3MUA5r7snLiuTjicDFwzisyKD5HMiLQwDlCsFzVlKG
pB/XRIfQTTbJRHjfEG3ywFso29IJlEHQj8CtVFayuayQvDgH6TMXEmkPU3z+63hIPrRMnkX91UAV
p3nvhWy09RBixd2tpcUYU0lGYK2IwLa+ir06eg4K8siyjPCC9egO5cOsqmSNSSXkWyoJrhiMPjnm
YOqibDk+TBZE4ZUUZ9W6f5YXesvqgxeefsLZyJ2a+PIKJSn1mR8DFOsJxRKG3hUS62jH5C3DfeY5
RHzSe7N4DhpErwVE4ae7IVYmfA/pDwy05IAiWpYk/Pk3JGzDDLm9MoS+4QZOxcoXruGzSn05kQTb
IynrQYBO4sWcLJVV1AA2q1JC0IB5v1iLNBOU69FbEEIuj85PNagDJZV7DFqLqdStnFaPNuobTP1z
4hcq0vfjBP9B77p6pPlpmD4KT1WTwA8k/31HVk1aqAfW27rjB9+/VjVx6H2q4Ld70uk8ym641djT
O7zttk3fMPoW8LFTI9sJJwYWx2fksGrHhcpT+orXJYoYkDwO41Dc2tb6lIAOrTykGf0yiEG6IX4T
dGJJtZ75Dczq+jMbdTSJp/XAxm6YewcrEitgBIx1sQEDx7+PxUviBSdLC5lBAUkzOkX9xkYUF1wN
oUcMX+IlH3GnJKQvNQXETPAnNMSnGEozZjcVOKngI/VhuQpcgwGF1sHAkuP46wqrqBZJu1MOILEr
5vAO7wxe5sXzzHsTdX0lVxlowBi5/zBLP8lDgRAKmGhsvmXbVM+h19A/ajv0NeSdIz3gumvFAnzz
y25/XBMCMplj3B33lwBP3ar5cUTXH3xVgzKB83BlN/l6L781KfRJEji+VOn7vyOkQIkQ/LG4VkJU
/jIa7jfrcmQmXvjY10YQRN8W6g1hXkNzH2yUapn1ohi8ngsuvzsmt4ctLAUn+/d2wLECIvbl/Uuv
AMFBi1pZ1QrisXrmlTvT511Y/XhcQw7N6gDQui99s/09rwjNDn2X9fIVBkPBiuseKjyvKv4g6BTz
zQCwRkv4Pc44saCCs8YxbUHN7KqslF3wG25AQTCzba+en4kjjiCiz1ioTM/qg8i03v74V1WmusdA
lr7s+9DzyniYIm+Cw6tWll2P8u8ciNoiVvydHXU0CTsemv3RPtc3kDVmy83UD22ENr22axp1JcY6
eJYCr44FVn1f6btW/yaqNUDl0qdMEaRjQteZXq1OtYyq2KpSsYkQDBLHZ2MaPUdc1hTCZyV0Beos
ivCP8WDKCAbpQQfE550As0vlo5si1BEgsmC/sgrN/jgaCjvLHypFqmDPre3nD0ZMow0trgHhnJrK
PBC71iohlhOwAlsvyg5sCDAu525tw2shyO6ZMoGWAyIs3tYI94JGDiCQkDEaoPizhYY45rDyY/ap
lMOQYGVO1MWQQxIy7lG/rN5dNZe5x2rQiqbNKcHsoiJTcfO5360FxutCrcXiIGT85umcczOIv3zP
i146VnDw/CAJv8PeeNuO0g8g06bm3pj2w58iEmJxEkyextIfzLMGN0SeFf8kUs/tpspRAz08+m20
InPsyDxq+sP0L0dOiaD0yW9Z78jFpn2fJER1yn4fViGGZGzEKedwpImhT5BJxF7nE8NbAruMTk93
MKySeFClfPTYhZws40+IDPaqkICptbCiQmy93CN9ajOyfK+YJ2EOZeLp6ogzXuPksxtNv1syDSks
BBUDgAjMzsoZ6CfvImitJ3sY/CKlfca6Z6BN2A2VQcJQw8Rtr6yFE/8vqkMDXb07o2Jq5yO7kDKQ
0yKMOMWy3M0zicQFAXYSxUdBcL56qqeOz0qW+V9Eg1irXSKEDkbNoUZdQ3vxZPqsWx/zoutKDFVQ
I6/MkCoHrXDqJQ3xYU4GPPK3i6K9XhYtRb17C42eJPm18Xe+gNS3cBPCQwCrMhRJtaytSm3+mNYa
pnUbAU/UkC5qZqpvLmT2yoiZMZ0Lf4jmlORek6+6lYnVw31UGFZ/Y4ut8nmtSF2vUg9NaGq4rkVs
eO0WY3fYFyPH0hdJeA1+9fR2/oln+mzLO5P9dWJJ7jsq2KFQ0WpyE8vSYalwf25AgJiLLsS/YS5E
FoiamQQaaQnPcZefUCFu2oTuwGwapFEhV1a/YhhyImnKepuoErPIUCOc0Mb0vN7mzdv6nwfyLo6M
XCcNPX+qqusdvxLug8QUosfZEm9k1/Z99l36sXw4uC051WFCvFSayP45neLaRKxbqmeIKqclWjac
8/+xaW+7WsGTPgHG+F3id4zrqw+1gvwRY2dM6ycGXsAdgnlkQPTB/WhOzvgJ2gBKQwZujrTaxD8B
oMQ0GgjDOQNhMuVx8zld9Cl3ytp+lvARd2BTaMJwwzK0bjjmCYSAvgMPav2sLtYmopOYxR7zYD9o
KBecqMuZUIgenHUn/kcaU9JRjjae47p90uIWB03dqOmYfMizWsKB9km38EFp3oBalp8Z0EwPOE8h
g7fMgrPHKHdjHC85fWxB6+eMDUa5/pz4Lb4KzwQXiiRGhI1+EkeL+tqTU/ihOFXovOIB6cvTelxs
hGv13HWB+0vkYhL5PNhkNRPq9Ix4edczqScKSeKTyQwtmOjXWLL5krEqFjiHTtNCvIwHku+fFXid
z5QIlyn7LyASf1xIKjpcQVKCoqKNmM3QF0GHi0EFbyYB5W5XTkwKr+el7tAVY93RxxRs4eRUtDmT
haCN8KpHn6utYr2HhmyLPy/l3jChx6KGIDwHs1MB5VNdU0wdJwgZI/dVR0GdG8rH6Y+2uqch1naU
VEro+CeR/FdehNCwI8KsBm8RBt3lG/lP0N+cJ0SXKwTkIfsOI+Pa3RXxRclXd81sp8OoOQ+jrDAI
xTOiYiXggZUser4VbYzpY3j5aN2WdW4Vyt21kGHh/cpiCNXV1T5lEGYXBaIOzaZHsc0I3778n8Rm
BhH5H1RAU1n95CYD348/p1dmS3grAosysHId4xvT6FFUWc9R5FYHun+Fg7pw2n0/n33T1RN2CEIb
6atZBvCPNN3mTYZLcAiJxEdczNtTlgxTfGB6Y5P9uRJo4KtdnIzKGYhwogf/+uFBPS49P42Bj6kX
WGoJxgZz4A/Kaci8+L4mZLiZR/r1SU1gcOR3K9bTXkOzXMmQmU+Onz0g98Ly2SyEYNT43BR5YAdk
v5q5J+1hCZMCsfzKTCx8ChJux3vZC6HV+NMDYhCFK7tCJeBoZ9IvsKfQKi5UmO5njeQ1/VRq2VAS
3AEGHPtT0Ukp0M+sOnJ2S6E1YYFmeBQA0M036SDzzD4sCMdEPrreDWYGnq+1dVB584PB2Z8QgfNJ
jnArM8wYBRe7TMCRj1x0HcbJohUU+Q6EasCbj41E/q4fjJ+xuwXI+hqJOWkIjCksHU2dMakMNv84
bgtJKFHgYnXL/2eO/THJMkFhhOQEMwLI8Ts2UF/IRlB7JOyQGdPWfwZwh1NVoeT31zWiph9jaJfn
EJE3xAoQRmL/4cn5qHhkC6ymrRIERhkWhSGruwPRBAxonCOknaxz9p+ghh6SPUfT6E/SaCY4MtPT
KJA5eVmOA/SSrV4lG41gkJ/5Sl4und7Cp4XqxnAk4sEGlEUgJi+mBSrEWI2vvrS+u5VkQMsPnvXY
83Fw5IW44WUDGUhNwU56rQMheemR2jJGnncOBiQlHkE9eR4qe86qwBmugn+onppKd338CecfI0A+
kQW0WuHHADW2uOzRy+uIZoreKb6q3mwrhTqhzwqnhZ2ruhxdeqami6VWoty5LPzhMyfhptv3GkPH
gxEmWOKfnrnXggaLIpjxng6Q61DA69EPgKDBYNRm5SQRcHgBUcfOyWz7UrtDmNH4TFXFddXXQK0S
DZ/oTYora5VnutXozxgchJ0KNOHENtXG3Nfmxgb8WBVbBWgRdaDcFbSKBH8p9yn16EUq4oPLQziw
EjtDvTduH2USc8otSeHZ8XKPbcemZaUhEP/vlykl7czdFFHXsqvP0ZWLSBFCkcm5+KF1pSOFFgTG
od5akQ1hkrJVNdF37x0BVwxoGSnHOEehOZvjgyDab1UCGOQf5HmAR6XW1+EWGw47ntCz40nC0444
SIZ0rm5cRtLaH7Ec/cpuFfeiU/i1jF0l54T/cC9RRo+gY7B2QwwUPgSFXMnZFIhxfuxTZ1NpteoS
lr1BAFogDE4CYWLm7py/+HxfO0D9JrB0iVmhnvhpyJzEYdomMLU0GIyRxKweGHcVRXWjxcSqsrHc
i4QoJPoYxU6zJXIKen8eBX5S+9RnKk4lMAo/TCDdiuPOrxhN91LPCmNTBrihvZAIl8csvH0svwx4
3eBu0wisHgmFwXCV23LFJb8OHI8sJekmexjGkbqi0CgAIa9UiuwPa4gQLin1DsXeersFz05o1alK
MT6YCU473Yn38cfC06AkCat+puFdDaABOsrtTgMN3Lr6RaQIo8vao1Fisd6U0lHIJJBNyOUybFuJ
k7/RJw8JLmk09sHxM44L9LH9h2vjd1Fw2QCO2hftZmrMpQC+ji60snMATPc6mpNluVzvoonBz9H0
Ze0ACxLC8SQuwj/txHsFPSSzBiAQt7alU3dFnPlifp07+X6ajz+vHmADJgH37ihWdg63Ligb4kY5
/dl0yUjLTkDKdhfALty/0jvSBD1USzSPWqjHa0uTns9Bp5NhMQudpikFOl9+LhUpF1zTKLCxj01m
QAY14Z43wOn85f+pxtklMjjak3PEfCzEx2nXGoqepdnzlfRnsj4KcNDKfRabZspO/MLnmdhwN5MP
a72TnxpaTvIJPf16BGr1JoShRwBIDqJaXYnNQmyP7uDEdrq+13G8Vm7+Wwz+0P5hxTtcyifO4P34
rgpH5jy69Muv2l5c0m83lsOVAUkhDL1HDNbsVpWohfuJu+4odAfgH7oMK94NPTk+jxAXDp40ievB
oZluw+/96WB4Qq6F+uTFHlnDNk39Xbhreaz6woZjmu+qXNgNr6B3o0d1VkOdkH8RrBcw9+aHG00Y
5UHUFnWa+T7Wc/efzXuqtfcvq3VMMJUgok4sEqJFe6QgpvMyt2IK2OHwbixiebXSs88T1VANS3R1
c9FgU970O15D/Mi24NGtRAt4ZSrF3IdRT84qhH+k00Wr2LAG4OzrP0jfjdtV0HJwMDPJWSTcVJtS
Pj9XRv20pl65wTDkmNER3YT2/Was59mBSwyWp8cPBNeGlCg9/v7P2MjDgXcBGX4nu4wCHhysoiRU
a2dJRKINa9s8MKREI52wOrVsahnv0MhqsS9EN7IFX9stF5EOmKx9CUJaqxmlMSQfG5V0X6G3QV75
iStQqSM1mBUd817T7oIT8AUQbNhg9WFG9cIRz2a7VHw6VkWU3IgOfCDOJVpz1mZLJA0PGaAzzwqX
SLuPkbKWAxGljrmDfNpM07HO1yXWxiJ/jWfJ25zBOE9q1C+xDUjrhigBO704LSWKCtMn6BOn0OxC
cpONV3UZVYPSSTiEMLDS1G1eaexUtD0lmkZ2goc3iw5Mt6SsCnFqVf1qvieTnx2MW3ut4qNYAo/e
Qh2aVsnVsGy9VvpERQf8f04M1ckqqbjvW1D562prdR8SZXtBKQPcUb32V5ZqKHddpodc5KW2GuIf
u0pTbMng+vDZ7clSD8ruI3oHXU1YGuQrh7UaaSd2JP8KbzIlyK/hZ4YYbhizUvTWjLRbBN3p4PdV
SwcsXn6D1beThC0MXgJmvTT1TqEb6lI1rVaCTT98VDw/6tT6YO/DC+R3wAx0DgKtdU6x+THdyocE
Wdk4wM+yrgcFkS6M2v5fHcOR6fJfp9Pfs8CuXq4O/0vVMasn+FJ4N539EnXjdOZY50RRA0ZnCydQ
AWITfdMER5DMfJrbt2IeS0A319Q6aalHx1yJXgiyYZ/TjRpeknvb/9pOimzTcE2xZWu1NXMJBLCx
fNvuD/Vp2lyK84qXBW+T2a7sqFEkBAIWj/7C5V/Mq+uLdkruLtlGbyCNU6OaC36W81bmxZgjCE8E
dqwdjHkSwXAd1vnRpbwUNVAM9O+tqBiE8gL43v6JzfE0xnN/Kk94w/h68y5hSG9gAH9/1xK3ecG6
gPEmqUaRsvXI/B5zGFv6uL1Y0VSL1SazEoFwFDeI/eDBQvtmk0LbC5ed1fyR0tDNUyY/Rmbc31wW
+r1CGZ8IeaOOQuhXcKNC89hxYBz28gA5a88o1x+btD43Y3xEhju0U5PdcNsMXsb/ipEV5j+cOnVv
UqtmfFKcfegy+38Gtm69P94bonaLAioGFgiQpe0QoKfQfbRXAKvdaPyCjComE1qC7Brx2IAT7GGG
UosnQMvdmVlMUdcPf5JyLecQ+idYqsaR41ymkH/C6ZXBCdnrSPTxg0b8MiKYWyvt8b/6gpx5XQ3e
qUIFeq39hq1288C5OIYAuesB3NSqUYSpuEMEgy/WJxbcm/Abqk4X1N0eqxffVc9otcDdmA8GT5Ix
Z+kHPPgervVUXJZ3fuONGj+mM7tvIbuFAf3wfVcD+ANqKuZG8ViPugQmea7wO9LHxq2uSjksrdhT
w6lGnF91uJDJvkDNjaPUcp2zNosv6J7uLZc4pCLoA2fZSNiDdDg8gs2IHZkpNxglinXI0M/h4lTJ
JyCvthOkDVCY/IWsyCwpiy6jQgAQ1RlpYIm+TKOAEppgk5n4hejfrSA6BZGH42aCDxo/ExZXtMFS
BMYdV5HJvtvtoGf3r5JxPZ4bSZh21g917yr54UtXDulzX0UCuVggyIIN1UTu19W5uK+zgVfeWcxO
oJTxltGkA4/i9MwDKdSg3DK784/QIVdjyhhv+BpwDo062krfrh55P9jdcM6Xa5efxl3WcJ+oSl4I
4rNrbN5wkH4LVdEj5PoykF5u59HpUoNXc6JVzWd1Sl4dqkq77iE0W3JLL0YNEaYXCrxKSK5WgouG
s3bsc+jxsztDKnom0T0PShBq7is9BdEc9t0vTjfLbTEpBx9JD6Urj4b1ZfbSBO7GIO4SMS1WmAGZ
KfFJKJkKVEHHZ6wLs2DgtTvuddZrRbTdtjw1EYxt2ivTQOfBe6Qp99gi0Ok4Y0++/Vw1zVEFOGdz
zF7MKXNVc8yS+jYNS0omo1KCNTCGpfgVRrq/wwYA6SHYdTDwSSj8bYq0yAQcBcoIw+XL1tzw1PkU
6rKeschN7PEH919yPg5SLsKxVrYpq9QdfFHsEWDhSqqeh2gCUtAG+U0SawuiRPJ5FhCeq0Dvuw4S
tk3Hcx+OboDiwJkn/5qZGgsUHMmc/WOi+3uf9QsX7LLemuepa/9/NXnkJwZk+pJBEqRCWdXqZg5N
PbV8ORKGvzPwzaV1XhjztTqxdiY3PjawAAprbDOAc47xTyPSK0x2Eli0QSxEEXd7Q0m8U3W/LV3L
MNu4TJK+kIDjqazqUx8hsYjTAvIDVjtuWHYQot6EgP4IfwtH0oGtKuwcSgNA3uAnXxqHnGR/6B0f
69W7/tH0GVHVN1psSdnYngF5lPC5f7nAOM0Rkv/GpAdkg5s7HHgNPPmJ7yHc1BC9yk8CBPndsthM
AkBjsGys1X8e1Meu7/OQVK6Z6P2OFKCCLXiqvLpADLpTjYIIfkQSyv7csIVLAfH6eDd34v1a1E+9
azoV9xa3YIICwus3OYrb1CeoiUjOu81ezOpbxMBmk0mmt3oxigWPD2ImYka4b7UYO8NrOwxwJ/XA
KWiqy1cFshyxhQ7LvoxcuWPjSDfxXpIOuvbFO6KctRTrgydz7/aLPkSrwweZueeykVrCTr7Z6AxH
BDJlKBMJE5l6NUpGbE3ChfqbKh4dhCdBVoyQSKb5kXNGkzNYu8xTKQlC2vLWSObgST1ZMfXtffwW
XY1gF7/ldOVw8II71ULOnpLYvFxNrerQXJm6Jh10i/vkRmNSW7CwKXRSlxKuw0/QLedxiuZ6iVGe
fwf+Dw62AnO+iJ05mNWEzmUinfPWRf3NBsfmXtnKTFiTh8OPRzh3YA20xbjwaIeU1pQv4Pcy9A/J
G+iBC9XYdo2901HeCuH0S1+kZWsxxHtKNJ3o9qCvfaLQ0plX7F/fKxomyHXZvSIlMvn3BdLz2DNt
+TWIMyHjzmE7ZeOqp6UO/nwSdZ9NX1gK9zDmr659Lk8fzVag+QkkdBEWCMv/j1+rhXCa6tJjsbe/
mI2O0ekBezXS3d2j2uMqy3jkyQkym06Bg7/aPPZf/2eBrLbP7A0v2xeFbvFZ1WHMNH+gk7DabI1e
IDoxQ9SqeRpC2qZMDoqd7VEZaZz+DQQn0bkQQqKJAcZvn8yjd4safu47zRiW9XDgy3BEo3oiwQKk
bAxh4Xe/UWlNkkG5Go33iTDKQlxSkVAqaPX6WSJeyM5+zyfRqIUXJH2WqVbct8qAJkfdLBuhQkrA
u1sq6O/6vnBg7BVp6s1rkOOSBNxQzgydnfCxtj9FcYx2aksawIyYD/fpHzZ/1taFFFEsQEUgBVeD
pZwLG+Ex6QBSRU9JbuC2oMW6FQ5qFCOS+4VFd8s9H+etopLQ+pU449uZvWYustCZNklKqIW1ORfL
as/z3KWBkI6Chu3okegrmOLc5YBLc8+nzBVeUItBI6fXr+WrmDC9dLIwdTHNAzOt3/zy92xXNm52
qQoMrOX4WKJJ741EJX3OnQr76XB087pnJX3xFnDz3JQh5Orgb/kun8hHQD1k1+N1WbAcc/WQVb13
FdJlqCjbqhozSinog6Yk20vjXtTFns9HHXQ6Y1Prx5LFHFybYvR4F+eEDFfNJt25K/H32kgL2AZn
/smLEwxYViHW/ho/SeGTduZ0w/9hcekJeAyCagOP5pVvdfzhgdkSUTQAlbO9bUG6rv2gZ3qSUUUW
AhisjM00luwVVsUNy+yglr41bdvekJb2AHqqcIlyTMQAJk9JKxKuJA8meye76NTFQ3s2325j68VH
juUHrJr0bJubakKd15prWsKMpMG3KZ/46s6OMhoV+r+FKnY7NfuapckRfblJE7Xi1VqDWhaasOl3
T0hyC/+X5sMsonNhvUrRkh/4RYGdDoGA7bn/u+J9yC+nwmDTAMx2or08BPBUOPSDD0XFlOHCqp0H
RtVS3pYBvsoIBAaa0vvgJO2r2X9SrhiCB26GWzDjk0nOBv6i1d/IpMRmtvfAkXnBqyn8oEtIHmL2
vQY1uF/Kfnuh16gBAgc0wUsPJ012mwQYRfHzr4VwKWfw6mAI2fj5MygF5IzFtORtHJ8TmrzCWlm7
w8fgNdoUwguRAwPUkr/H/fPBixDiKZAk8eLNuKyiKhoZZoJoXm3EIaCNT/lOMqaOTcMeuk61KyTQ
rFAD7kxFZTGNnQJrPc05lG4HnTaeUt/imeE0DERB6zJaaQWO17uaVR7EH/FP00boXfkN+SgX65aP
QcMRVwi8sqdu6HazF9ysnRCOrt9mJxWbPPy2f8s6gX/JVvcV/q45Mu4/CRpK48gwyP4y8ILvKhK7
SyzBcDYkhr1k7v/Ui7WjzXuvcsU10r/e4iDSnFyNoCI5qI11jCqkgz0yS8MYKAqec7XyTpReJFBr
vv+myvgnBPO/AHrXvFer+LLFBUIc+vn+x+3CFgjcNFtGM4dv0uw1bcP6zwUhvMFASzQV2RUmyC2p
EJE++B1LXV/RyTQRCa7EdqWppjvmnGbLHcAF6oVfdaWJzAT30xsX3gkudXM5Tqhmg2SRdAxXCK43
/MpNxFan+ITNq0Mj7KwBbJGpDBixIac3z+d8fYK0nzAaOXQs2XIbkvkAAjsx4GXTSyWdIJxeUe42
h7HpkbbGbJJJzN8eqvhhWTEJTH+R5+KMozMnljxCILdkmxCDudC4lUNVVPCBEjK46vakch7PZzwc
w/hjTTHyO+4WuPeq0quVk8XH77LOZYFT4t72/yc47XSDllbjMtm7EsdyQLapkrdKVCnHVyvb5oAI
qUY04j3ki5xOF+VO6ebUqikTLCpkKVw2vSxnfzjtlepwvGcA9ksl0vmPhhUTYPuPoL2LGxAMa9zc
i3WpQkj5ycx0/7MTyWZYff//gSKn58eNgMFehHhNLsUR31oOSl6zcbslW5ZOZRVg5cCvDrx9n64T
O4tWJvlQQrLvCZ/QThwPKrewHCAxNcrPrLkJWn759/WttLjCBdVWgEl67vfDzhLvO/2QFkWM+thF
UVH0SNZL2q2BxN+IDGkqZxxR6qjTNLPfgIYiZG54p8N28S8K5qYXLqKKfK3BSEsE6cyG0HlF5/VS
CFVSkne2VD6vwMX7epv5UM8353HEjhAWyNTfNl1AXCtHM80qOzfrHQnSmBP6rHdpM5y1vEY6/2NM
8upMzzRoYI8qAIaSezO2ClX9l2Pfo0Agw43CDTjlyktQKSXfaYnmk7OuLk9aBbWT7wFWZgo2EDcp
InQyipKF0VA6BohbJopTRhh3yUPw8cIEIeYB7mBb+5jmwIlrXqXfd+wLusShjxP3i4dgsxYuRYRl
DQZr7Quljeg0LR+cJL/0VOUPeCaBYIO4rjWEoPbMzARcknrubLM3Km0Ualh6t4VFM6xyl8hIIZ1B
DSVvg45QnYy2YkDUQSvHW3n54Uygf1rlDGrPf7KSnGxwyoQxOgEOXXHzktmKG3/FuwSGAsEJ3NY1
0plSWLYmIBBSvcaz2G+VQWMFgx44gigNs+ki4cPaXWO9utpwqdf31gDHyIOy5Vm+DG1N5Kzl7T3F
NbgDHN2WsNz4RKMlgsiyDV7bua7sjNndRbUbWxLkkJKgjUD+3fVD//x5gbzkls1hq2PTTgo+1Thk
Mp0xTRaTpS87RVj9kJTC4f1XSn522nU1alBYr8XRS3JzrUKnqtV/VOtjEzmTxBxyPotikpq9cGwJ
z5aIW8p/324CSXwKxkHePHZWrub2mIeno3dHLMVQ1AJJPnfJHZpfepL1MJtgpPDrB6aNWjEtu6W8
wPwhvFmB6utUHz+oriJjjbY879OhfU9N8qD7TnvOP4c4FBfZUvYfQFzmsZBCmy1VXNshOPIePfag
4zYl7k+25Z9t6PFoAoL+p3/Gjg6lyPhbXmwqtBtbgM2jqhyLD/hVDVIFfvFNMaPsJeb54ZIztiea
RF9cLdRDV74TyaAKwqu5o2Xgj78EDNzdMkuZQ/73TYq3W7uYMmtUw1N9YFo1PbLn9c6tvk6AEpjC
boFkh4/DNkPmtHWCzKpbXUhPgH1qYo5y7+kmxUA/e8o/ELflPK7pR2r3rZChjsh5+lzztyrzwjCX
nG8p8b9hrAdXPhUAvtuIx+ex/QFBXLUnRgrr1riK4n+V0htOonEpRZDQkRb6SNmkJXMAbr1Is+P2
bG8HMq7KsOY0M0uVs2Fk3bFz5clcCEQpMHiKWV2j9Vck/jD95eLlmxYsOenSH6jHKC8nLzia/nFE
iIgNXNEPQPwwOfZ2RDl3edwEKme5dQ1owm5+WodnBnpVnPwKnZe/aJa0zJVaRmj/qu/bGvyXYzUG
bVMTo/5dSE/q0Q7AT9zTs4mrmYAEDy6PowQrbBdrY/JQxceVNcTpgE/DUZs9k36QJ4EhG+6n6yIV
+iLGkvvun798elry8I7Y/XRmPKM0Ywj8YPzM99gxWXaJpuoPGaYzPAW92D8JgnBTrGWtGawqyp0m
AHOjVRjdetDMdpvG9Ayo4nz7clxd+kFsHd6tqaj9L+qvBsR+zcR1J4F8VDnEzH7u4HhmfEPEaKWt
HbjP0L4AThJrw/kiymiL4t3juGsUgCzfkjlG/HmO9o6bnGzKuFPO3nbEt0khmkygm2Cz/WjNqJaJ
umqysMHoswPW2MYtnQZ9pL4QHpxPxAHsW5buO9/HnprUncA4BWkuyxDuVa1OEKM7rjfwyHDaBaN+
B0KzCswV75u+x2gxURGpSJxBfjo0itrkUTNqWfinYsBQKM0nYYAstBhMfvYOu+OP4o6+EbsQ/xbx
5taTkBjJUJNc1XKfV9KX4MRKO88Kas3JhPHmjEJCfcuMsPlS22l6bDr1qwWFMGLTYrUtZ2kdRyyK
5NRhP8gOvknap6valh6nafOfhpbFLszoNeZcM4ejLxUcnI8IdFt6AUb5eNF3NnYN6b+eJQa9oPCK
0fbPBnF8kpna4+HqKcUAtuXQq3FFvw3MiKrL0r95Mr39sVDiR3c18tNyF+5+H3N18IIqngKRwG5H
OBMi7flD14AUgqFuTqeuw9ZgvKxhOHikTxSenLSXCS2VAZIA4dOpZJLkztN4zPq5gUzKs4zaKUyh
NQ23+68H9WvAcPj95Kw5k1hYFUmKYmA0bNFqu/aD5qz/1p+/vjyMzMKhTtw1qlSPIuMXCpeygAmA
3j9VHStYkxv6NmL54j18mQR5pUhOVKIsmFF3eObrlXf2fhrmBWF1lCuDaRCi83ALWFJhHItggZ9N
j5Rawt9rPVOmXoUaNt6XbCtZEZJjhvEI001f3lOICs/tiBcLKz+Vs8/RI+IDBDY8v563PYCEup3s
w4tlZ1awSfWIf01vBOyn5czjRVFwmFpmv7Bhml7Hh8uqQvNzrCEYQHHlsyFNLHRBX8NMZXfumQZ9
Ob3hE2/zPKDGbdYaoq8AOBnKnuxNXaD1TX0v9RXtvO5M0tgl96yP1ECiAi5Y00REyXTuBOUYblr5
5Ui1M+aWIcBz3fuxy26sDK8GWAM9oUzszJOL0CUHw0d99l+ia7xQEjGRenJKacoAzxNDaYw4uCTE
etypYUm5BDxGf9ay6AMXcVqvtW/yjKgADeOdjPr8iSdpvL3SdplVIqALJr11+594viSzgxawl8cj
g15pnrhHGxr+OSg6lWW4VJO7vIZ8Ah5sAOPPaOOyCCnN4x0FtasoobDx1IgVpxSl/B63EnC5y6/j
dqBgsfIsZhTeLrbruEHJ0NDqcP0VBUwn8t5hHD6apoMyeBmSlYZv3fUwTnj3jqNYl6K3eEouYzou
Vr21lPsdF+rsyGQhbtbfFTCWAiuswkJvbKWzvB1tK29L/eCHvjJVWEUZgbOkw0v43n98YsSGN4ei
Hi3c12wmTBsLip/glSYToxr3uoEq1ygYetYTk1v6e9UxDS012kAGuFBBY2MKg2WKUe4jOVApcO9Q
YNUiPt8HmVduy0pRsvO5v72AmoNPHow0r6YrZKAxw1otWeSzwgDaOn0ISMHmJGf9FxsGV9yiMSIz
2oy2BCMTbXjCEsWY6P0DlqzSxI08UqYc/GnswYMPptfnADnhbVkWafY7VURxZ9KHc7Bw0if7ZSY+
9AUWKzBZRtfn1i3811s2P9es34GI8UgE8+I/xyD0pd9OlJcMWPF674SCV6Gh18tIOqjgZ8cLk4A3
64sT6ih5DIx4W1hs6t9aQiVMvL8ttcC/2qMPQNIhmIYalvJHl3zf3nMGdNQzaq+GyawPQD8MQgZ4
mhI1yFV75as+ZgOqMibOH0A7xfJ2aNOO2q/KPc/7sgwyndt9BcmFAXeRebe+OkqPBfObPG3af26h
xn2Oq4umJERlEo22O7u7H/z8mpbCASZ22EU+LDIpsW+YWYHNCj0DFAoiN8o8H4B9kKrCgVvp+cbN
JeFoZMds3qlwFKAfMLiBBfaNvxtoXYDL9FiEpZoNE305YbvB06vR3NvUBxrLAxlAX1WGiIjTAn/h
YAHoJ9DURLAI5i1QrNv0LfVuREQr6cRZ5ogqD+QBuiVICnMi/CYm2QLkQdjFXIABzEh8wI1LPG8d
DOW79pxjHrCaDw70jfjJpRF4V5vNuzoxBKwvHmOmb3D0YpJNmdI2Kl/AlmfnYIdG4ODD641Iohra
KzaahQxY2Hd5EMz+Ux+9bxPzKGmdqBhx5+5AXZhA2WaXixFYve2SKWrp9uF9ISmzD4G9OQbk+WyW
2/cqNBzdyBFhX5pFpdcP/jZ0XPTHxda9VvjJrw8PRFr9YkOX8fiA9Ezk1Mh8z2W+DiH0405jZE6w
dyfR42sSs1+ZAxJh0GvxQgBQUZrBBTRFKdJziQjjNnC/QNSaHi/Fe9C+eZNboAlOwK7P65NLOGW9
gW5cB2W3NiJ97JFxLPHUTnCF6gzntGxcnYwR2P13Cp3klVan0HwYpsWaS+kOeMqIpA0d/sDy0/gO
MVoFy/ewDOFSCHhS1O1mv4HsiSpR4wzbRi+dARrmUsdl9qM9ja02dTWs18GldAZtZQLCHH0rIE4L
4RKEsrGce4asKwIDaJvHL2lsyQxIE4uHJ7RswsxuZD8MHn3+/2wTsxNhZh/9R43bdZr5svhywxyA
4zQR+is6HwfTFj5ju+nPWzPy4Tvsf0plwvPdwYvxC1jISZcGc49A4gvzDDg8SOv4fAasMpRcuGLY
8CIR6PqHUwFmlY1ZceC7aJi6vCc5ggBDW0DHQOejyRVJMurblJLuv4v+p6hN1aEUCLkLAvzHnYBv
5crbq8K4RVfeSRMRwlXc/lXs/EAiG4v6YpHkcZ9ko/V3yxwqdfyuIhWy6XO+YyxgsMjMn0DyTW2J
sJapPs1HGGzoIJhyFVLtcJKJaIJH1EqA/yKlj2zOTc5rCMnFoMU6h+XNYZXEqImkY4wVpV6Eykvz
44kK5zHHJeDwt4KzhI7aCm6uJIUM8hkBVhU44GD+Nd/HJ8CsIgz88PC8b8Gs/U+k8QxLqMUPxRVQ
touNwD2jqdywpPwNwrpVWUP/iRspqHY4waIerOcSDXL3sCuFT8PV0XmODqqGQJ38BBd8TcPWssR8
g1Wd6omEAYtcQhjmRajKTK7Q/Y3eSzVRPPjSHdN8LtXqoV/OHN6iitWuQzTmnvmDMTokgWW7crRZ
TQFccNpH53OTYYjTNqhy5DwxW2Qk2Seshx57evPEK0D7i2qFoI8Zv98pUgU+7lZbenBBCywSElKH
FEshxRTc8YPJ5c++LhY+E5XDWyqlq9e8I6W91HoV/KIpt4Pjv5HIWU4m4kWYw9XwvSBVbneqN4Wp
CTjaj2iv1kQUiA/gXgxnAND8UBq6elTDv85ose9i0GSwiT8LhL0zDbG9NV8I4jxWAmayBdq4rGrM
RHL+9F8j4nLrVarxfM3ONPSWBfdwr9LxeYoMEJhOFG6N/LLL/o8bjmHNIaboUOAZRRo126GEAhZM
bXYRS5Q5NosjQh60DkJByWZ1cojpY5/aU+/96qrlnG+GKVHTGWF0XgXcG61PVL2VziPhj181/86K
nTpFu8qCQHZnpSwMrQfAtzvgCy/sm9C3t90Xje4d6brZj7ZrDwp8dMX3MlkRvIsEL3mARswisflb
9JqAfawGUNQK5OgWuZyUXOXTPuUqCMm1DI0BMLkFVuTxS0G7cJ4rGtE+954jQCWXI5+A4ixWoRkO
caYhc59PmdL2EX5SIL3xWWK3lg7vWEUTqPvX7/+Jy9UkAtaLJqZg4rI+yUcKDD0VsEl2bgRypKpM
kMU0a2KYL++D2ac5TsMZX+blzy3FOIV9ZlVTdwrSQGc7nCQNRfImBb9MVYdOLaKv2tuAjt3Wa0yl
sE8EAPslwwgodhfjMAwyvweNImmoPn+J3zXD3TxdPh2G9/nhKoN4MB4inlGXt6Gkmb1hUuiSzcw6
/o13NtSmD/1U+esrGcdAG98yfvKPecGomzWvK2vtpU2gQYpxurAPuTuIloTR8kx+a0tQ0VYQ54//
Ks1bewVCKW8IHZn12HtYg+M5wa4uyDgM0g1n4cc3k3ATh5brKw//kA/1i/R1abLTRgVhGYpwaHPK
NyODuUELLErgug6uRC97a0Gk+t9OKPLzi/pA44j+EK21C1oH2yoKk/PqLMzpJi7cETIhWne3Dmv0
DwmBxbfvcKT0t5Bw0620tZiWA+TtuIqCDWJpiKwHpV9eJTN+Zg6WFj6tfAg0ft7zPmjzkCZ+mg5T
Xj5tURRtIOb18rsolXKEJlOFYVNQ76yIOBf9cbsXCdOiYfVtZCW1Jn2M93+MKTmaGHYTdfnlSbXv
VxN0Bl2Z3NpDHcYIcIG9reJIYTPjBkTnr8e4ZnRDDv1ri6W6/htabU/d6+vb+g26oXcwVnjIHuku
1uuy9BRHl29ODkOrTIKEbdWXcxcwEp0HfKoyxUUQhgeVNdQmRwSnOysZpFkcUXojZuZuc7GSGSGd
tnvTPg5/OHmo+YbJjxMHWDP8p+VxNqJrAaZlOUVV1ZNT2kkkVS/HF4uPimIb8darYdxrAmf35hdL
AQhTxjV9ZcK2wiq2RcUieBFfEddA/4p6orqqH28/Ji16lM/1Bis26zJTtgQSP+PMqh6g8CKTI/DM
cCULw7dg1hSfJXx5fDl+ckvoFuznEsC9VHNyw342OXZREr44Qf0kxjDGbx9xRwCNOA0o/hMq34vG
4LIceEuDYmscX/V8DL8ifymJQjB5lM6tRykzpzDXE2c7JpaEt3IIjgemi8sd+4KUxekucvnkMnvc
vW8cYAgRVLYeCnhw2msxC8CQK6zrmOR7UA05f+3JdlnVg7RHgIuzSwA3i9eGRl37ZNAC8EQTuq6x
FsRN/4DjKncoU6Qne/OjOXKUETvO2VI2aQwI7Js6ToJZiQoMAqvuziU3GV25me+JJO7eP2XqNe3c
3ot+qAWRvQWBToAmHHASosjdu9HmuB2jaAqZuwLUEjbnbW/6F6b3DDw7Hk2sZID4Ub6F4mPiVDYq
gw6l6npk+KXAtozvoSyv6C6SS6+TmVIUvCmGdRfGUuUKcAOvIptGGP6MG/AXbJ7lz3wxSRva+Z7o
XOGpNfzDy6cNbRtqBfeJGlGiY93JbUAaEX/GTldMvICQhpzKWduq1GMid7FmDSunb/FLGGdwRuz3
r0xGXKmXdbPpWxxJoCKTrCHfwUNbM7CNIH0wfQnkJCXa2myaSaSP6ftnUUVZ5ti2duU/3lOYuUm+
UWhJ3yBOi1o/IBW8Jn5DJGUJf5y77n2FKpiWmXh4ru9ErajU+UROgthVmqHpDE2wq4VRoLrhszXX
QqR1vgienufl4xJMIAjTn5jIzyl5hEASr08FVjHcAjtENum+/Pt09WDKKJkLCGATjlIXGvxu1NXV
cnpezOEP3eE7RzwxAw7X+TiLwnrD1fxqawLGhKARxxxGYviUmrQHGNGTVFrnaRl/pP8ry9A8S5Cj
gHF0qdleJCz2r/f/1vbV3h+GTxyHWdjIYRPxo5EYyhk9ONa7KuQP3OHeHe3dwGXt8QjZF1CXy0PB
kHP/l9VS7ETH4qTlKPu3DsMXc/HqXdegRatzGJ1cVnlhvPvR+SxlTrtM4d6gjvAm+L6fdLFS26rj
IvgR+hhkAbKfqG+7exz7PAqbXRE3R8VA7N5QN7H3qR4GUza/Fh+5yr2Oa3j4YXuuMYg93Rp6xqVj
AS/rep7WLq4sw2LC9lsonGyHDMEIJ9YXCippY1ldGIXPR2bRdRF3Qk+w+yuijcLCWkXG+ScPaFuD
xSGItWdXvii0qtbU8ku6xRJp5StanTUUDC+9udLMl4AMgz0b0nDhzMbeKQeMWOD5Ba6SyH+2kksr
shfWUCE5z+8j8VtTUQdnEhKexmmdG2N2/hi6HPXFJ/ZD/12Uh5OmUlG3/n6KLmc8Vlz/wgmgAFQT
KbfG3NshZJkqi8YFwUKRsedPFgZP3LIrc6Rf0uBCY4GzW+MBZ0DfTMKSjOLdDgZN0FGJL+m01Vea
ncP9gBwIT7WD6RqBzrfDD/ya21ov1pnxSg5AzU5N78miA57q1ZfRq9zlYRRaMWRlAf+dT7mio9oN
2H76PQb/BPTHz2Pt4O6pkJUVAGECkguaKQ7/0cJvtpMtoDyHoMu4W+QklLKqflkkWDFmz1E+uCTd
IECEYgdrry36H3iuzy+HpLOmquZp2QthQlXxHqkHhHWFzUGBj7Aa8hSv2qIDfA6PTpzPY/35LlTM
Tqr0VUMFuOn8vZwDFEpP1gjlb2mYRAfcETSyh4FDRWHqf5t22zT7sn1IBG6cn7mPPr/C8Yu1nAcu
7daRX/nkyHBqcGjyHbJ5t//qwWY/kcUvZHRumX7A7txptmQTGKo+NiWnA3eku7uQj3SlI91HnLby
Rj21N5uUrO8DM25eoge9OD5Y1tbg4pk328U9Mx8r8fdNQKk19BNRbGRAj78uRJRGgijNSAKpfSyu
sDtjSz8V8ukMysvWNCbKdjyACrwO8WbaEl1KQXQa09+YiZ88VGZlfAjo43lDiZd4zNWln3IWb6Uz
rWXRU3V0c99haUSrfRYymIuJOiSMJvYgm/ezhesWJXTa7U2o/AgBC+R0QrqZIya2ts9KAv6STB6z
hfI5pxr3KB83VOYmGMMhLOHUwjNX7oNtFRPg/Dr/UoO1dzsY9yyZWTnZQlciEGyJNRT/QikEjpqF
nEZ86bzj06sMAZriFYLtYDh34PFSqKn9/NT4U0abeORQ/Gc8LTbsgep/ElFfQb44LRGTQ3uePLKo
LoE6MHzwUPTufjQPFagPIl5BTHbrJrYPGCTZnxKuWt8hv1849/X5/hVIeE+VWbEoFCWSEaRziUSt
HGggkWX9uKA7k15eBRyJ7RP+7/sR3HvbeyygUbattRHot+Mllf1J/TkCewaCOlL9sejxbG5MQbOB
hsPuSP7MI+9MCAxY/iFiyyWK+2FMjDCQ6ohmp8vH0LKKJExrCJVFhbbmC5vAiK0m9FjpAU65diGO
7y6lmghOc4dMeysOs3dxqVgmKCG5jwvs4qlPrYSNO1Z9pmxjdYMnL4t7UhJibhM8bDxXlB8NHHGg
KoTIAUa+eUDpBZrC6t20yNmED9+/Bd/myp0viXqz9QOndI1Ty0lsZf+WBuBv7ZRZUCUebbmDcdYn
dYwItLDtG7DBklg/iuEAARwcdms5XSEjzToP1P+GoJhCZiaRezyrnOjIISwjGHLsYjSY/X18B1CI
kf7wXNfSYlN5ApMh26Wk5Nhx9HTrv6l3pn4CAHQQoEt5ZLZasjt3DddaHQhLLbpcEJeuldAOJ1r4
wy5a5tXarngVm1zWnCR9E0zWemAamkj7sj2rH3iAZSp//9b9w6ipa+4uRppTPS35W5qp0Bx6awtI
haItcE++x4/e/53CkGF87wJbfMVegMMPDc+qwMRvr4NHgMrTzqSk+Cg534khqA4UtlSyddCWeQ8v
BvPFHFEs8Z26MVdUMvck7xCgOjT0JixmbRP+urTF835f+ypPyluJmRtfrsfaYrXSo6/PyQfHIJ6r
lzL6pxkJs/VNE7VvTxGp69riUS6xQqUnloZeh2wRjuD67kcc4t5pUPK3Oej9kXXSKAHp5j0j5wU8
077WQJt6Y7/euhNxhlvIP6GXs5iTDpn9V8KgVYQsb8iJeGRbMQMzMKP0kcHYP+z4LzOIlBaNDyI1
5gXWLGGYDgygMXAol7AYxqYTO0TAHy3ak9rxziXvhJd3PbwRBwRecNI9DzFUxCCQkuwdJB6JHVwO
VAE6o+L6FUppsN8F46eKrgm0EQR41nNKJ24xmn1B3T/tVWgqnHJNQPlV1/eai+loatguzl1zV69W
bA23/3oG+nce1SEPhUy8awCWhH6LLCCM+WJd+HFG9Fq9qpsPIQvJ2NYUvkmQwru8Ct3Mc/WQJdo3
9LLKo8gJ/s2NvjnTYDCHjrbqMzdQ2KIBTYee+tJSyj1xS5MhHjTe1Cb/dls9TdCy/KfaLUypw08N
xxLocv/KL7BhyCTfFJVEIbMVhGbcmuuDQc12SSK2sMY4Q1DMWExP8yAlBsB+Kc5+VC+QYiQ3B35I
fKqgrurOJWh757+08l19WzS4IpmYQDdZo5h9WM0op2N6sRYdjpHfLnj8FHyYRiCdUw0+osmpP0TC
QZDs8sJC41x5Vp/bW4hq39akg/hVQKDchgZOmjWxaGr4atop+76uznGbHjJL9/ArYtEE8hBMgqQH
Hpvt9zomoXFXHHidGvr0PqeZ68hz8ckDloaRZkTdxcyCawMAOYmAneFQkj5PZxrTk0WAFhz0pSL1
1bgLDa3hDxL96xyrHxMOtFVwHVQlIKwAPBLN0GZDu8ppdoLsfPzSU08/ZncLYiuM76hUFQPQrG6G
Kw42dqzr1NP8o9fItnSwtUabiEmB3ZhfPYqod0KEkPGDUBmFpPwMfOFIQtDFLn0uxqIW4CgzzYzt
BqsjsDTeS3LD56KHjZyYIEca/IDqozJhRMaar4rD4Gou85IZV5aDIsJJR6NEPa2JFhOgQPiqrWSW
mOvnms2gQbLpGybgg8yYNaeoUXeNAIi+NYWEhXs5cUQCvlySTiRv0J+BnB2AEt7oGZDRJlGJ6YML
knPWKUerBHfATsXRcViqQ07B7GO0xjflphSW/UG2BBY6peq25u88phkbkdGd9Y7i5ef7JbYfMvf2
yFj07OAMaI528Gm632epeUgnJs6+by7uGL7Y694Bm5lgH+74yBpZ2TqdcrxusZVoJuG/gCcz3c/L
Di0ORA62y4BRhaI6vuiT75wxWA1pontYFJv/8JwH7WtvXPvsY4ZtJll8+AbrqWJIHfv3A0KtFlIx
VduoLId2ArMpTRE0G3j8633V+bdW1c+k/rFmNYXgYhcfLblRPPeIL8mIp+vSJaO5t+faWKxKl3x/
YMeD5+1+fMHGuN2z1c78gAnbT2WzBJTR62Bf8A2KtL4eV2SB64YwcNQ3UB3aW1adqhoC2WmclUnL
530Kv3VUu5OGfAFgjv1zirqD9PaxoEcFkeqSrNncP+wqBrYaq2QTlEY46/NOxUr4J9taEPjFvqJi
LUfMzuj1wGR3wUaK4ur7FZdHH4CT+1k9G9YmceRD1rV4/ZdM95NsbgrkU7tA6gtNShoHaVC9O0PM
ZiAzkwUavw//1Zyux1aWl366iSB50XoacN7a8MrA40MEHX8ceJ86FDFn4wkHTxtDKTRnQum5ogZZ
U72gHcz9chjxPJR1ccK44vQwh/c7K858nWFAcXVVADhzhtAvVDWHx+9VZe900nNIAndUYwh0d9Vh
b/ZXeQVoAbk1dtnyNXNBkQ+je7s8Tz3QklEpn6+Z9LqC7pBJYFdGRHKnLWtovJgEXiYwlw/iD5/V
w/SkVIMp5mIbJBxOVMA71LOBpzG4vxBTd6KsAKqMVu4m4aP9EVebpa6qFXB9ZCjIzknOH0Mk0Kf0
Znh5JTNHRfGQPES2OV9WR4feW+/xFasohy8YGTPa7ZephRQGNFnrtzqbVAEYebnsGMmtQPGah4B+
a7osmVGD2A3KWZxxd3bFdeaEa5QNjJ4W2X6lmj2o9iewHVmXGt7nzbbdNm1rbeGahS9Yqt/R4dMK
4YMv1Lw3hC0RCGsY5j5OlVAi6yGLnEIiuIctJijrPnJAe4ya8JVaKYKv1eX6XlCUGVO2tir3c5nn
a6AVlGpJ5U0yKJiBkCbyqd9+rIq/ItHNzl+nJY+QWJIdbD0unz8AmGhGL9CjU2Wl0KqTn3mNr5Kg
/ysFDAeyGqL1bF9amFRAjUZ4qrH/3fc1/iVnT+OYgUQnswNe2bbHf5bMa9kLGdesir1jdWUaFan9
lM7QmSW8/6fmMxAfuaWDwrEQZuGA8VfONT/MFgJnxImuJmZuy2Bjrr5XBoXcx2+2K7GGdaAM2uJJ
I1uj0TFtszXixgZAUZfpJKzMfBRScwasHz4VEaZMTh98qeu831wcza7M9e9cAtscg16cW1O1GbpW
O0n9YXeOd8xPWfuAJiXVOIn0pGg6Ya8JMjmJaLHBEpsMh2vFiWKGLXphnuxt7OC/Tx9HTGxZW4KX
m90lGgVJl1txHo5xBg1wdxBv2tJktU3x/LyFywidszBzoPhQKIH9p7Up1OM9IXtMb653M75i8hxg
urQ79YdJOWhOy+73CCWF5juzfLZ0ovxxBV0zN4Sldtpfm+LWukX2ljcSpyrpI7+emvQNyevXQozd
aiREOCRcXQozBJGe+gZ5uZduBg89hN7Z7OhNxEWKkvCL2d3ZFyys11Tog+0mJLAqDHhmMrMzEG6+
Kv2Hyi3fOdPjOxKaUPvrC8I3bXBXJbleGp0/5xGXX7zyyWLeyzFksYPnT6UUEXOq44adN5n8klV+
clmERyR4lAm7QL9iZplSNVxSax01yx5hupKgV6LOI7RuE+uvaO+jg8LXDqP7nYt1eX0hwCYtTU6q
SultotdVHNS5BZQ0vFR4xF/52JNbGsg242MqQ88Nfy4wlgnpVC0j2iYPHbK623xTf1ooXtPBoBoe
MhzhElgurhESQvAM4zn09YndAEnZB0pFxtZ4/u3z3bkerNXkbVFxWFTjd8dKuH8VZkxD9s9EnLRg
nnny8rsl3kHF23TV9YlfOFyl5VxHbeTb2s083d0qnF0E9ogqP0ExQ3pjF0aPcVoX58hLEoz9m6h5
FIZ6AyzVvnYwrX/RB4Ca1RacVwHwvDnIVsc4sXeQ748IAObqa/hw/A1V4XVEuXLuwZ+t7rQ2nMB6
/hJ3CCqWU4+QH79q6DgU9i4KJQF/0dgOoPTX0hOt2kxQb4NkrOOOrGZXr78gBotAH5+YjCbL1/m/
XEJC3JTbdnuf58IcwDWCTgkCrVAwJ2zMZSrM1kHkYCxZHvrqSsKQwU/cFd8vcxDyGPvn2WnCwKg9
84EcWRsQtNCEfbUaat+yxNMajydhjaCLoDm4zMP3RV40C2wtLVr1UVXIJ4CU5ZgLSR3zT+iE4a2o
t+zjwh2mMUUKCsLkhSgCVTECbUhidS2kNgUeS54VbC4YSYO7gJqpEr3guWsLEnq7wcm50ZG9ZPEp
/PifvmwobWS6kzmSbgTb/85gsRefMRfw44q3a6Ps1OW1t3wGtlNNmcipvkGsorJVtCzTUh5vAQU3
lZ0gMH7Xyi/cTHTV+3wvivRwnf+jGbkDLBhQK1Uy0yBzAnY3yIoLOXdRMXnf49IW4dhBlAZYDzWh
0kK3J4OELsu5UZLJY8n2fPdEiOb0zOqUuwLs7bEaTUwPR2LritxthgS1liRQA88PF0zqk2V3JJdK
jxnGwSvCJ3ihj9wrXZzB47xsuZ1TmjegTFGn3J3cROXWEkhU2IOJE9VaKyRsB3MPdiw1nZlzzMvD
EfjdblhVq7wjHJT6xe4IJjdb7FyXVSYwOIgHts1NIQvi3HI9jelqp7jtGHZoR9/ZOjZUSOTcRO0O
HQANSxZLleWKz9rHAsMWPbLCZOcm3mz/q/ELITpVUBRnoZJi3I5MbUJnJ1Q/eGJDxKpa8xwf/O0X
Jd7EcKLSc/cIbsZdhAr4BNsQ0QnI7MIVuD/nqXwnjkf2m2slQ/INNrMDwjsBvglfcDJPon89LUKM
uNtuBoIrP9IFrshpxA3yamqnGk301hKamVAaU+t3qpXel7L0xCIr5whi5xAGU1rXaLoOMI0KRyUb
G5dWywrxrdwyAiAMCn3CPSQs7eluEHlCUDpfZ+uHW/3/S2WmfEOPcWKmQUnNpLnDVGqPMF3tqGVT
20Wtg1oz0N8bDE9IrSvJ5UlGLpVpmC4Ggg4ATINPFs0Z4rpNLslgDrfk8DPEHsYmFBXcsO1DpebP
616ddpOFinf9ts9wJ6gR9Ok7bJJen8T/xyIumq0iH0X4nY557uei94NtTlHbrVW5pvqfsZfI5rVP
JsmDfwpqLvBU8S6qpd6wWNxddqAZasl8JI06V2w5LYcW/h7wWC5P49rfOUIJ25oy0D0CCThF3iyu
512dr/hrDXnTAic7HKqayJjvLv0vszbmJ0ulFAzSwJPgcQFbMEkNneObSRkEXFuaNBHgQFsoSuyx
rpS/+pcHBA9cKsWH+E096pAm31lqom9eumXqvbZz+Lm9DGtB5mSx7xXE5Taj583s0UTbMzIyn4jw
ZyDRrCKt03fxllfVe8T4/7IdMi6VECrWnJ3RH5D8mtrChyl+aMR9eu/k6q2jy6Q/mvlafstKCc5V
qzSOeCqANE/jiOEJmyWABaHDt1x6B9ZDUf23cdnnJomqnt4YsI6OOKi6zRP0Xku+WDuhADasKovW
UH1Tbvd2v0NkPZLTzYCZqKm/6u4AoQs8zM3sU+4E4aa+rQGlgBAJ8gn6tLfpmB+uSMi2p4hV1mz1
TmTv1DD20lKWG425bo4BrspwVxWSHcj9Ca9WI67dEPRig4+8H+p9JTG40XZ12MT4fB3DEJEXkpjt
HfMGsCgCKcJ/Zzy/puIyDvGu774C7TcB9o3mEA8cyU3vGm2UV4QfyqRIuURzrFYmvuxDlBUG5ZHi
5xHl5txA/Iok5nGQ2j+u5Ot3DGRMO0kgWCaAerAWzzNIQ4BoTvj2eIepicj82Ul69YQpgv+f4H8v
9tPOouGhOVkRNXDkqUqV34XkIDr699JhB6EcRVlyKOJ3w19GvmfL+xZBuyaqodt/6IjgsdPmQzSI
+92d5EbORIzhtf4FwABV4zA1EUlA/nalOn2WF7EtB2C8G29PiOsEFSJGjGIfFMm1j0+u+hS4Mir8
zHuy1ffjc9w97V/Rfjlm4ZY+QYHk8IWwOyn1jbqGCXWym/bfO9SjfTFC9uBKZTHVB3/xdAn0BJvN
Rf2+W+M3ZRTXpQ35/Et05ZNb1hQrvE5Q+DRhFZMfIgXuJlEv34KPCWFun0lUN4CsYAspl3sqZA3O
Y5x/gIkKIMcBUuYquUjzYsEFiiC3JmLtY94VDpUMWck6rIDSlcw5DcbvNVqCvAU15ccSzyziCviY
ScijlYJOM4pz/mhJwgstGPd6L+nbra89+KfxbzgVah1MKJzzL+/PZvG0RBRrXxhi+mVV30qrepcG
lfjqFNeZMNBdvtEaWW16rMxidCRX2FfX0UaXRGHIarVDqNjVnqrk4UnF9HQEEvrv2VhmBJTk2u8V
WvvA+apr5xIxmtP3XPy8hQy4NcFnvFO7EWi16RV0hIjVg7NyLU2MxVDw1Gi7WPhJrLoYT89Bktwe
lYFzORqrp5G6SCzoS/KWuWkt8sIo3K2q8uwX7T2DGRaSSiCViLvD/F+sOUcAPRRddLoWY2QH6ZNa
4igThgkHfL+Wo7dDBwFKuuu5UsvsrouUye2uIaRlgfis2sIUdfiMLEi5u8sbUsbIkxinlRaSvVit
qRDjq8ibXq1d/ccQ7FLv1IvGNn2U5J2Bbqbschwoj40A5weX9L+5Mt7IL5nwkfVfK+jLLIahhnhw
Q9Bq1cds6UsOPtPzu7PblWfZUrEWWKfSK+oU6rVVtSfwnb+CTapUHdiPLrX7n0EU3TPfa54GqyWU
u5pBeUtyNC4niLMz7acLrZTHJf4AGu532wTBKUpM3hoX1Jq83BbXAScBMxEPrq9dAOfRyT01Ce+H
TyWUP2YIEz93kiV5XH9ojYi+3TTIhXWDRlRUxRhqhcnJOht8oAI/6Ile9nPswPtXB65R0BwO1JuK
vcoIPIbgCLjN9u0IF7LeEPy1cX4DoJYeN2BdycZ1zGv106ZOt32ddbC0FYo15JIfJQR76gPybc+l
2E+iuMsUzLHBIr1VFsI6PFueeGDAKq8aq8lfHUip3Sl1llY8e8O+IWyy6QLRC7ypFa1cNLCSd1eh
2PRnSmu+qeIkIrOCCev56IF6quykcCctWpofhHAaiQLGo0r77WC0YKw20sPrp8nQcQKULrWboZQZ
eP2+UHOn/3tU3h4d0C1ANVdQRdhDMdukh6TqrVraLtvNlkzz+j3IToE0j0tNB8GyqhnT1BR8Fzx3
c7AZ7jqPjLZu/R/MP1VGxRyCYbtv45oV2fzTECXCauks9eh0SbGdl1Zi4OuQXCB0I8ZQOwnV5EX4
XwGryc0RfHH6XOSltOwyj49uIxK9BzrLI0JOTBDfHYTTkF8hJ9oIoAZRlDQdrfO+I5P1f0hzm/6B
oUmkkFMfrH1nKbyFy3lTaoz/GbAhl8m8KR9mr78ENJGZ9Q+6OYSIKuoxM4n34H1lPiqqdoY2P+0a
NVPCqItN9n65PNi9RCWNAZhXT1Q5rTKSJlhRnXu2pgYGXEtbOxpTuEfakN42xuEnZtJoQHLfhwDO
QoAhu7QjIXAnf0oGm2kujXZPHxCmOslkeY/d8bi7t+aNutbb0dUeu4nqjR3XgIdyehaDvYageg/R
8J3ayUexVvfcOUWrURQdaB5bq1GH8p0ph6hjwBUm9W7WFUcGpCizCPTZPOtrpHcLpUOzUnaCp6PB
PSaGfwu93vHCAlwpOZwd8PviQR3jP5Wp0A9tHVDqa9tET373B3bcjh3pL0+xH3AZaj1vwMNSz6Xf
UtlTjWPvN/Etda3fSh3Nq3zn6pDDMqhiTD9Z3thGonOGA94YyopEDctRbcR1IWU8o4Y4PZUMRhAx
j22OpfSivTwhhmWO43FTlNtYN34r0IPmD04BRi4XeNCwVJHtVNj9kI3z2qIL10WA93ZYCk7Li4Z7
8OEJkFXpYILVr4v9gC98172MFLLSAxMkVwUMo1a0R1Tw/mrZOJKM4UYan26x98hRW9TRKlJwqA49
BIsURxSEqN6eGCrnHjlDyM6/WPHsMEjCUi7iQEcDfjx93QqKPTG4eZD6qj8w4X/292df1YCFIW/Z
TO1EUI0lPsDu9w72EU8BvXt12JVZifDSIlIxbrWi/n4pRJLRBhSD0hBRuALpVZArWdU0tV1nknBi
679AXoYcGSbVeyO6TckLSp4muawVltX2h2dPPdxnYLCyUMa/X/eTUFcO0yyNzDYopLrS0G7t/Rw1
sHHLUc6CoQsMTJi1SfXMRqO1nFCzWA6g+7hwr3F5dsWklNJvf4NQ9oVkNmYcxnmLB/Q9AOQCPz85
ddya9tPg8I1ZD3NsBBducEHHeYEKo4b3txh7EmFS1pzCu4hlZpiUL1t8WAlCKz2HNuWGBmlIib89
6IOBUTv5VlhvkO7nYZj13QYz1NrHsNalNbXWdTpMqdOVhbqKOUPD0S/c4IJhD2hz+MEU3nCZCD59
JjnpSySV9MYoog8vS7e/TaEfct3y5jYGNlO5ZJidserEEGaxRA3rOPBga2lrzlv75wpRO3X3muiY
VCifRaRvGxWBVAc6UQo/QN/NgY1ndXptX/8MH0vtoQDcfCu0T8OsGfXCrQxylsD2aw9W10BauRqz
Yimx0vXxXshZv6FtKLLEqYHZC0pjf4u5gN0tZOAcOXlVz5SceLRGsSGg8oa0994uqGJBSsIdFX+C
LDe0R4nHMfYou4Jkpoi4GAeNjien/7CWnhD9F4Ma0O8v8F9hcLrqQ5Jsg/AsFfzzwOGtXkBO2LQX
KPCb8UJLMu3Xu5sq4rSdVCYO0b778yuOaj6NbQ7qHLhAKGqXWDdXcsPhdT93iQNxTjVmo1dRL6jD
95H782fIBI6325Wwn+f7EFmFjoSVfqO5kbNJBxbhUxwvV4LQENN0Wg+DUhZXbQauLaygmLklGzb4
6++jR95qQJN6eGQtGyZshr8XfoIYTdz+pdLScwggC+W7PM1xZPaW7LKSiGaqmkzqCUa3vRuPMyfa
75+55njqL93P+5wnUgbLZ7FYpn07njwKcA/I7XNUzGMD4Fg8CFuIo99fLu5Tkvr0p0v9sZhUWwxC
BRVAUYJ+xcvThekJXHPgsjjxHU0PIThAayFFH7DyWXoCPXuFgOt34u4eE14VOCDzHrIcmmRkUEAe
8UP0NCHELvhkc+F3cZSMDXkw16w3Gt08nir4M1Zosw85xtcQTRqo7o7xGA42YxoOP9t7YsRi5FzM
SL5SjJKnHTQBmvsd2951e4z7pJJHyGOqxf1Sjy5sMcTCdL+Xx1KS/n59NHISdjS14QZJLAumxnm9
8B7F4WltVx6O/J2T8I87UXJBU8wVxqPc51iYYXxijSc1ugFgEd3jjzq7cbdaj4g/cBE58ubxVA8B
szVMSUuWfT4M4f84/pf5VLHLJt7mnirE/Btedt7lfFwP7pU7mGqGhWejippEc/gkBVJ7ZiGCrsER
kqZaCJ5gQorQAzdF9NuR6Gb3QnoeXH63nQuVRhj/fJWsDo303VqeSph+Qy5AO9qLp188Z7PAcuQn
T6oXy2WMQldGcSDU7gr3rokctLMFfZf/pU4SzmOUWqMh+2SBJLsJy35sCzupq98mv3cbOZgFh2df
+TeK7QC+Sa2d1VnITaYxOY8x65H1diQyD1MF0guMgfL6odnwG1SnmulW5bQxBtSNjJw+8f5Jt7B6
0pP9FNP0e3AD2/0ROjCz7uMxyL05RYggwBu1ylQM1CnDdptcmyh1I+HNXumWbVaBIJe4RFKPja/S
Tb4hTiRIfobq0CZyQfoNwL29G0sli9z9T2Rqoq6EDobe49S8GA178TYEI0ZIqhERZYC9hBQRnaVk
M+NDrfGAJuq8k8U8oIPCQKhBH7tEMMdROBhdm8C6CMoNzO1g+YOvC5tz/AZYIeK6uxQ1qW9l5Cr8
uvRJN7yL0LFUpAALKO2PeB6xVWpHfGlkrHpSUbfI5y9fB+FzOySDOxS3nZZhv6GKyglQVWuovp9/
yP0bW3OIDlQ1DqoWL19dsDKyRWbLQJbYt9t81h1ylfysyARU5mdyYBg3SIEwusM/wKy3m5TpLmjj
/O+zgo97T9qmBrE4Tt6gPLXoD94SgmVmFmu/4keiJuS9OMYZcsJTrKuXhYfUEVlDnSvE/061t7zV
feQTFLXun1V7TpgMDcnPuYo7JoEAU8B/RiBCI/qkJ7VTyM8QnJqi8RdjqBQp5opdejn0mxTxvXl6
I4rljVvhDi7Gc0xdB32qIfy3YND6P8Tb45wQXOzxfJCD0NfnxRI7XB04HlpQ5MrvWzlWa8SFW8EX
resRgXOqBihsOMmMgwUMK9bcZtbG9Ur0UJnGujSiP1Z6JCragpJfy8/Ffz6ahkuXE/Q8Nmk37VJT
/FbWR5RZnrLdLoco4euF4cO8OMFaf8As9idrGOCY9UEWOX4z35iUbw2jaQKW7mMW17I7RZOPakfk
2YFQX9U1TvgsD0IXQV/EJ5f9VjNwNdZSUx3CVSgIOZk7l/FBzQKhwznkFSpPMA+6Okz+pGhHKiDB
Z3xL5oquzESip8Bb5GtPyC3BSxa1BkHOT9nh04B3hJ/f1QGRQvVOYg1iDavhUJKNppPyjCVy+7yg
gdk/xO/aaHx+QzABiJyBYMt4FJXVUzyKXMYMBDoSxgkp46CSLVKQMZx2KPFA8kBcE9mi+vyX6qHm
Nn+QjiozZZpr5pmg3tTAm4pKKdW5gVupuD7UZ+QyO1phrZNi7YgTTsisG1QqxMvmE0M1ia0tz8v5
/sZxWhps+RCUPBijlV2HcG2z5hM5jay2pagHKykiDdZpdADOdHh6z8o5ccQfMUbKZzlnabEMIJkD
eDJUNJtPAXEQN73Wzh70LXNN9wjlHrgew8L7BE/+4/7F6xGRp3HwR89jWdddoMl6pbP2GXHQ6GF2
AhKrXDmInk/2kWWOsm3+EFV5dK5OZEpMDq2VZOeDpasQlgoRR7jQGv1dEOP377R+xt4G+YutYoUH
PTAaNgDpf64rUD+H2McGHLQhgfgYahBt54UXxqDzXkJCBVrAaJEdi2VEn54auqi/0v6rWkDKkyiJ
4AnWJlj2J7RHyl0ue6MUJZZcJ9c/SX4R+kK8FYOhi78F/Dng+dEc4CXKO95fF+5dEF74dTJFQoau
GxJTphL411M2Nfshz2emgHNEghlR0Fqlnz7yqh7vKQjDE/jX3zSn1S0spc1wXmmfrlMK+ScCH5uw
LrI3rcVA/ZcBZ8HqqD3166tOXhG5tTGt/BYquVUO4RW7ihwMuW/jKPKgcHw6ZUpQmj1gZ6CkAF+N
DfZn3+I0vsBVEdN3MuNhNucGgiqkbCPeyEyUQmXsjy8KDc5L6GzyCW9SXPxmQf1fw1T4Q7/z96eR
WS5WVOK6051zFLaJ3VqGPIcdWZx1dF0Jr89BPVBe7+cXhjqdDEtgON1WSsXPr/KcECuNIDp4Z6wG
x3fJYo/P0H8BkMv8Mt/E+Xt3JAftfvFAMfY5h1J8bIJ93p+n05EavLArhan2ZYIVegb/YDGpsV+b
MEqlH5vW14zOGElH66GTX7wrghqwxBBfCD4IrcelU6tYZhWijNfY5ubqffe5ZR8LkTYJ9S8DKRN4
n4QTScg/TTWjI91g2uIJG6Di3dP29am+FJldLi1Acd0bAAQkyJPE1Os7689Ljr+bKo784pWfmQmu
arl5ZpLbXufCQQdNZ4uHu2oVvm/1Isz067dvju7cFUhsvtkZkMqaXdFhXbgKL5u80kLPx6o/mbHR
6oulKRGpe5ZJb4h3MPDxWiY+gr3yEndrwBK6ALNATSqO2HXz3D/jympSuVMjzrHxvvzlQr5l3Lq7
Jx/3VP8G4IbyW7f37Tg1cS0N11FqI0/fDPagj785T07TpA7RDNL1h3w4rwnLQkPPTVpszL5YV86+
xHJg/nod5ZyZbEE6JY0u9peap+3DQbjXY+buuNk8zDfFILFgZnTEUt3C+alqLo49uk0tF/MzXRb7
UFFyqWq9nxBTvO6JMADkpYI17bfANRHrDPv5pJs2X7OrE3+oVDohlvvppj6BFtwsigHlV8YAW1+q
lQZZRejpm6CcCizUriONe476ddj98AzeI7W+WtxvtSVnaVKZfQC+wlXrS8KT01N0KFVtap53Bd2A
NyZ0V2OR2ZmUB47It1mGc0Ea3nrSF8FCiaaXu83WYZSRl9OgsoO0aNm2dJKVMnwp2flG2KlHVTn6
V/wDxp4oK095oOjHgjD215dyV/v77U69PxoclUEv+dZ6zZsvAU/teHctmyMrvhEVyMUmsxrBEG5H
FeGsWdBD17+JddF60vdNpdBLGFwvDDv1rlV47QFDnEJ/QQwJFRjW8L+aXkaTWl7dheODtSkeI5+k
t5hijN25nKgDFRO/FlmhXFmTeFSQIgpYKvLo06+qrnipPmz1CBi3in80fLvmL/7MEShck5CDaAoJ
QD4A9OH5x/QEIFC750XIPFDXfj81spCZsey94TXwVL5jkgLyh8FuPHeMsFfW2LUMysoDgwmaPMBx
FBOLyAuhn3otHkd/GEMByCMVkNHb/k40s4NE/uQaUayNRxUZQ7E5xapesJXFuobirV4skGqfLKtn
pGvJywe3ynRGFAm9DODKGxzakbcG2N250kG/DFwxxyM7ucjShoSm27hs5D7P6nFtpPWqVaP9fWoY
cKOsnDkkBKfQ5Idmd4mDyNcbuCQugv2tmH0jNePZuxtUUfm5YrFG97fSCZgh5M9YGANr6eIZkWYN
MqF0dkfFGGekD58iF41lKVANb+4tBafeAlmLe+rw0QX30QW8xRUYZd+J83BPeevLoLg4uha9b10W
HYpl6dR1g8gxuL+vQUhd3/tTCMiMqghV6ScdLrXMnPtpGPSZkD/ot5sDYe7Px0Wkl/fPUPfA5Kqy
e6QYTQ4bLtV/IYHUb7yt1/N6DKrlv9tEMXPN9mrYaEj92TC60xRC8ZKFw4kYswDBjGIlwzLmLAEe
+K7mumZ6OLQKAImKbEbMKJtuFaY5c9o0BuqesOWiE6o0pqaQOf3j5rm516U+8PyAi8tKtRt+UUal
YbnV1n8ol99thv1Q6L0S/Chp0ikM05r0tQdoCBVzSQ4p2DrVYesrV9+HiL8jKfC3twvkqYIc3Ytc
8rVnZLMZLMTCHQzB5eptYu/rPQE5DjczDhgqqaJ3wlbAkXIhoxQOXBMBwn6pmdgGXBX2uFJgIXwq
cjDJmIGUo4rwiESA868Eqdiu9cVlQ4d4uxsH4BhUiUri0ddx8BVwuNAWmB3vCH+wLk4R4lMQaIQT
j8umGnsnUZrn8R9h351wNtlny9CKrvFa0ye23EKuEWjnXX81QI4up1lbQgf/mqJhuI6+I8pW6jKK
s4EOCDonEWGODtLYcB1m3/DiE9tATqQI1YYD1w7TxNw3XXBv3dC1FZ3f7tKZcgZq5xI6PJ83gCgt
Z7th87jjbKvkx6lfHu6zFeOBfafUoLafccS0jvBHopbI/UwAqj9U/7jA+xivhzh2Gsl1aSI9+/Fn
H28+h5miFsgOsEHUVZFFEWNJ4Qko0zKtgZID3RVIuZYnzTbX+nysO3Hubc6PYBrElVZbXYyw3Zo4
PiHYtfa5spafupXRZ5yMi6GJtjYmUoHd50/EYpcMtUx66QfJQNTOjLcDT8aIOoFHcpB3mAqjW+Pn
USvxS9TBcW+LDDQ8UloC0lql4q8OTPMfRKtlL5lpt2zRIw8I0LVq7VSfje+CQlliQJNkp1xsnd8M
mNb/ByVvHXcSIbrnOxL2KA3yZr07aHUSs/Or+I2DozUBl1jEZ2hlnGog01JEI7VWIzmQPxrvAB8m
xqDbnAKkoGvGVKlLJRJ3qOuvS6Iz8hG0Osgtx9tP4Qw1jC6KpPgrX1INZlcFC/D5zmEtfU9c7vyV
OrThzKQksgZ7L5ylh7OgU9ipTBRLUPmOkHaO4fBZ7s0HC3VBFQuR3iE1gcbfvMySuccHdMdZMlHF
Ud5SUlIHw8iUBjj+GAXYegLl10bKkRlvLZcNVtYgEmCQ6ZUg7XDG2zt77AWBunwk4Rlz95/qzg3d
/HboiZApF16ZXlRs95tGZdDYBiXXKDZPCjn6zV3XPU+hsWQqyMGQ4VJnqUvoIgFbfDCLGNvOMzcL
WSUajhjTmd1M9lFbRBHDzAlOh73sJmFV3PZq8s0Omrm8TIVFEFTVaj0rzdNB+27TPIpKZM3M9Ic+
kQJVvASKwnBdZFjo1hvw+mqbNjFcE1DYJDdsVlhV72YH+MG86VaLXhmQHq+Lm2GT8+ib9PjPhSkE
l8wVYh4N1NrR1IwYioU7sOZGqs0kJxY+jdHf7Gl4Ch+JwjffKIiywGKcYJ2DcxvFQERewPK8gVrG
uwueSQJU4WYodtTllsDRE2BUbH38Dv2GmEC6d60FWsny6hIVBb/51m+k8iTtJpPIjDJ00qruHPxg
8dF1qhrn00t656dWEQ9a7Z7akK5FeZv7QXWmsLBLg4oa39XyTDDI+vOXbi/4O5Lk9xpV8dOoE8Sv
Nkk4euzwlVkI3KcEmcOw3HBP7V0Kiyi+IEZVbscjeDK1ZUCE21hD0BA1nFB8J0XqjN7wPA2vnXKG
Ju6Ypm3J63kwXl2TkwrVrlyEMhGwjKAJmqfQh2Tzdw698ydoj5QDfBJtbvNQvVxbFdQdrHwcL5ol
yMith4HFHIXHsHcUe0QXWuWJOiW7j+TJ1IP6j9inZ0hS9f3qlapsAbb5Xy+iUoPoWeiGztAHJxQp
tpr2vejPIOeAV/gQg9qqjdAAld5F7XG+J56gfNY/XseC1FfLeCAZWDSdy4aEdg/+hytgzakyn/ip
OjZ49Kiyezx4e+z2LJWKmFmQ/7u6qW0OCbldHBNH3Russ8R/kc1LXcE7ZZ5NSCR7g3pYZVOHKNgD
rkJ8eDkWEA4TA8/dj7FQnJkFvVnB/CdObyM9LzKT3qJTAYib+XQpISogJwDcytPHML7c1rYptK2k
lbmLksaSrN0p3rJQYGrOEmCS1mxLPtmqXCNGh3wfYOsYCrP9jlDYYdJ7wsjzcAzXWFEIdTkCpvOl
MIglO3ZrmcftWcINBhxLulr86DVe+8Huz7JMBaAsaH52/gvnetp6/tQUHkN3B0ixXNkf3NFzBPOG
glEkXcMKg5SoMEksbp6xbX5VyhwBm25ZJtdAywZoRB2ZKUHB8TMm8gsMNM86V5It86a4iQywHQz0
tPRx7AUpQHS4+M/7fJ4UeASEGzFBa6IzO2bGiKGkSBH90sIGDc9OmwT2uqctfpcEWcNgrYUPeO7w
aMTyZ8wyKX9mjxAZZwqIQlNuOjZLmvWIEBlZmKMS+6QTCzHJMB337j7L9YPeBRW0oL2F+PeAWsS9
CDGPRVHucVPdGbxqh3E4cWL6ashxkC/W0NvkY9LoAMDOMT9te4Am7ShKLpifOBPzCTpZEdEccORM
2npj4NAIDmWJBn3nWjoqLsTtn/hoLNjPbZzmdlBc629NZaFQiF5oyWQeqRUCHFubPze3W0Wams9W
KtzHw+nPwcWG96xA2qj285A/eHlpsfzPirzijSbrebw5bAx5pmvnGnwHHX3IlvkTBrl94gI1KFt3
dripMp0jBiXuY/tk31ANIpQxaKkUcGyHzRqr5nrbLGsYId5nth95OwFfIH22iWEgjP/VzAeOvi1C
R86IqBj8PR78EnDc63j2hK8owkG7xXbAK+DvoJUsdzjWcn51O/4/bRNr/L8Pb1ETnY44QJPgZ+1A
HP86dG9TI0G3F5dqEHbWxzSA4OXljWyfl+TzN1dmDV4uAFxR340qG49zMmEeS4l0araaY0XtNP+b
9NgvnvTiwj7YEX0kw7AvVj2h73QxHTvUUZFKsYZOZDJiqTgc7HnvC5eFswFcqyQdFotZ2bLPZm1i
OQWsdITlrPQLIF7zLSgNiIUap1yhqI2KSlRVHJMdNF0bXB1b4dLjAniVpN+YIKkpcifr4XFi8KuO
dDXbs7HfxKA4lMYO6kdlNOmSkRC3XFqkyrnS5Qon4Slatt9XnxGJ3zhYXM9R3uQ5paDWGeQOmlMa
fmKutEXpSowcOpwtFls2m37U/CsLEEIjDe3OkwbEB5ivs0s13v9TYnJexOFHzvYd3AyUpJTSyfcr
ryH94U4nuWbu3mgOASuF1WrSrcXJgNsZ5zPjG0GiMIxAGMv2fhoEWaozRtvsRxARPtPlBkKe4QBK
63jmG2Vjk7VwE3Lf3dszhLD/+tNPBsS2u0weyvFXpu2bNsmAczDfoBqRWN5NhGZQUBdaHev3P1bt
oZdM1G+hcmduSlXs5a3AGpJ9F9OjDEOA1XH8MZ7zO0BkCBEOnXLzhRw4wnxubjbr/0URbxajCf3x
qwvQyXtKuMQlEDJ66jNIqGE3T8S+Ak3t4kaWErPRX8X4lnQ5i1ueA3wchNk6Bs0yzfF1zvn3+P0/
fdCVzg+pyeWAz1i92fKhsAXy7Kkl5Y8n2LiJrb6bydDp6nnidXsH7IhaSa7FHTxauqLgXxdkLqj4
PGCAmg+FqWrhxNma9GCesb48KDjXDOLXz206CZEYKVvR9Rsdfcjo8pmIqX/ZBLC3IkOGXFCmuZLY
9mwVjD9pvWkPVlfhQqEJ17VPoYvt3D6ymgoR9VE38xFVB7iC1o2zHXsVGkFzb4c1rUtzKb3UJk+B
hBe1OI1p3rfZhH53eSlyhVq+Xnd4cER8Id7Nu2JbzWpu+3UHlOtj6d8OcEeom0h3810b9Vvg6csY
vhPv2iwC8lM9lKyltxOC8Xwtx6cMSZD9UXdYTPHoq15f2k56pJ2P4HZB+bXnPfIg7URwJnOmL7qS
SJelbEuEymAhkSs8q1+bbLQPxT6PURIRIMnYKp2nXlsxzu8ErX4IkRVqxHZg8PxP2R6MbX3k2K9f
cohxA0Air9QJg+eQE4qgFKLa7kJFqZ4P4/nhv/yYejbBJZdB1KIJ/V5yNUGhH7yKj0ehsYZ3WnXZ
pJ6q97KuX6iDeLJJxHAoOz7pyeb3inFmTbpgBsrfwACPxQBqtgGUMvKHkryxQK8O9M2JQFvuotz4
Z9P4mQygkr7B364LCUjPDoIyxbiuHyYzDj97AUeYiwnSdSuDeCil31cJwjOi1s8uBzd3/TqvPJqh
mfqfZQkxnLxhab1+Is98kPiFT3ARIBd/6Hv0QawOHVwUdfSaQ2Wajrgw+gmPxuqppUqtEDEZ4Zns
feFdh66Lpi9SDJY/mA98K5AHfKqilokK4XO+ZPnp6G+YSMgMwgwUB5cfUx6W2NiRGdtJGtM5gSD1
NV7sBo2BQqWLYpxWuy0h90lDpEDnoeiLZl3ufmUozIQmcLHkVM11sJK14bkX4ufGAqkKmAozP6wN
SWq2QtpON6S/Gc5qhn9gWXlFF/aVnyJuhWD6dt3r2iKFlD9h5GCpAjP33Au0X8fIw/ao68mAliry
A+tW8I4EdH2ijwhi/SBzMUsIxTNNtCLDk2TKGGpCX4btw9PjTwuYm3qBCjMVmBV0F/x5sMnH8xzO
VESCcqVawfp5Stea7HNbY6rRVubiaGKcgMu/nHSg2LlpO1yTpjoIQ4rpg/5QUtBq8AHX4OVPSge5
BvDqr0P94LdCykHM/qlHl9yyH/PojK5ACl2cFDOrf8xAZduWZsidmnAfRIon/IqCR1lY+ckS0iFG
Oq1tvuJfH7PwZDwfl4YrQ1ax5YJijqWovVgnZcr7grjHWl/N/6LCjTGv0iKhgVM2W6A6bH5/3UXK
fjOX8PV7UuEQ22Zns4OTrGwRpG2D/hW+y7IU8x/4tBrmgCnv7C+z6kqyLV1EpTJCYH0HTd/vweEB
jATYX9FgdbyAnVOqKjDXzYsdpMVuJTjbZuwHXYR4h5wSFdbog3RFkFc6ZvRFCPC8jmDuvwWm5iZ4
RpIJ7vUEX3w1Am4arzLskAhUVGvbn3zSl+skoUoUBk6Ig8zPC3J5wS3xWhelCPXOsQG20B5DdEH/
hQAyfLAEuNQYepxn2lJip9sCu2e5IowolfklKyqwuiqoVSmjh8qrmTmvFEaiS63g5I62JCiFM1db
2ZtozQdcVYR0K8MkHYpDb2ldnsrFvrxdpaeBGp8woNYe2rGTIvX94ZmC0fZVujnUvx3ADIlI4Jbk
+kiQdZtJa7ymCxYXl111U8RCA2TD38eqBz37uvHZQKIDOGeEDCesouTmpL+NZOCiDlw38UPGHDFZ
zPXi5W2QOBWoDF5aoxgHksk3RggOorrr4NnaK1tO3vQKTIah/k9/n75ragJHnl79VUoiqqKB+oW1
QF1I+37QeYVTHeuPmsJt3s/N9LO3I7hcpw55J5ApUZmcUCJq0bx32V6IMJR6R+B/uGmz5gteqGnG
Ic0RMZVzpMQxf7D/lNn4egnNjJpdWDdRIRXJGpPsyEtC7ggxrM8w0ZVXisutlcZDOXir4cZ4eouP
5VmxGm97eas/8L1rnB9/6VwiqYvGOII41kxCYdulhZkSSQSZTXqdpIZe8lPHAw4oEjGC0qaw6BKo
BDYH5PW55B43UMaIfWaqaerL48YWUd3pO9MZupMVWSHPY+q0Gn3+5W0wZv0qB0fypku7RKqKqij+
RiHKRIeUOIrHIQj2aMHsLAuTvTgjThe2Y2eX+vzK45tuXpog8UZGtguVdFCLHpQneeu0oN3dfzIA
GhEVj2BqFo5FjBNtsdoO4nv3mSaOHfD4LYIwyY4g7DZWKvdOsVPR3+KF6HGIXs5WBdZ+6Cs+UU/c
84niNLxViIaQmDOBJ3a5nJIbL7OUqESy35SeU3C8aBSSWRTJno2Y072VVbe4xfrN3ux6bLy4n+N4
+Hr5XfsAH6MApJ/LSMyIZeNy40RjC2G7NQTIEfc58C0u91gQRnYcxqMiTtPNBPYu4Rt//SXq0iOX
F8UYRlfaGj81OysK1dl0z53qEi4bMG3rRAGmpAQnsTstjLc3HYE9VybMbagxhBGXytGiOWs8DoMD
bnCoX/cwQzRL0iJcnpHX5hTaJhWaP+K446ZhVCd9ojubt4d6iygyi7Z+hksCORrDfjLm3uj1iEuP
on8Hkrj5r0GoiNEV4xpSQ8cx0a0uGb2cwJ5jhuS96ZhwgNoY9dO4ApSHJF/i079VcdChOgxPMo6f
+SGR2nckc+iiZ+upJqcN9EEfVDgk0SuO9mpVDrS+A5ef0h7mFldXT3mA9FlKieKJM2aiwuB4RwMo
IoyiEP+r5YA4Z3KynVDaXC6iky+FjGuSAoCas15jy1YInEt4aeNPk80rT6DKIiSKAsMFQvkmd2th
DmXQeRc6nPrQ35xJ5Du7qmML2+prtlHCHv059YOGdvMIWQo9/3M5atzaEs3394z6ldwQPv2pXc/f
m+MkdHcsJ7EyX3YA2TCo0Ei/pMBZ4jmZHaM52nnTSes170BzelXA0FswOc7pEMtuXgwun0MZbY/L
oX/YlAJjGKde4UDfZ+N6gZnWZME+693SotYL3mO2O3S/r05M/h6du07X8p0+gOnAw3WXnO9OrwVq
OhC+OzzUM4Elf33VlkL4IGANgTjXo/C09CrwitCS6S0cVC82F84zW7PFaceN7uc3DMJI6fSwh1Lg
JeXSX6g3XG64cw1mh5Ur4cDmljkdS4ODrOUAH7MCO1YhE58S7eMtPuh9xC17SJOsQ+UAVhO1/fbA
OTl/E0/5LXymSYeVr/WcWdxb4LGmZ4HGTipfn+HF4tV6apyATbPx6vkUEinBsEStl4uGT9hsFuSb
m+2dfaaxK+UI0wCALBQdH2VlOPGHDY7GgsPhGbPjikOy492FYOA31DDXr/xObAQGwwsdRwNSLeOx
GGPgJtPudzOhbGiesI3rYG/GiCVKw+uSQGCvWENPPgJ6ftLMlWIX3Es+MZBf7oHKd7RHf1XabbYQ
rTo+Uy6vjv/lFT01D6byAlcSQNo5qgnH4sz/fcF15Tjf4vkdChnHCsy+SQ01fjx0GnYBSt9adxQQ
mYxBdNymcQZWuyMWAwYTwMPNyQX/h8UbZJvzJHnbhkQbh8NWWCNibQNDyb7jn8yfZ84Ase1khyH1
0LTC3tUBF0vSc1mHM9LmXDO1s43eNIdvW1dgf3kP2SNW3MJM49zH7CfGerUQ0dfVxSKVDLr+k2LD
hE76R21vJ0gy/tFeqLS0akK3I+5QvRdjsxlHy/WAK8Jweu80m/tpnk5vGlPBZhE2ufNosH97+IKS
AowwgaTKYiGvfn4KTN1oFXO22scImweJX5Yypv7V7L5AjstJfoXRPHjG0ge78bWKJHLlZD2M6lSY
f4DZuuD8fnBSZQRJ73UEPPEFNChKH7vRncS2vbhNTIsqAd9yQTexhbuKkHDmt262UCl0+D5NDLON
RoPEMfM4jluTcJgcFeba5feIglGa7bguTl/oDWRb9tRn4XrFmVZV3ESpLV7vyg8xwXtWjU/q6xLR
Q6UbEgH22Bo7XTsJOpK5zYHuvOSlS4rAY9i5vgVO5xkCg/yqQDDU8WbIeP25xxko2KrM4ufcxbcd
EtUDUzgVtJYv3kvq+fUUcA93F1xgQXxHnOwobfogkYY8EHw2ZQQdEKRrZEapKrwYDZGTR3313t65
D8eIqx1yORDEAbLR9yks7DTAdZSrDNqUeyyFtokfsD4fP/Z8EvpK19dNtUAjCQWHBdTl9wDIn1yt
uDmp9eyusbIFWoVs4CjvF6FZ4wEB8hGzY9nStFA+jfkCbO3Z0gK4BbUifNbnMo3PogaSHoRnhHUs
bm+2m8Fy1Biv7hUWCu4uv8XI9+1586to2TOghWvoSvxgM/uMzWILPUU7dlG30um+bDGONEZbwCGY
OmqjCJrIwShu1mqVsr0Js1C0fFB3qzEnIAn4mOzxGAFpwT7aiZBEDT/Onef9K3QUNADDxGlsglop
Y5eh+HZ4eEcIIS/T4CFBgj0t4PieM/QhAwJBymyEsIr2h8pQeh0ULTnM2KLHatOBYKQ6bZmRaVLb
wOG2Dj3N/hAIYTV/y68qLDQ6h9yKxTEbiaMJvP2Pa6OliiHbda1MUQuUP18kw53bQpBEA66swuE5
CD+4F4Amu0wRDG4mD4DMNwM2KfZLI+tRNu4okRceZlP3+SUtVMXh9gv6jqlNZD9++CrVXmN+pfqO
ZJjyGzMt8GljC3dAKb3e5JjRGbnOPKW7iRVdTYxTT4ec8yFGNqnpSOOHSLeauvtuaFqXecGBQ+Px
s7J/dnIcAmVNhpscXflzen5uX9Quk9WNBSA5FNI5U0rr5/cuie5wzwMYSB3lfL6Je5tjQSf8oQch
1kDG9U3S6OHCtpaV5RfXqJRagcQvKFpJTAKD7Ci8OC2cA+A4rx+wwq3Tplh5uS6S1kxTjznrjth7
1OQTI0I9A8qbScChfnzcEUGfwMh5B6qsiFF49UaudwQpLvPXecUSfznjgTsoQ34ZN0EoPFpVz8sy
gKGwpnp8vG5TKSZ0l0eOl4lVq4UxKzzhc3pNPCy8wYsXoyxbS/GeG2TJ9Iop/8x36X9m5tsVxPVx
3leax04vRfvFe21cPXZn0Qz1C8ghxElaaTgc1LWCaX+cZqpUIruDNZfKJFN6aZiUX6vQfk3xPQoW
C3ejSCtDasAYyJFnmt309ryT0TC7vvIM2WVwxv0dOtHRfLyNa28FE/zqaTiwie1po6aFFZKMUlSX
5ioZgZ47Q3hoi703LL6ft/eL5tfrxBEPVsiCsngYHHZO19C1BTHwH/r9Njhc9y0tkWc0TJ9xYksZ
0twkTF+2d3mVpwOj7zjLUpjMVLqvsRQQA3s63ICdKxfJs6PFRnyGIHivmer+GZQEp3DCtCfzNidW
DGKjpDAEAtWVexirPXP7t8v2bQXGyOx9988dUI1jSXN+hHSjcpoJUG/k4Nv9gCx+gmGsyZy5KrOB
aWhDQI6f6xiw0sELEWH/jP2cZE5JrZME/ZeNIHSJZBwJXZePRrUebKkPSKgvREF+w8JXNOTn8zRU
ptZIPw62jBldqBrpS6/kW7zm7uDvCPhLgk5D7zHHXnQkAiMjIOfyZfiw5c4eLNYa1lMboJLuuyRH
yeV4KN9wXW6mUIM5XBMPwYnAcUfASzbkhRPTlWPEM6a1+QLN9uiPqbweOXOZ7oFp6nAb9t4UV6vY
2vVc0BpNx6332tC29WvNUggposbc27V+9c08yVC4ddPsDPnSyrcDx4uSC+Btun1acroQ1LQ20ADD
ywFZAt6W1+1X9hFrDpxcI+HDhngzxUxq5Lzg1G3LTGQj5VhA4fvxlGuqQ1vQbW2fOE4F2lYusjzQ
mo8rVneuScXkAr6LnuWJ5CpTGHM1LPNRO2Ky6eBLSloJ4sZmHD0Psok7GmbeqU5tKpS43mAUN/Zx
Vc/sE1e7/V4b6BImeTwO3Vlq1WKiBd+U7eucrA1/cvugXnomngBfdb60lFYOJBfcK56hHTJ2tuFQ
Bki1ncWAKLqT5cM7Bj6Omo/dQ1U51pv5EpiwEl+vUtbk88tDEkEDC+yuFLkCEqMf/QlCfZ5k3jpF
unJV0qxvjgBUH8EpgIwJlsJH/nXvAE+U09ASpZXVLJd6+07O4O2lessJv/9yDJQhpTVfj1B5HaoI
C+m39dXRQNE82twMCOe4jv7ErHo8Ixwc/Jh7dvP9IDDAOwlFfmBiQKQA/mtcsPsdcGyf/EjBDHq7
7aklY6rHw7gkogGDvyqCmnjLW/DMTFSd31oRuFbiR5fLaa0bbpSqCPD1lufd0l+Yj8Q/CbCMy2uC
He5HDKf9XY9BeDyesgW2jQajRdwTrFVpfieAwvdm4HogmxBxzTN1+VYZ0V1V5b6iTKmw6k6xNm03
VQa/XdZBcl6rHWm4JWFK0zXcWgpOa5XUR6koKF4vpES9vhcRE9e07UJRWuAn4Zs6zVS8bajmbo3r
HsQR/ecDFwcQVQCYyoyF0OAiw1zrf94lSG6KFylFTrZtkKGmWaB6al9l8sSqs4sWh/7ewm71BTFu
xdlLchQjEdABljKnvPV7p1J1OuSBFVKprS3A53RL2s8Zf3J9BXSiMdR2oyZVUJkob3R73cAh4iZM
+vOIW/Si7W8NdY6+vq2nWaZCr2OTV6y/gRU6P5CjH2OMlYkMhggn6S59T5pYhxQE5DqcKtcgLMfn
19Mg9ZM2WzPwqwwSDGpBPqsFvcuADYLsluJC9XcBbHyjev3wguQRbKeO4yhYH5Hrxdmm9iIabaV6
sWtZKwiuHH2xdtfcGf+05Ou8b9a4oFsax3PJErxbvblsnfAo4JxQ+gfC90sbHHOqnJJ4Dnsnoiia
VUxAWBhzevXqd55ulkveYgDkp/y3045fDrbRzEOI95EZLxc09X8F7zuTX0IyLFU9DQmZTXt68xXG
/dfLuizXTm5Hvkz8IvY5JxOv4y5SLgBgFVacuHuOVWd4+TSCZQVjkfz0CJNkxv3IhTHZ32FCrs3t
jrmuJ4j5EKkCtSDHte8cBgaLjjQ7eMb3bmADLyK6O7TIJ3WHRzpJnBX4aUaW3S2AFUbcY5JJ5AFt
wnhQCzsUecvfVDJnLZnisUty1JoeyJwHSrNQzdakj9U7DP/XuG9Uy3Ew+iheXcH444f9MM01bFs9
TyVIKIbZ7q72v6PsSz4Aib9uit6kUpV2pALsOUNfhoN0uRHtP1jPQ/NQW2GroLe7dKraBIG2eTP8
kGE0cp/vzG4ck1XIvBJVjkWv8UdApmFU4ZGdjdyux3/FH/nqayFJ3msGiCx+QqZsBvSKOSaSFcRX
nKMNZLk1OJoIJ90lqcx21ZdyhupXBunerJYkJw61nkkU6JkQ/dnDJXDl3f/LdTtYsHu7GeqEWb1m
g8r+hqsWqPq+xA2QnyQBx69tIW0Q9sLh86zLCx86bc5ffsW3S9hdvagrg/lnot6iZsBRrAlpluw0
8UAtW2rK6od30PVYyTsGSbGqZYjwCa02TNJ4WLyDoDuRsmX/ZgxLeygI/FHFRT2+PBWNYsl/er+j
5R2MRShUxsqARfrruQdoQgqGNvakCVGYE+8bukr9VIcyglKmtrN0KsHMlgAjK4rrEKX/Ik/hJc4l
NBbdlNFcf4G3Qp5ljU8FW/6kQJODErUeP8I9q+8xHLlisUvypQh4mr2/+sRzZ65xszf4RZCgCEEE
XokufM7W7PQd/gj1RR72lyyxEbplSrz8PuyTPQmwIjiVs+EzjfwVKKXNsul4ZGv5cROZV2vEI6HK
qDdMV/RG4fWmWuSE11uONqfpHvWXPTEh3llwzG9vOQ+zpHZ2mvrcICATTw4y7ST7KG6/hNKKy8gG
asq7q93/mP7FZ0FTHvFdLuYCLgIEEQelBrcN2BtrhD8L2/Amax8m78VscHEW61ScLQUessrWEosR
447m/wWCkWgIbWTXxapKZPfmMOGh6isVkjY8vVXx5prIQXjnX0oKt/AQl0RcmusAjsi14xdqVuWW
c4QWFaf1h2Imp6M4GKNdzrXWjpcKrsmMMnL9ktSayNhVpDDQ7IxlR1n6aPWIpA5JofadBRrOt+SY
aq4J6BJRPrfmKhacIndE2g6mWLGlFJgPPstrkBgKBwQ9TydF1EPvxLiD3W+fJyZFO5tGueAmkkAN
qVUcsFh7SOl/98jqbxp0tcUubvg31OUEqKWGeD2utvN89UQWiZOGBv7xW6ZTYgO3TT1mT+lJejzM
lo6IOPwiwj3r3LK1byhPWACgcUgO6yaAoTtM4nQ5akp1InAMo3mc2eQlprMwu7ptSIuraM6LvkbG
u/KeLBeD6XE5KfmlVFihPXZXMXpuflTY9kqY/wAM/cJJgnA2wxuNDk9LWG6fRmH1lsw8PnFYfdDa
92FmSt9Q59gVZ7OW1ot8ucn6hfXutlKLi+Cr3RJeTNVZG8eN09mduZCRgBvvTSowvppysc/1rHv3
vYZvj6+JYxVtZD/nU5R9kLPLUf55HLn/TAfgP3nAo7+gBrecqWSVeAiARI9YlQGC2E7Ns4uCCYBG
gv5vyzb6H3DyUMCvBbDv8iJExH6bb+nKhgbpu6atfWK7SBaSTag7XDm+Yv+3G5RBS2sLJ+mqfQ+g
rNi8MK1qXt4tzSAM0jwa7yZ8LHO7Iz7gNFEknLwmyfjuriXwv1I4DSUb62QMQSu543+CyjP24n4+
HDvxBRYiYwo5Nsx+h3JfeSXSTnzm9+twb+SPOAPx7nopNvoiqXVUnibkFVh31h4N9ClWXH4LZlgc
+XThS9z3MjxmID0HQpd8jaiPgmDhhlXAHmQEV8BjPccvpoZosjuVXz8M/dAooaXcAFxnFVvhelDD
Xg8TsraiOfZFnL2U8NYJ7BUVbXqAliw+Ba/kp28hJak2WedItlATIe+gh5EbToTGjAcg2zKCrMGF
Q9fvUr3bhbfc/UKYSt2QVtQT79zZDhqGu7UwfrSPgIiBgPGLTH0ENDRd7v5rfsZbsW3AeVcchnM4
bUD7/xk5qYeJBgtGxmumdcDkdEvagg2S4FPUKXYXB4tsHCFQ4oaqOYvE4mGzE0xujQNVlzIowCac
IBquHq29lenH8NBV4idsmO/ZhJpJoMFdPO5NFkhNbhUhITafpZo9562r0cedLTvIfJ62QSBcPhQs
Rtnqrq/OJwCBdRG3tg8QvUp1AzWAV9GZ0rc/C4BzmXKAN+8oQtV+V7Rqvv3ulnzCs6a7djAwRWjk
eaEdQjTxfVIHWlEarJCVLhzaRBUY1XJuCFFV3A2fqQCGr8oRio4kmFgND0QN707D2A0gfu9zPhC6
xNqqNq7hJAuhuHst4g5OFI08vU8pM9i9pmOklXDOM2g4jAe+8Ywdh91nVYxVYRh9S3NF8F2VPpn7
LeYsAsbFRPVvezdrd5H0xqnEI1EdM4x3M22cxPPKSKhRq2aqzU7/ltw0XJfY5GPoLrFi2n+7vGWf
bdWbV74vfub/QpoMp9oP34/iDqv7fzy/C4yEGxH/lxwJ1KpQLnKTEI+1o7purhbAiFXsetRNF88F
Vk7kPGt2jt+8WhqWuBdV2veVlbVnAkGj4C2flLtcWoYTFd5lPyj29B3hGfeRcuNtBqmFYUWFZ7RO
zyy49B/dCvOzm7hL7cq55laXTEwDIq4u4qe83F8oEofw7eJyJb+v/N14VqYSUUkUUzUTaIkui/24
40JvzgRDdG2Tjcuy1McmbHCZpZ8NFO0vVMCZVhVvj6rhNBCQu1V2eXy+C+uoUkd7WMoIVijwxeBz
1MQ61EnESr+qm6bJCNOrOj8nvOTstXKoDJL8NybE/9Vx58Vz80kYnjImazOS+ZUUUybNbKTWCZcB
fZyjTm2hc13aLIkBl8qCOYky02WCoaDDH19AZubWZLI9sQ4xstxTcvNTwzY6WGQUBAJGseu9eN5x
taGLhqhLujyoYsuyvZpz3eQf8oxjpTR2Kt+ZoT8rnErx2rxw4R3iMd9cwBM3mdvGnopCcnFzlomg
WbmdH5e2DtJ+oCN0FyhX2cIun8a4J0uzv9jNxbS03QtcLee1WdgCnDsFMPIPKFqW2TG6VUi6Zpg2
B+wlUWVYJUJxXDfWwxJHa/rfxF9VQs1qZO6NnzWe2ZFf68EpgNKAyqpm+59vJgA6euKyI37Lu2Yh
z+H4dZT+Zpy0ty8Uj/lii0cOaQckhzZyRQJ+k9Xp27izYoopIaTS2GCzDs0QS6A5re5jgF+h5zfy
qoGTrOLhU5PsVOjcwz8ft84FYOPNCeHnfu2gpBKLzxFsnzzS9BCxi5n6AIXN+CjaCMeo+1JH7gB9
kc8Gq16pj127eTQwj9s0RpVWDoyAkYbkckaAwAaXNgUcyGK0JOcRmeGF9hqBA40HDd/EbgqESsfL
kh5l8bmcfhogGHjkax7ZnUdMtZiS7kJontoiCbwzdlkIPb0CQ7Oiyf7+AtvyY/S5BSsvdmLCx27R
YQ9STE54EnyZPgTZ8GtShDr7UKiznYPBH7oGDasHYHCpBveGIkK1N25E5L3ns8f/K7vpsU1s4f0K
jeTwv4Rcq2umtiOss/TJnXp2Uz3899ChFNpwrtqq+uyRYqldYNgioRBex14g4EiP5zHD/R1avuuH
ebn6YJM6Ogjqzend711q2L+0CoMzjIE/HGCXVlwkrr6v0L6tP/ZTSlOWf+wz55KNYMRn3kJOYQ7k
2DxJHvBfLn/7T22TX221ee5tlTakHyNuUPL7iAQYkBw16Og61KMWPirehX04cafS934SKCovwrzz
TiCZOx59H+paD8uGxn3YARYBoKJz2MvQsI13LJZoWsAdI3AgnJcMAhcVq4e+pcxmHuCRIWn9E3TG
3SHaSd5RkwtYBSEbrgaR2nvQ4W6D9YqKGlOrj7ahfcjns0mfUp1E4WQsj6jsN5/HfZmoWi9O4pGI
oyBnWyzaDf7926yBpxFwMKNvMczKmjhMXAwTBCsWCP48M+VP/t00lHm6xMaTRu7qJegStN2b6OwC
9NTqRFPAA2nqME1mn0/Hh4ZUrrRJp5VjmB/8VDHEfDZYKUw7m8iVw0eGkujzjsobfcqHFZFTkU9c
CumZANtg6wkku/4vh6zMrD2Bca0AToKfIzxFyr1ET0/Zju1W8adr2N4GR5HHk5oGR/OgP/16+v1D
UOlejzmbIoQLzAyXnwYx5vqzXHCcpV4djWCIj5exbam+r4rnat1LnUNR3VDVclKxWq9JsMLINTh1
/U2IeKegJzVhM9q+soh3lchkZIPICtUjzVYVcW1wMApca5G60EcO4aEFnez5jA8zSiGJ/gCNUooW
1sGQxE0+Qzie//477FcOl8DiaMqRK9Nt3Wg6GICNm3p4vmtF5gBciz9hRs0W16OP5RFsSgReZm/K
2z00/rJzFooo9W6Ult4XL+r7qaOdpwN5U/gC1glgwjY3hCAcNiK/k3ZDErM58SAfb/vh+OR1HIV+
WpH+8/dkawASgOf3y+qejZIOf+K8hYy80yC3tZBvCFQpsRSJ72DPq8PAB/wKFSV0CVA+v57cF1Gf
wqy7R1OK0/qnUj0bWcwfy42IeJ7kFeEZeHs6R7jR5bM468OXf4IAOyhw3w1om03QX6ZMy8UsHqm/
JbhYfWS+EvmzhGs+FvUtn8CL4TzZk+moroftuXSkg8C1wpLmXM1UcxY1noYRz0j5EZSn10vnDQZW
xQ4XNMMWdYnkReWa5ALzywvFcO/ifmMCp1vcrJYZqAbc4gm66+wXrs/31Sk3iH7XgwjrHh1/gLZb
ImSaIvMknYAgmuWmNYKetPR0NfBHVea8FlPErPsl/1CcDgIJIriVIY6Wpq+nRpTCsCtAM7gn1NBn
ycr1f7uENeyy8fnYwJTJtwom2h6zPnr/n3zFqKeSU2xzaDsLWJsGUdQ/rUqPa9rO5ZqsFCm1qFen
xBqKWZ2vsFqBBslx5vj8eA4d9o75vqVrsNAp02bMWYiwtPmqLSz64EvzEZ40Eh5JTcWJjILgg2sJ
UWB8FgCFIIzjlA7Gh14OrfY3M+ID1dMwUw7wZDgxPCCmiRY9SH+uVRDkRUBxoc4YwVpaq1HvHXys
qEgwNGffe9Px2x7Oq+VTItmfIJXWMtck9YvdaEQ4qlw00dL6vUIlsKYPUQl2phxz2Nm6phzGPDS3
KTnRTjWggzOuMssW1IebRwur9OzB4JgY2bfxosen71rs6i7J8gPiFtWvTbLcSrRVLW1U/kAlNbRV
jpW17fh7YMgGRu6EycosLF3Bc6g/P/NnVmSd62QQLxCAyA8k3UDjR8ny3jtNpzesdNe5fRUPCRJA
scoLh1MxhXd+7B82rG84st5w6TE4oRL6nH41y5vubuDJWX48dYY/Cn+QZLRcT5dSEwpGPm8uVl43
+8Vyx/xB15HZYnbS5E8t7Vi8gE/13OxCua7MoW5zoanCxdCw3RJ0zSbxXeLs0BvDkyCpB/viW4dF
3hB8nnXu/5HmeHZMV87pjK1kmG97OwonXiqrGEE79dUKL6cVqOWPjrqDw9RNPtMlSCknZw1Ho81x
9JtoiAmKhv2dlkmbPF/TKyKTz75Nt2SDAx2xpPy3ylpvPyb8tx4+oH7AbX0WgwLPmNwMTSxpnX4l
sMB40ECAZRRtmUs4Tdeu90cBiT79qUWCdMQgDeDkCb46ttnZUKcHv+Ioyo/dcOE9is28akXdBEHb
pSeY0stnnRHOKfmU2k3AY06bAU6SbEJYBvVI5ifUsl8KAy7GrmjNPet5Uz/RRD7qjCEKq81/3/+X
Lu/wIP76FEZ74RX5S7lCNTkCsHt2hADgoa19PnIh0t/IObYLtZak9ybGa3n5sV9ynB5tOOEofpbL
FpgswUEWHUifJd3XXcuLRYo4iNiXvQ4NL41hOvJ5G3X5nBt4GxDjdutGqxcmruMJs2ArGAqSvEUN
32RBrJy1zyR1BhKbU0vGElf3Zi2qlIl2mmo3WMBXrRtxBQ/a4eWacbTWmIy/323cMepRUDHzgx+k
CkYUIWQugajVxtIZawGKk+FCu8c9b7UuXkhSlggmJzwe1CNwQyg4wfc1fZmfXpREOFJKmabdJ75X
YlbiyxwaJwJ58iHfOfE8oYml9TXw43ws7xHzSLnnLflItHGG1ayOhH5vGkK9M+kCVgHXuvY9865O
aDDM0tJqACycjJj6qiH+rDIYAS8Jry+y6EBmVbY1J5dxQJ1zt1LO37fwuQIjO4wXcAw4WUAbQqdZ
E30k+3ICFJs5gW2J8ldQlL3wchwQqke/SB5YhnZ9SCK7rNQEJw663bVuERbMCze76mt0FGXrN7UM
82Q7VuxLbPotWZaah3yRmvBs1QtX2rMDwJXxyAcpNspTauYxod7g6qddQB3k7M4hbBGcaIMFOGzS
JNO2W6myMibZZzmsiDh6842fgKhpb1HZ2QVla3MHOccqn+MmBF1Aab6PsMzbKxZ1JDSILiwArSVJ
Uyc2rmQCErV4gDQJIJtq9LaKLsHHpDyjr6BNa/CPfOA6CLr/Dsd1VGc+33eJFH1l79yNzfdKMHO1
J74O3nKJG4UfLMklaS0DPRlNLJa1GHuBberOvgTBaJ5+BRm5sC/zfoJUrVio9cTHKWvnprsIAFba
bkVsrkbh3PaoHUb9iwRLbL/GOpAATNZC3DzU3PeDfzQH8jya7iwEK+QGobFKemxwmNdz5gYsHP32
P+A5XgIVRdnm8GmZ0fXm7ISmiV9NwMNY8vf5KTzEYsdyW0q9LRQgpKJdpBvQkxXm7NPIdIsmxU1A
zZFZ+RgGsg8Ar3m3XgRm/BL5yzfJR/zFWoz81jOmH2JGQJjbidb/7M9JSBNoL5nK6bM777oCE5pN
9EPfRFWSZYO1QuCBewgsgVDMmgLsqCP6wxRPRFUAXFrFsgj9z0S0UCvWkbnsc6DQSDNJSZXlSesX
7paqN5r8sivvDBy/ztC29HwmC2zJWX4Bmlvym2LSUUgtvLC47zz3pUmYF2AVF1ca0YDTufRNHGsk
HIYK+bmuQsCRWPfZL8zdy71tCnq1UF22otqCnqFpGpy9GS/C9P4KRVgaPAU7ZqW3/6zQR4gVTiel
T3u59sa+t4EXbBH2OAd4pdBrbbdYSkXAjvQEIrl2RcLvwTx+c8nC7h+NzJQXqbkBNBxIfe1pXcPo
d5e1rJ7UmpyzdGoEQ7yqdDi8OM7LISuLNmECqTTl8p9PX6Y9iALnTD7A1M/wh74Vsh3ldik7Vxdf
6QanEFtEaKer/pvwMH1xiHTQYh2RQe4F12V3WHYzfLn6uGQTIWiQXXqmX4e0c8laVieKacV3yPM2
b+aQiFnKr2iUGQN1gz7XI6F1j6KR49Ll7k6+rtcdaOvjLRg/QJIXbbytCetsPcYTpVJGjFO2N8BH
lh5MiQMuCrvYFmkYoMYkam2m1uAkSVUAn9mOuYykFaMWC4HLghRYQ7J7YaPY+sWRhB0d6RFU7gc4
/yFLQW4Kk6PVUySlyqLh/7IGrHCKu1I4w7aPIWKDje7K+Z/yXaGqIzfbFdzvcoj2WztYifzwst73
d599dMpQCm8YbRgV6PKZ4GQmC0k+qNxJ1j1hoi32J9/ptK4DlVf7JeNIV32DCtWtUbWRxgzjD8fc
iyiIYqtYiqs1AHn23C0hd/aHWTyWORI2joTWmxQYhJYI7A/lzKLhYoIt+JVaevFmSM03cW/dhVHo
7mrjoQNP4gNTr7Ulhxv058ABi1ZfeYmVhfD8O3vaem85M8zwbQpS+ceoEvQ9+Z6CP2VtpmEXvfQk
6tFLxoMlTtm1cXIcYtYMIyzaQWK9VXWBeBfmwYJQ2Q26lq9DwSr8XgrRkGhxOsHMvDDJy4h2N1W3
k2QU9bm5ZtI4OjbCsF8OgVs6wxL7KWtxsHooxnIO01TR2kVY6nwG1/ZlDBXAo5YGs+dEX2tc0wdX
IN6uO+zbap/D2g8qB4uKdCunPl4VvBqIhnPiv0ZiYLHz4OTMd+DFMdZ8Gm2eqk2vJKNKDPGpaz4o
Nj2naEN0Lq3zq4LJY2P0r/aLxEAmZ+UDR1u28ixIIf595ZS8R3Kg3rpdO8BmIUoGpoDFDqIGpadp
fuaryHHJKWZhPbthMUT2DJfDzhB9mMrK5R/EbbnuFjLB27/X6Hd5Zd3nqaTFOtM/3wUCo4Nws0vY
x/01eebHd6vHTAZKWxCZKyLjZLMWsLJIi2PCjhAX7muL8xcSJjloFIPNUuO2RhGo0e2/R1KZPm8A
aYWYvWvB/LKCR9xIld3mH8sMvDVfvzGLUWmKIant92sYgX69DdxKP7UNdSr6SNqWd37TXJVtwQzD
gaRv7axZnVfVakgVZ/r1bN/04AoXFFX7oFsOppGKLVOU/X72ZQ9kWZhVABGd7S5A1QW2JqDQH49V
3Kg7UGXhQdNKUF9pBi5wsL/zZ7b0Gtov/Pw1NiIK705AmDp2m3G8ocTaOy8qjmyrY+L8Nk5dtNhO
ktCfHqUxyC+J4/oXbc3CZW2vHrbEAhX7j0ptMKS1DbEgjqOoKACEjMlX1XsdDf2tAtgmSC/aTKQH
xWMtb//9gR3ND2EaUzF3FD70+WwfLNXZdQOd+egbwsiqLCYIp13pRilHDQedSnfb6HWFKHEDV88p
GqBP1b5RYfWJPBA2VpgsmQWO5hUa2HJCO2cxtcshA8KCpdQ1gVCkoMjIYTboh8V+NKETvVHlflsV
v+huQhvABjMcvs+0OY5u6hf02EAPFeaHK7Agstt1GSyT8LwiJL8N7mZ995cWaG3MQ/Yue6LeZcwb
3Tj/Fp7FraRqlFHjVfAs4353O31QdZsr4exuSYgJhQiN37FajTpMJIVZj8NDhIBFieJgKIrmcJ9X
Fu46J2sDwN70S/HZ/yU96syPnZ3UxSef5b1wEavlY2RPQh5v3/U6gzpnQoG1GFsRs4kyORtJQL/f
XEaV1w63e0D1JK++sgmTxM3bLDzkaRAKr/Wwv5E0oZVX41kVbRc9e6sqMINJxxlOERNlc1N5S/Jh
atptch/rMuJlCMj2RWRcsVsWdWiEwXn5zoWvFp8Jnw74/BDsL/I6BOXzLExbhIXWvU8/fxfR5f82
p3sGyPIQFQ262HCD9mWOzkcWMYhUzBzB4nYU/BcvBdNpHLChf5k/rrBdXBhJJhpQ0W2aOhjG/wQs
0CZiHDBVvh1wy3rjb2oIQrVntsXhJp7EC7a8tgqipecXC589+8c9NNGpR54/WxND/8yrtoifh5OU
71S7DOwrEd/aSJayh/WUhPrj9Ic1rMbJTpZkiLUl9wExlziR22hgvuh2qJq8WJwXJNyKvYl0tpMp
8gEDqFasVqfMaaA06YCu+f9zRfiBFv+xQE8ZPDWXrzns9OUGo7GSTwmAlNLiwkPBox8ZXlubD6kA
9ghTQfd1fyv1zAGG9slvsOn2DGLqd+U8jnQff8vrbr2J/WKStPAbbW4q3kOiMjcybg8/UYWu2Ii2
Qdu5YgoYVWi1L5gqWW/KfLZ5AosBUQu/7u1lOIo+jpyk23qLQdc+XIr1COFvMY+InK8/BnO3telQ
ypSbZ8nEj2VgbW/6ISOqnDDSOURuJ81gnS58vgxExvbIzhf11YrAkn+GNSFagohn0Q79E3J6hP5V
ljAeeWZaZAebBW8RJc0OSLVVDh7VYonon5QDcB8INz6qMX3jxkXE08SsGV53tVtSkdoTl6Wb2Wf3
+K370p6T9Nv+ysQcFreeQWrFKawagQ/JnybTUXIfdj/U30bYpYmhNUf8Ht+n5JBeJXSV4WQqp6k4
/cRAb93RpXqWkATzfpBUvL/W4FQg3oMtYqww332ii0430nHZsDU9rk6DO2goj9QGCo2eLhtdwjxd
miM+3LvlJIRs7jP30IH1/AByVxy8+sE6txZKx5zy2LcSJ5SEQp8k9hCFTLbIez5XkepgHIEXNr1q
TX7wjTtwSICfK08WpO6fSTQlogQ17VR9yLc5wo13KvBue7Zp57mBwQ7KONL/bUvuJZoQdIf8oM0E
z2JYSn3kr4dcOJaXmQhA8YAF9pK4M3XTS6KINyVjoFm20/bQx+bTgDRRphUkE2aez9oa0GNIiA6U
Kwp9msqwXDaf0HnMoknLb7Hq7H8/mkOsUiOiUV0mslqSc3Mlg8XXnKvOp3Rhtd7ISEucSM6NAOgZ
Y/+OXk2irB4BuBmRviRu6RusRk1771c8ZveZf1SUKDIOA2GOH6YYxmTBqfHlKcrQDuysMjUW2E0d
+DoWu/2dvGiQNhjGOYIkOi+E9HGfv+1yLMVfVF/JwiMMlVBvjVvKX1wDli2eqrbEyUtn7DyLso7l
3s38SO4fT1k4UVnUIvgZBOdH4Zwv13jGgWolgRIqPHfW6RK9NAfmTwwe1/6yvGZpaMoSMYXLi9NC
iXwYQcCYhUGJ6Elt+vhjXWYvMlcKGPFnpZ0AAcobwT9y2lGglUyKeYs4yWHPnB4+ZF3/Hv6SQH7x
UCjiFw0jZXCBzcpWMibev5CDwd0s2ExQeuc89QWaOhO5F4RotEkcj2+ktrvqhBKPj8Ra8E1mGJNE
cEUDCorihkxdwc6nEhe2xQfsfqRmDuVUHEDg8i7/VHr2Z5Ptvz3QrgFJRldmOE0dC7TAV8NYJguM
BbUVpYwCMu0jr4+Gw0W+9NxbjuYUftse30T76fuVYR22mSBcwUonTJCs6gOVRuaA4qMJIkFy7YJh
lhZzXkScBdRKEJdl98qeKOahk3slskD9fkQARvpvyJn08I5oh2ngGh5lT0dEFjlq/57S/LzffzzM
y6sVk1D+KscHJ8IsRqMCGvu6uWQOcKLE21UlEbzHfaBhk6pyHLQVPdWnPMND0182Vm31WIVR7LOi
mM1I+08NmozPdm49P5LSDhwWvPp9jt9TcnGLLKCNYR1Q7GU55yA/jD6milOLAlXO+2g8Pr8v7Ola
mGx/Sr828sc18cqAlF5PQdcRIdnnAG74BrnAANeDXxZYbmrkLh40Hd6Dgx6OMEsDU3Nd95Sa3WBi
a4MuIvuM8Hrp2rdydIxWlfaFyYmMavvkLIIVHAlxZFuNc1B7jzQxUhg+cK0szz9b4FPm8o1bWWC/
cg6K5xwMqHZGsCgHBEPce7xH/y10fgRyShIX1Y3XRNxFOHIeodZBJ0jqxR9/JObl/GcMKFqMEEK3
2i1ueEsoG8BNCBt86CR6jxcg7hh0ej2+9NhN/IZONKuFcFD8UTjEGfZXUtzMrH60yqYeunbcSHuy
uZ4Dxm0uqalpCV4El82zhEf8HbVeTs68crH1EK1IbiQ5t/B3RNfw6Cq4TdVvRv+Q3JDcdHVQ0SGq
/Vy2Nqv6ZdVnd+Y7pdh1y9LDy9WQfI2vL8r+5JzCntEbv1DSBe5czNi4hEVorrRltF955d5i4m0V
ucpTh7s4hMfvaC/R09HuIwQ8fO+k2jFVuwaWoflP0Xa3GXiaIUC+XvE/0PtE0AiF+E6WPwbEB2j2
Dk9F58EFii3Twg1QmukcaAUO8r6fW+J1hEaDjW0Od1Iri0pX6BNtxTM7d5E7skAMuj3B0b5vW1xA
/U9C321pGuwHFsSeuXs8TVh6i8rUxCmRVAzpIngeN6oILyTyl+dl+sjgWdAvSxK7mTdFc3qUyqfH
wdqmVjDAyjGrwPmyrt0X1c51HqkU4W+Zkpap5CeOqdMfCFDoYO33phv6cBYmTVerTBKcWPdHT4Jb
/h9wrZqSMW4OutEmf5ZCrsh/+uDFIeuWQsASTdYjjGa+WGNxy6PJ1NNTFWj5s1ldqzzp7r/PDs71
A2EsF0zWrEqu+nmK+z51KGDelQy0fqa6ceBUFbZuTYeZo7wQwrZ0uzp4MzATXsr28gFn2iwm2Hgh
yxGyxZG4bEHpPtSJUkROwy6U6xrzmTZGg/3K1HLpXPkRqLs1eHf9yT1H4ktrraQy4hJxw4dV3JBU
Jw6IP6e47W/QFJCduXsgBdNkLsg94Ar5C7ixPbW5aYDIzaWYlIhZug6R9O32f1ifu2fHHNuD/cLo
cXhamBguqzX0o2RX+0zQlcvanV4mU9mVM4QleR3reAiVXpSzn4+vRLYOAXVLobKhKOFaFurqWNGP
c1bJ3A+XRQfL+cnrNmabfoNYn7dNZLxCg6C4Dm2CnvJMIo7vRyxcqAXiYNZEmJDr1puVJyOmiIu+
kvZYAGg3gnHKJp0wvqL9b4V1JvjgYO/MVY+iEAr8yg9kwIMLU4C5Dx+ppHl+lufvrIrQRYD50WiF
DAluAQQMG+ya0nsTqjw54KqMi5+TW8tfoz/3vRG8OVfETmiPL1Wsw/zLJwCXYzqaQr/jDzIMF+QP
mmft0XKwJ8EUpq4A4fSjXnfm1dN3L3aY5r1klgZrT51RUudYJoVQnKe0GnjLSRXXPk38agsVLb61
mipCvLtEYF0vfqorgc+s624zoMRoNX31+fU3LeUK2/O5NiPaXqCGCe6UThGxX3VnX0MlrpYJvI9g
mnZARxMh8S4802c1/Tu7XKRW5Soey4qkHLJM5glwpRRPJkP5gPjFGoPJfc4w6hUzR1jcppHv19wl
LLlnxFiMo4Lh2OZPHUyHsoMRMJ+wCcLWlyxdfzam7nHTNE39WU0XOm/nRO5JwmcXzwHRKNXbncVP
Abxudk+jG+/nlFIUwBUz2fo7hAjnwNCk7fTSWCmR97Gd8qZFLd56MGtIwkplwWfFTSfFVDcqqWIi
tVk2jRAWeFVvdkkGsdPd46u6BxhYT1VoBUZbkgdMjI9de6jD3sS1iilJliMjcumD5ObjTZgv7+11
QsrJT6yAyGWkYdpJUv1kO66q0Oe6BDXmqdmHCTixFYxZI10MCt5kdVl1L5I5TC4s3dLC/aAXN1yP
XF3tRJKYOFsBIbhTrAzcNQ7b/d631I8fpWKpWjt44ax3Y3WHvcL1RgyIy3CnGteVMDxD8S1HcCzz
SAvadoWZVbbBGsAJsB1FQC5sHUwzXiKNNgx+R4bw3JD8jXy2Lj6/DRe9px7Xpp900ZTluVNVeP8k
ZzDaaxNT89zT3d4h2oT9LLzWqZ5NNpVduKX7ZuIAEVFRAHsGi25as15bV91jZ/TCpjambwAfJ3MJ
mJltWalJCbuIbs9FUtiGsC3PtNQr9ZrKdzMK4x/ZKr3KVWin0H1QWxAcQRUDaBTNxmc4DeZjyQk2
cpefx2X5fXCPGyX35bgVsxvbSdLiy24XHYZXJ5+BeTiykc298bfdGHVR5v0IKZuSjZgSK9D3SfLV
GcgeWqSOrogT90pfVt6akcGr0xWsbJ7mgVHJnvqM34r0milXwiu8quefMlBRi9tt9+wsii10o7cV
9sDtJQ076L065xAr1nE1AgcN/IsGMjtcGW3CNDOMfqpgE+sH3C1tuEpL2d1lSItmGT5pV8wK2mUe
yqMRF55VuBgSLnInns7eejUsxUEUged7p/vFAeD5nSiXbLda8me1/ATDSjBFOISqKFK1dEwLhvTy
/qu0FbykmC0HtngWvos/NkngssIUJljMsLx3S5/dqvBMU96x4DrsD9sFbPT0c2/fbMzcIt3dImIb
RDRIudX4zPY+5kGrsv1/6VFX7e89+1f1RNQ8nrX0auV8T++GbncYjMT4IgVzXrbm/bRMhwtwUbg9
z88FQ2ZKniDrFr6mjzjVyUHmKur9tQAjJMkgqEfH3j67+SHmEIE2GY9G5mEh+nvY8IpTpxJp5MZI
jGgnvd26DydZY81uSUmrxj/sCHycU0entjEULW8AQu+1Xz4wE5Rh8B3mysIUJiyb98R5KBqpHZKW
3e8YECjc9jMyTkLHoitOFvEOIyERhwXl5yO+Am+++e7SREUOxNsjeZwfOjWVqUCQGFDkjb3xTVo6
8lCvU9jekcc0Z0CP9EpXXthroPBS8EW2H/5XVkE1Pp/emO6ROYqFSQc0mVJT4llOFPexajEcdQkF
ts7MKuWiy4KDrNWISkXFdIvKewpOW/83Feu+mOgVfa3GK0TiCLnezFoEAtb5R6fUR081HKqdLE2T
3/o7GGTV873Pryq+dqbJQQBKjDY2kM5P+VOgtAbO461ZmHtHV/kmf4Ojb7ys0if2y/wKq6pUyPqj
Aar0QWEcz3RcN0OQQRJ4opwTzTOKKT1YIJQmvbL2tdK6/BcrwLJNhqYlHuQvTzXC5xZ5Dq0Hiiuk
8pVPKc6AtPriyBo5x4vruPPa1pDjClzcdi3i6uj9LEOPGSmRknavwhFCcNtSFAlo0alwPsCPi/3f
q0ZK73wQEx3uEba9XajMVt0mpoPNsjpV6vAofKqILMabWSc57cD8vztwC8NWAlbb8EjLrCFl6PM4
zfKs9eqQlU8X8eldQwoI+SK0swqGv8/4r9yt3F3m81H0DR7xZRuxOKjUQ/2VNp7f03i4yIstZ6rU
Y/sOdc1dMeeHmU357IZ4WC2UwYuUlNm5qm5DmOKcycoSoHRHDt+u4id705L+s+8KuFNlyS4gYCyE
Z29jZ40OU8rJWt6190bCPxzTTI9Pp1JjCw+DNyBoat2negQ+C6CrXVHDrLPV7IwiVjhXk70FicuE
5Wpeq8/4p2bzMoQUHxuZwMeto7PKidhtNI067EYr8GSI1O6AmfJr17dt49GABk+qS9WFVzusbw3m
5FOyL6xLGK6jlM+1BiK21mbnT96SMTPmArFSHmqMflQihUKrSZUfXct37NtRbZmybPUbSWjHVlYe
YAEl7hU+fHysZTZjeNo1oFAmAuwUBO6yOTEwUg6sMlIBN6+54Q+MVL9zaz7QoKYPeeYZ/VswSM8s
NtB/EPnmZ69BteDRXKc0zuud632l3l0XAoNuYX8ZvTIK9h45i5p5hjWaHNfRXdRfqkxNimDl95H8
U8goxwcGsNsWuvNlwSeXRmDi6DR7bv4jpqhbeVReszL3GqlDobZ3jW53nh5L4haDFXh8qpZ4A2Ax
ddAvtVNFJmioL+4tFT4rMsTg1dXLrQuOIZ3fSbpvPNyN1S8go3GbYitXtxZKt2943Ki++bMMAq97
cJp8FaK7Tdrohds+7T0b88+1euLxS7gRIgDlpf2DX7FBsOgr2L4zcCeeuKEEKUDIOrtJ3MDk79HY
Hkmd+QT+3sAAMRB+59cOUAS2q0LK++UQq3aS1oTaLk9oKZKeUgWQ8ls7NXc11Rres1vee8UvGR3U
Mvb6QSK26dMPag/YjH7/kAo8YaZTv7IZg6TVceqCunzmkq+MMUlO+jRKXIlDaXGibFvHffo36h+b
esJ7akYUmFr3Y8TVt1rkYPdEE/G9xE1/bRb5urigtZLVcy3tmYq2sTJnP/mAKaji7r1OWDA0Bf5T
CYGFFuJoNNb8NW+epm60If9I3hNm1MLOJG+8S2UcUfNyMjcTLizGHn44SaUz48zWGOkhpqkDLvUj
3JD/YpHOcBgeeoUmt8pLQsyUkaRsU883HVE+rZoFPsM5wiyPevVF36l0Vn7kuSh0s+RFq3H0NNSz
kRqWWMCIUrC7UtHD6EHCR2KF0rjjah8BxNVddDlP3+CBAOSVQ8dLmvSAjUvObLERxbwWDtAwsK8e
P7k444VkY3LMYnALoSi+xigP/HeY+dRzNcHzsRPmg2t2YQctYxGl4YdcP4XUQ8wD66btkx4MhIV3
GgVonrCpPuPHoDUiuSMRALbokU38YT5An7CZDtSlAha2Fmqca/sYKq+beufQXtvHbH04NmBo53hW
xwPzrbJi/LClIY2XZG/NZ1Uoy9gXt9ZnCDnGXndOhJ/VUO4eqhddLz/IUpZG6/+wISPA+0prePWB
FNyEfAn/TyQVYSOv5I5coqDYP+RusE3XyX6Orzm0rfLw3EB2CqU7d1xUuTJhlSMI6itFdIsZkVJ9
t7S9Svy8/3mPvoDY+/7xZnww0TjkaHdslRCOMAnxOzxDJOP9UmGHLeL8Lcr3lmyRcSta2Xut/Nr4
vCXpSTXsemPVXfxDWJhGq50lqins/eNQggLXimpnLrrCTKEIdoS5FpTjcrijjILNqhuwFpBZGj4h
1n4df3VfZCGpHF45aeYOIyCYvr/v/LgF9yezJJ/AR5jAEMeEp8ynaioT9kD+kI7g/xp2wCbXXyIh
TAUTIQ/T4myQ34LmPG1CjIUVqhGKSXBX+XZWgq32+VmMGkFnQOd34tbRk2forQunIMUpmuYtAwcX
UzukHgobh9MrlBcJoRpk+Zzl/FU3eI5aNoLoi3enaa6T5ZOmQ4qUQJ91eKXhg3vdhANq3ohFkYXY
f5dr9tsLGRqDFQObGlrPpp545YSljKZUvvOysbCY0tMmwOPMQjHH/XTgoSGGe3TpR6Al3yEnRRcT
dEpRMU9d/9d662LvA9R/PlPHxqNdWFOnZvBDBY8Arh9pudGv5qcFMJ8TP0DKO4znpI0iZirKP6k7
r3Xm+HzhwpdJxhko8+L0yCd0pKGn0b/nW9J7oQxMceaNtCTe6g6lSFl/rxvEjfnIQRNEUVg10XXo
OYqw3lYEkw2zUiWeKtfJI1HBLmct+141Q14qTQjD78v61cv+ff5bSXSmo88zeTS0uHIEcyHJuxw5
Aoxo5wH90qmDdz0fQiLLid/d5oxMlE2RhVDS3eTK0ydWsdiD9syBFCTd8eods3LKtGnVRvoYU24i
UHh50HzHacSMlcmRbhxJTw80Go7hJsvcKdoWotuYrDBX3DSmSCymfN1g/FuzJAuIcWHID9mxqb4s
l3ldAzpGM7RQ706nJWgJISl5HIdSxgh/9YDsqLDZLsTqMmZ854xox3aJrMwRduE0wvBeY66sl2PA
+ki6B0WZXrSKx5Y0Aon6E+2xrHb36wIvS5t7UoAgFPM6rNw4qkRWikZO6sxX5MCArr3J8JcWbHtq
SUw2CVaJcIX3E4A1hzM1WvO33PiBzPgSPYgd3xjCphlkMsXrNbx2mnOhruCu+DIhgPR+MMAnSnFs
lsTQ6ClraGocUY8NmY8KZUUwfGHUFwSwaRK4EZ4jKWfXaIow/AN1PcorQrhlgkbrItecgmxs8W9/
GB6PKi1QCvwe66h+j1NRpSJb74sQjod1/VEdthZYt8cDDtKKV7wvrhjyKz9CbjK3Ax7HI3iFTFwc
LqPBLxUr1+BuFomUAlOfVQexGa2R3EHm0P+WHfkLNukrOtV7dc99QoCDT7y4TLMXpYRIuAZ7Z/k5
sJ9sHPYA/T+/B4Qp+v7IDV9hwiTFqKo1aNzr7J2zcPDya8UMvEMXyZVHeEW7Xvvz4zHW8ILRecfx
w14ZVTzuMjSkotaygs0OIv825FYo9KO5K7cW7X43KcGA1CVGqUBC7Um6V6tTOPnJuHsQlKmd3Qi0
7trRke4a1rZdSgyZ0c5TxAn2RAYIINU0a7JnLsMCIPKyNNUK2q09LgQ2eyUkXe+uaEQkomdHVea6
gahaFR0UJ7lEuT8z097GBE7uaBgeN5j60J8dEBLjgFwQ5F0ShPa6uCYF306FqCV9Cmc0EUme/mXY
mWOLJvbK/zr8iwnfRnDAhhrDHlCPOLnDjdXuSeuRU1fjdsSwdIv6nQ8pafmrC8qKoEiXvRhdSnou
b9DPk9SaX9PRdx01vw/cLe1qmCBapqyhhyVv7ttZ3/t7xTgaWDG6HkXx+V4chQv5g9Sbsn9WHkSq
ot9Tt8S77caJkTkpS/rIwaP49bd+Yw6YMlxS1e78k+rpmV+X8EMieuf1L7vJMbEN+uayfB9ugbT5
MpRK5iLdT7fgYUdXfxCB5JhL9qO7RORkq1AgC6OtycmoVpRepFZBvd9J34ype6k96K3uDjxXnLOp
Z77vcueibw/N4qNNsBJKbXZoEsxKFOPpB5yfb9mQAxLVAjNlh+XeQQHqQDf+sbWIW1cVzEfH4qtf
C8sqQNOIJfG4z01uycO45DxjBRDhm5ABBqUq5tPSkOvgqHtXJNu7kw5MYe5My2DB3/iKXGBRRjKG
gd/VXBZm2JueWHw1EqURimW9xC6YfLPzO82R6kL4Qkkj67vf2T7fa5I6sxqr9mpbUsW9cLLz1sda
Y+nzPt1OSHHW32zyYhapmm7InlXFzFXskrL8OIvuAhPEuo8zzpyHPqjkhL6B/8FSE87vM1KH2oWL
xZCCOtfPsmUUh9PONkkqjY+YOkhIJiPDARFxGmAKW7orLsQP9dgw4Ao8yTJ6qrtTRBwldbaTF7yn
3TIpFNx6Ff1J/jNSc993DRDLo5siunwhdB3WGN2XjTQWiEorKoximiF6WWsNRpUolQSqZ3GXlSv/
g9f0xV4WghYuNbiDQAjCA4N4BILkRPe5S4fdRVK9lwowYQsJ+HPXzfs+y8RzBPGgDqZrMFVsXOKK
7XrpL/opoCgiLhQjdvFMZOirD0qKVTW2Cb9Z9jfY61AB6GBrMMkUAg2vMacz9Ox88ZI8Kukcu5NS
6Um01ObyPozQhH3kI8Qeo3AYl9wurKEWrOGyZ4UamsGcKpYCcvbAwhYS7LjjV7Se/XI3w5j0w8FT
WTzFyaUfMDL6PMbPtaTbWw80X+oVRi2M2yby9F29tIvNbIkE5wHTj3NjyyQpHkEEVmsqnyQBbTjT
WeLH5eUOCXCyvhzUPhYfJDMy0WvjgIWh/hwuuAOsCMRgOooJe4bR+js78jnqsjMMlG9KUCTfUCy0
pPZnZvt3LtUvac9/aeWoBiw90A6A4SL/qWcaL7FJqZyz2yj11+qzoVn7GhxWnoJFD02X0G7UvEkU
0Sem+YewSYTrTLCZddFWUjqD5YG3XyoHx2jGYACufz3hQm5iEC+Q/sd4jwsyLjMeCeeSy5QJ9/cd
8L32zEzNcNJj5FulzHz9gOx7Ed34V90EzJmdjNncV1M3CnF16v0JjWQW+2o3EAx0/SnuKmC+jAJo
6DtqfFwUSrMlFyGndJzS77mC+EmtG9xQluM7NyRbHNX3bIhVsY/8yd2ZVJqVMcsuNhJMYkDX3T8Y
M9r+qigz0ADsjUr8CsQdwS5fitoSALjfJ90tjDL4w7iqXCLXyYlmxKviWXlZ6Dm82K3FzX15yN61
RKRajwKTGyVU6SVEtItC/qf5LxJfhWNfUEY0uKNkLoWBxSQ37ZJETmfPgMl4QKB7+kgvWx+dLq0E
cm28VPjr5KQbWh1Rjkdd0xoRcm+2LX1FP3xStZXGpKrpOavR/SipxmQd6B02H/LbE0x/w6DccyPq
HWVCGRF3+tfN/d5mUXb45eaU375eMT2HhN+nScPMZry9p/dJBot30jhzfE4PqTO6vLKcd5IRzo4R
3gtJQlnpr5ukrTZhsfy1zX9Fdyf1n75ln3ja3THKc8aXoZz/BxGU1WcVb3lXOTlJOyd7WGxRrQSc
8hOaOPIhcDeNnIaiFjqpNuZPcz4QTHGwvCytAwQR19QfCPlSNaUk7ihKpAZBBh8ArkdTZe7jCHQg
4x39L8zzJuX7NIy6rNxPp4997xDpsII5VA4zasip2uj/OULgl4stxuLvYvfusFnZjgtsIke71ZRf
8vR6tzfqSO6fhuoWL8DjYNJk6VAKi5+FPOUbgXNRyIyJLiTubmEBKQY6f4wwvnpD4hs7hZ1L5A+O
fzTdS/vTuPHuE4l3Mfmi62hFdtpSHV8q02LJiIpMB2bYHcV6tpiIBel4puIY28HKc8jwyLcyCGA4
89EYRXUSrUwxsKRMjibi38W5KAPRXOwedr/vwTJ8f+PzZllW0gG6Y9Q5LRYa7JIwg9KBE+1zrwuy
z9PFh/kpPwcEVazLm63n87St7Fed9iLx+QkdWKwTBqqk46sUZP0GsW0YZyuYlDfs1LV1pG4r5u0Y
I4OiM82aU58XtVRHtaPZO1+7IIU1LG9MAgwBU+A/2fJNg6SMgUDoMVLBD7IFs7ESETttJDm0ae3c
erlVmcP3ohoANJIXDap9IWt/O1FCdmUV+N9DJWVnWQd5P/CmZSy+yikeX2Kn1+elyqFRvK+4I4Sk
9f84CYBoG7nk3tBMlNkvnRVNceK+js0ODqKHWTLpK0gu6IJNAIBLtJQUb/q9DK7Q88APbKM4UM3Q
W/CZUNeBsAJNJ6ItDrK1tfFZCipXOujJI++gm4Kftj4tZCkFnPZi0dBflHze2ocxexIH/It3QPw7
nvZX1AhrRjy8ib3gwfUf2MBqgNsuY3hq0PDUB/Zl7uxdUBzQ9URvNGjuYm17vXPjzCtg09/dsWO/
KMT1tOV2jzVPQKAozlNBBjKW+hCMFwxhfz24DXU+ZvUbOlK2uMX+G2bxfUqCbt0S6fNPKX9bmBg1
C9lNN+FaKFDC9MkVothScpoBfqXg+AvqjnjtdI7vrMl06SNy1xPgaAOX5C7AJhEw0YfCT9mgfMhz
h0liDMa7XoSkrXqxVGnBcSofaq/C9kD0q9xNCWOEO4gjyWnEUOj49BEIJ7L8zjPRMiBtKqBDs4/w
NS4gZSNrlDd7QnnL4uvB7efQjwYY2uS2wcSQhC8KTmQo08hSfsSlkhikajLR1BNPM27zg3Z3n0oA
i+u49UlntQbg1+kJt+jWKgrObMlmU0FYPw0Nmh1B/c+mQH1F9JI5i9f8h7nqfskuWEFRUoatAyck
wAgu0FsLuu2k4YFckZUPMgEcjlujxyIlDon4/q9hPKi7LcU/3NC6yDEa3XtwO/T/jLri0KmBrjSm
xXRcTi1nnsfzNJBp7Mcui5XOT6UX062oe9ij9KP1CI4XOH6B7lofwXkyy0rzy+1zbE6cPIWpzoKi
PWZcSoo4AiYTTV3PZIMEHe6AkaleOet9EN0nzaj8QOqotUAaOHFZc2379hAFAC1ZPDWm1CWpco8r
k7dthZnQoZDB6lLz0hbfYqD5WsKyfVFhej9Lu3C9tZru25NrdhCwmPEIiIXVvwIYqgejAD6ZuZn1
wrx4hzaorzyFQrb3zRiPYLEsJM4LBoVkA9KimsDeZvwwBgibZOTbnGFNpefFfncyRnWiZHOyX1c6
N/IcXEugGlEdmFwTVM8wZ2A2dKCMna5S3As1ZKBfiivhrjletZIJNbuvsUUD85amAdeNdgO48VoA
DWOkfM3qI+1aQre70uef2E+l7TYiqXTt6NSULnO8JA/SArlFly3DNgpRELVkIwYdLzJWLO/zsCqe
uPHJeu9D3KHh4UlVTqGrGVTedi94hxAVn2pjqe2gjTh+zIBetpYLHpEeudBfKCczrrSWQdZ6NM9N
eBebo7c2CyE4AhswWbsQvuafqjtnlVsADuBPJRgzZrS9MgoRd54UOYJyIQ/9UFNhPueCnvbRhyXe
xMaFg5ugUKOt5/gMEjSiveVCm4a2yEv60S0Niys+J5DRrt97GJQy5BXxfy2LFztZGfh1uqPQVrO4
6NiK4/+YGX9vwhv8Otbvo4/c7DBS1I68iwxk7ISAnEDDqBDPFGxzr6mc4/UNEIxxfIFdqQb/Snn+
SAaHmh/QJtd69B5BqBUJRzNGtm79rJYdaBrb+tgMWaqbM/g0mVqjGsqFUnX9Qg4Dcxa3QGxYymvg
9cdX1hqLdjr7bl2tWE/iVKbHc/GWS/a/NOBohvkJF3gAdblOrCnEvOmziVVP1YBjMD+myNZ9SXwT
vp349m1yzdkFc/3/WHImx3BK/ZdendVvG5fcvHqoiHftQvhzUpumNfTOHpZo7Mv8nKU0vDjI9bEG
iJKrSMlW+yNIwxNB0llZVhxn6khdYoiNLsKsmpFTYGuQns/lwLgxLg6ZIotj+EWD738Ou4HMdvZD
SQ6rwXesKlDopVmdoG7r16JmjBuJRRQnIkWFzhG6h3/ss4PCV9x2jq4sYevfad5KzMaORzVWN/Qd
rK0ugFoZ3+o6Zs++bDY3xyj1zY+d5oG+LG4zupxlBXmQv6ZojzGK7KMVY5cjfclKwg6dTwcvEXdw
mvIcZmpRIT009Hzl0Ab0q+Az6LmjFZHdC9ZLddVvJJ3J1i1gao0VR3onFWD7r2T2/KEZBytCIH0p
QUEad7wB3K3uQ6+fNV4al+CcfRJB7JkSwtbUBRGPmMmKVDVCq9IYi47+i5hlgRDS7n+VlUN/d4Gs
F462LYqlvPkIkLnIFJGknRW29PekG7HG5JCOaxMpDYTnmexC0j8Ut3d0+h+LjNtSlsPple40nKWT
t9STEoMeBq4MhmYllr515BdRIEOUI28gMW9K8GLN6iVjeVggatWMbtgxFvraOlxgKXIT01GZRXFd
4lNvCXa0CWOmOaFQZadRPspxAk4WrMcrGw2l3cu64h1szANV6cY8cA5RhfgLLoIFR9+cPKC85EMg
zYbUwbV77wVZlSiOBTHfti8VfPIq2JNPjl/bQ1iMzzU6MpWpRtfY5/iwF5pzGZfJFa9a+/jXwc9u
2INUeGG09Arz0+DYJHu+8r0ty/WpG4sZIJAehVaKhWavj36mo5pxIzFcquVa3mF84vjDlJp9v6+n
ARi/K6CI5VjNBQI5/0MWgYKM4aqQq1tZT2CsD4ta0kk2p7v+S3o2t7UuLWP+nazyagW+znRqcrEW
vsJRl/163kCKb3g77FoJ5TC0+MR4Bd8yrR7gzGAArSkQIOOELi23bjxJjVQAKqmVG1qmPFoEvbKo
emGOdUbaaA16WLKE7F9ZhBg09nGTAKdGZLIPrrkpykLLVaFpO6NtjFAyyVyOLMjd4gj451J5ODf/
zWC2lfxylgw9MwStFbKyOKWyKkOvvcm90vmf7bBj8tCqk1e8+k1Bop+GCZStIrAi+biyi7EqTfK2
B1V+vjXL1qfpyrI5IMrs8nryrLcb2Gm/laTqPBEC9/pkjcxTRs5kE/YAOM9IkLo/dBR/I2sqbOnc
oGLGTDlySuq4n0/MqCkqVR+7aCIuFC5B7osxk//iM1JkPHNUvXWalmhDIkupAowqCZarhGadCD35
pPqrTuW8rhEmKodBgqv6I0FwpNDawFVxdJj22lbVFWTFKjCEddIn5Q2LOyqvjvUIr7DZeY3Bzuug
jgrkEXc4ZuIv+JHEUgkZY0wFo0yYEI47svpLcgRK+HW/0llXXqE0+4MQCcw9aqwoRBbe7ZQE3bne
Rj6i6m/V/xWAJJ2q5nmSRZf4WB7FmtXpkdySXGSFms0B1LDHiAMXlW8ZUi8D1GYJRyf7ZS0FmHB5
ZS7aTM3lHk/d2o7l188Mb5oMndoutGhY9daWeMekMPj79nNwpDvvf0B1aeX/9j2uLjWhuV608iGV
YVCwKktOcetDNRh/tSJehrRGL/N7TMYEMYd+iJ2XEaEQFzg5SI7rMrMC9SKQQqLbUpNJl0OiwZB6
TT36w8ca6LOoISooiCjEof77+RoHrn2H03j6mo710GI51MrwDS5/tfSZdka0FOQ2cNisbOXGE8kj
LetfqLOVZ5P8nOI2QRtq3DfirDsGFz/EvriC4DI3gi5ZzNv0j9VDD2hZWG/pGqaKw3sbqNbaEvcF
KlOu4p1YcSXC/OPEHmjBkqsYGgoY8Mfvqr40AdpTghZVGC+fuLNOLswPvG0TtbTzFqT4kXXAnv21
kyLk3cuD93N1lPT+/jnfjl1a8x92dxGlxvW15buIUsvyBHO5gVUIKl/3Mix+icK6LeOikvBcK8cc
78kQxCCTfpwJ+vwD8UzYtsubcfca0veXEJkvlVpmZ5xeWv0iuPztlNzEBRutx/uDfdj4kptbHAnV
lzRY2+Vch1PtPL72DHbiJtzcHwNhKyUqJzkloLGpIvtCwI46DhImJSZKxTgyAxSGWrhys6H0ftIB
P9tywkR0VQjzecLn4g/8m1E3wg6k43ab7SGjq93sRgU7FU+gf8QTc3nbkLmh8rMnEs53xLkVeD+0
YNNd4PIoEWKrG0W2lzpJm1vSqtgOfMb48BIzWH+q8UAlQ4gSOyKod7RqyJobCJlgVyQO0p18OYBZ
8gCvNTLwlVZVltcTohZwqSKksm14jMIEssdmE/7DsZ829+bxsQSZhP284M6MgPpqZgr+2oPjSEP8
MkRhn9zpmgejSAcl1n3DfGWPU3uQNz7CFADZdm0Gj3+15APDK8auhZMss19aAbA+mHSkDeduAqQz
qQmZ5ZencsL77s78pGejdJrTfFeEn44LbQMYPlbw6vEGyYCgYA5VzJLVFubBF0lfehXUXssCWSrS
BVSX9vWSuxdJssU9LgScxHJbQ14RiKZO4pappcAdN6qtSqQ3O3VE4eRrTcGyhdJzbNNgPZZjpq5I
cTbdthTV6RICUNilhNMsz8lwpBuLqfwDRVzS8rmc0QdH4JPEM5rBjU6en2dXEVTgjbp2y6yDUmFR
xxs5HRSlvhTlut5gu6YLNmoJtse7VN39ZKxSYMpL9ArABnKXP9adK14uucrkvC0RQW9WbdusoBuA
eEIOCdq0dyze7NXVYfnFfqp6lS4kphhVzknKh9NBqLT0P3cg1fXLrYICC/hCwOgOqRUsKt4rb806
HF3ZvbRGHr6LBGfksQhakRrme62KV9xRI6e2c+3FAlB/Bg4Bv3wT+NVwTazFULzmvcDbWNOI87AI
KIVGEDZU+GiihqXwAHHDVbKNny27KyuUKO8BwTsAkLGgm5N/XbeYXFhxTTHXqKRqKu0XCFebCFdu
QrUNuSFhHCbmLTGAhfCFjnsJUTyt7KytzOhWsES2rk4YbML2UhyozEUXzP8+yHs35XU9aLrc8twg
chBnTILghxY9xaYIVRMv7sm3YF7TX2/+vQp6jPLOrtD6lJGZoMqGxE1vmQmDPCIBv7fi3ILvEmEy
hBwahcnJbVdF+Iy20O8Vmbe0iVgJ2kxAn6hriuuubuBpEPwCHjE976cyQyfE7WzMMsegLAJcPBqm
S4RswYkHzZ6Tc3EgPGG4MpAM2wo/2N5qZEuqA+1DpEpiHI0x0nC5gyv1g1oot+J6pqdG9c5TIkQ4
9mj5m6AAr9HDGDeX5NuEHq2BBQ1s864A7EcjjXO6yMK0H2ewqe3YsD9D1fnAsv66DYPzkR+NG17A
d4rmhUmkq0ezgUKtXxFibxz2pRbEQ2szPpkfeJDYJfs402LwLIsvqCE/Ltle27sIx3em818q+ZgY
FM1wKp7uBeR6bMbg1+Emc6QJoomC8fbB3ejpxjt5hhEMZ6y7wvqUzlCiQIF6wQxS6iK3xrRy0b1k
W62RdCwUCP5ZCTvxWeWGohVKRNjgPA6kImD2V/RsoiM3m/Fjhugmv2oRGJy5ihOImQXjwLqPlepa
hpj6J6UJSs9JgidxZBhGEg4x281h84U7NHoKFgabiEpOQQfsso/wsXIM2jRzHtTVTLiyORrFLoId
5zmFafwoWzJ8gUPowRBuEnNt1KX/beg74pJDY2En8mGs/EJwexK5CMdzeKCmbhfp95NVlQTU8rea
FV3i9IRQrixFgsXGq7uRGYMsHzI2oUQF6jj/yfSQwTAepy0hwZy/WfcsZEW6yAV6imFMgPPgeiKv
m/Uw64aWo9f9q/5mGrwNiM3mHmxQ/h8Dz+HAbqTJPHsHw0gjkJMTLeRCCrLFxvzpn+rxoVrn0gn2
78jRpT0emL4/zapql3F0175crC2O0DGqk+YxWx2rYZVx381gS89lFDSmqw/hq7T+W5NTXJATFPOT
q5sEuLfXh2w1kSP+xxe2dH2JdLMPNFJSHSKi5AFVP2ZSU8zzMJHLcRo/jMiD9nEayEYdXapEslH8
8CaW1DBVh9yTr3N3X4ZLWkIGGa+whfuJcukrIHN0dd9/Onsr9XeX3aKFhBb++WYwIjJPILo1m49X
xBG7ixi8QLgN7Y8KnZlS14Ri7KvP5XMk4CvmZeVOgcQspBFy3Zl95EYsqJVLNASS1O70KMPscnJb
BXLnaBnM9ce49L7MCI0VZHaJORNsL+mJSSLyS1E7Ga+8vNNiwucrStAxylHeTyBxe5HFFoDllbHV
EqMS5TUkg/4UawZ0rPQYxzFeaLOFghc57I+vS4LMJCMk0U+AkXt9btjmqfyub3NLAcDxJmiJ+ZZE
TzRPp0enpuZITmz1fRw5vApnObaOO7OsHUHvjVBgWTSxBfmK7Vpx0wmO5oSXVCuXgLPerpl1oYbj
gH2JMrSeARD/+7yyvoquspOvqiz01KId/9q6MEG7RHovqZEp3Y+VyUGwq7DcDdFcU4cLYSkRbIe4
2XabpduRhstPcXAOfoJ6HkJmuRlEi8QT0zWvhxfdSn5ZuScdG0tOpMC0vvYL9eoEdcKKbOAy0Yhg
18t4rOWY4kl/7UEx49rK7cfZhsDhexqfF63yUsdg5jUHh9tXSzxly9hWjuMpnwkb7ZTgcaZFlh4E
F17YGJQGG5QW3r9klJRnIdGaFFIPmRUblJfV8rj+IyZgLy5zUnl5HjgaAD2NLOQWAx2OyinkYRkm
9LnXofERpxjubsBaKeRxNzJKgIW9ZwLtR7Z7rW+0nuh2wmfInig7DBDf6TxgccQ/DxC3alHvrSbt
FOpHl5zeKajJk10/3VFuzCdNUptHZ8LTzNwZ/+mbeH12yrgqyRcIyGvjjCB9DG4ujbmpBlXQjcJ4
KWH2g0gZ+cKOFc5T+obn660HE01VvxWDGYKsrN+aW81BMLUyFX2WpZaNTno71DaK72zx3nVMFhnZ
z2hvau0h4EXt8n4koGHACW4pheuxKrEd9xUsxilmtJU1bjL0GdhZvW/vgQrcxbIYFUWtGluIg01f
4jUYuSa+HJRm0jlkvzsOBSLWl/EdQLyzJYRxB4XTXyPQObUDJph2W/Kq20aE8+dI8uSMSRumrWae
BWUYTb8safDT8d4/qh1EecHl3wJUmIhsXwCGin7AL6cz3uhEv4tut/ikP0cnt8EiGTC6G6cv9qCE
VGXQtQKSLicLPzY/+I2jJTEGvO01GwNHDZA5RsZn/aOC21jk8eFufXGvsfjVMoQIcJto+8PyeBpr
NnhYUm0qwHrN1WRtmqnvSSSRhXGLWp/Sh9XOWe22eEAlIEYLqoQLepHpLwv24JTQ6Cpr5XvqvXcu
Le8GogvlP2Ew/J0mgzXrcxVLAh29lR06Bov5ovFIAYWTaYrUEhqRcOYHzp0jBI9UzAbQtx4kMPLO
lOU07Z1hkZUt57gDe9w/BTqTKGPYAw9OxkDMAOG9DdM7Q0vyA8HqOLC6NZCqB+4RfPv96Zd6x5vp
V/kiOHxKtY96sEpJTupXQjZniydNibFT6MlCX4cHdY6bVhrmxBxworP/ss9BkzDSqa6yzFz1b0Er
MaLiwgFlwPJi1mg1i5VLOV5HKEztgtm4id0A5ZQLw80zlTxo1kuIB4hgriR3JN8KBB3FsLk+RQPP
amuIBKxXKhHR+RMYFkGObkhxY5cwPoE9R5snOOacYtyP7xTbXkdaqYQZ06pmaMQouAUz8QLm2JPG
PSv5jSqlUM/GW8QQladxyt+HVMa55/kE1pJLDD6VK9M5AZXFzfyJGa1Zi48+4rxYQnl93A54aG2O
VIPO3y/yw/IkPaYeLTBa4/RlbuzNhGQEOGAn40MHOqU5OgIFXEQS0e9rKng/A7VG6JE4Wcl7kmj7
yiv0LkP0gEZbZJKqO/buWDVEfpWcQ4jOcj0RuXUWTBJVuDwTOgaUQUkud65dRZUguhOEBlKDwP2c
M1SL+tuTptiix9W0u0YUPqtvLIsCJE7hqhLsWGXwrWjtwobjrtN1r6iLcIfO6cM+UTmVO3LKh03G
sI+PNIgvbdaCYMSOA4xWO5b2ztT/kSF+Pbd9v4Udiy6CXunHYoT/Wiam//TzoibzSSnHNPrv6oZV
jc5HNB7yWIyRUDruI4VtA3cknLuLBTDXqgmjbO3J2uYFnBGltvewlTLfqEqNKVdoggrfs6c0TKl/
9cesg38OwiZ46dIinsKEkaiONbLIRy++h1GR9i8OTc+QnlkxgIZgq9817Bkho/Zlp2Io5lNGSNRS
iosbGSmj15EA/03oC2cbHqnHL5cALmeYaHGtQbfLbrZlcOvitqpuHwubPK3rpzTkCbPfhJH/UUNM
QfjsdX+4NuSq8NSbcznk6WfhHYYfyq7Ax5KEzAPXMF46995zZ7Qyrp1VY5mP+R5DYnYxMNBkmkl8
tH8Ya/XlCQQUqQPJowAQmRO8lTAgf9WyQfb9f6cigTkDo5L4qbH+ZNKBskyQ7c+K0baPTqkyNj6o
9ATLwbRKv7BoCNC2hOnsZTiZT++A43JMkTJXiNSYibUB0rl3rpx47eN+tvo+tlgtc6dBRXkSlboZ
lMCx2z/HGw5dpi5m96Q/aJfK8HC1PtM53ME90nXQ4mEdmjUkD5z76SmhCGv3zRvGoae6IMhz+Zka
87B0n/tiidsEvBsKD4j82GJOeUYnWFcm+gg8LM8u+F7NMNzyq662fo/beqO7rhQOD9j/MZm7s+Gt
J7bQJpRnlSFipOgXEot4mc3l0d5iu4FErYwRn2uqlTTdMKc+liz9UZK2Iu1ocbObRRs4OPJDh0Bh
jvPJUA5DJ02fL0adJA7IXsyATC/jnG6Hl/P3kOdL3Ftu2v1MSZWRAVjkPs94we3LXINsdxqKU0Vh
UDJOMGzc48sYd6Qh9STSu5ZT/a/Af9+mrgunI4z4NWfSAfCyQ0kJfQP9cIrzoZb2Lp2yMbo+Wn/F
COp/ag3NTVed0rC8yZ6esdhA0vBg1Vqmo7lU0GZTKJvXmPBcJ1jZ8fBA1iStGmgy3XJ38owuAE04
u26h8JPZPMdBXPPFgLgfE65d5bsghRHZUAC4zC1ARCMGqK+aMvABunJ/ODnXlIAcrmnPIGT0h989
kdI2peB7+op1wy9hJn59BTu1wvrGepRcCgIeZ1RZbao2tk26XMCumOX+ix0Cn/8ynhBR16B1LbH+
963/tFF7NrjhNvprOrlpM8kf0JKqjnFLFbIKYIU3fdbJmHYhcvLEaPIleu8eHlkVwB2lPxcFFqpN
+sSQSdPF0TCuiUM/sGCVdujvxr2R0M5qqCGlkIbGz2VvOx5mAbC2sLHfYHdtfZqO0soEJJJpkhMW
GHInTnDd/EsCLdgHA3+oA4lgwkLh2qiezb4Dama5lbUaw94bFnWMPFgmZlmJUoYe+Iub49aBVJyM
LQ6Sr9T/8QDxA5tAbr9vmqA6AbyVRPdooowxGzXzDQmd3IwtVZnfSFEotsshjkVFAdrx1eUbVrFI
vaQXTzu0ag4XsSeoq88Uz/0KDRU6LW4fCgbczk+9wtIV48sUA33N0Cyipqvbaf3fVI1BgSa60mFr
/Q2AP5Qh40Czd6+uRo4WUfciMdGueumFymV/U9Li4gtpkunS7IXBO5Hb8VhKw91k7CzQIKhz02nP
BUvqIgfzEfhwsv9lmyGw7h/BNXpcw1dEZ1PnbVKc94nSd5pSvItWdPQWtRXnqdPKw7U+OiUsHPVo
iPtbXRZliy8R9ZDN7/asr6XB6bvbraQBv+RcPjM+vV5kLYnbcr9CtcFUlka9IemTXo9s+F5HBVnN
m2bkbbgky8G+kopsZdmBGBX5ZoGJDmgQeTX4T6BWrjAzMLh2Ikv9oT8s/81ysmoFOFZy71HbeeRJ
XQKQUjk33bXHD0W922ZQNdFUC7KxsjNVscutXwx27uV566G2dlWcECFc/T7HSSWDWwFG5VS/xzkJ
ORqbcz9wkHN1palde7Q35mbBnmQA56QqvQinpgRsByxKVWbSAMh+ToUs5y6GJasIaWgsvHLHijGS
NX4C19H5RJfN13qDH0ZvN4b1RK3VuHmIO098Ht6CYiw1vO+E67oJs0XS95dVtEUEiq8Gi+NTGlEc
EqKRyQ2vh3NM5Tg28GfDuWxD1JsX0hlQScafpKkxfZIZ4zittuheBUxQEwSXUbbhoxIW1EIpqfDc
Ld0e8uYDUqrRInzXPqJqpXG7n06EPmHsRPb8iSDW+glr3SmFr4O6YKL7YL3gMTlav8ULzrv2rVFG
PUoI3pyTpwEWqEDVS9AmloigiYRfJ+B+t+A9Kqji5oO85J1uLeTYjuyEvwbAM13nMGu3c5R4nKF8
vkGVz5IVnjLLeEdCJnXDOFyDJPrvvGZy+uG/e5ZsOamv7r0xaV0frkbQNu+h+ApY8BzPxRyZim9+
YpZSD9Vih4VeiMuuCYySwhep36Aih2mVJFtNBaMf05IT8dTz+vSXpWJfA1thEtZ+yTFB9R42RdFt
vn1RiUGjeGL/t4d3mWw0EaSz9z78tWR4lvVoP6UUDKtiBAJ5JATX/lEfYU2Lpfl04keccKVQMqA7
+RgcPOAq8DVKAV2iuHtbjExs6hXutUCx+08Snqe0HipAhbOdYRLvvz6nxvlcbCNCOOYfZo2baAqK
l/G2nZFwVtWOPa/oBpJybAla49S+gZdoQ5Wtv+82fOTOwiELINHdZUVktM8hiX0j7hTu5pYVJqLP
M5DkCG4KidhqVXraSE3qcoHXml9WFBHY5qJcmgm65WvGNkl41EkjpamKHULeTvUAQCW77B2qyxYX
an9ZuU8OLcseK5Z7yTWUZh6rwAJcc4KM9hMkGhLpJi3ml06JCKUhCCU7FDFxEIz/xynMOb1GyVz9
Xv7/Fy7deoL5m66YhIvrinnuU7HL91iqF+ze6pPRJC7hTpT5V558jZDiODNphxihYGZcZIfjOYHB
2+J5sYsMFbjlAT0tt9ithwOK6Cgn0NMTqEhGz3IUcvn0480QEuIjt9OIFc0UO5yAAwLlH12WvLmZ
nq8BnEIyw+eePqMaabbxgUAsfiKaTJKoeqVxbsLEfsMG+BOM9sH5FoXqb0YOmnYnp12mvSo/hi4N
WVLpm/RjMIsAUlunCAMZgNb8IneJ8x9WRmM+ruGnFrSLZPk6wQUCxvAU9oLW5HAGMvMYGLhZSBBE
mee6CcF6+Z4o+phNQt0FJnhzfq0zUzQ5HDhcg0U8hb0uOIAWTT+6QCqcUFGPy2AsGzp2op4Teu66
4iDYsVwrH3X2V/B7oe5a4+HBUTEq8LGnMcvuQITTZbbTduJETNxdNg5EVYUfAhDCWQJyIcx9F7A5
lLkVHsXxfyEkJFnPZe5xqW6AHLt8t1hcd/hTh9RVv/1mP5liLSGY3qKoh4/lKL//i1CWjoM5I7hs
yif5t8QAKeX7e9bH4SZuIZIdVQ9fWi55FT0Mi8u9E24PhZxBPLENOOzkucgcYWs2YHMykPd3am1C
aJu5+C7dbdU21iEeAa2u32JAkds40hvmy6gGb48BJ9FLvGa2c+ge0sjNvIkrnx91SnQcAnS6n2AC
kyCZYn6s/cRVJVrU1Nk64r5qgHqNmnXESzLw9XcfLIE9GDds2UU/yAJZly5ADoSl/pNGIa1J1CM7
2MTeFOiXj7NimVtsr+93frKamKvjvXSfBeDYURQjXaL3Gk0m08K7ly1btbbIrq4K8b3SMUDVx5f/
dfQgvyHEqfTEo/BnM+9/pZJTc9ekmABirTI+/ZTQHyd65Q4nCkal62mbjK1XXSaSPLxMiSpVoHuY
hsUaPUXAU/iu5eqzBVgyt/tl1qIF7UV4hnjtYXT6U1tAiQ6YqR+40WwGJAOgKlsuuxgeSX56W1hR
CQarJOUeDtRXdzraQD+xa0MOvEWLQQq99oQFLa5Z/LoZF4j5vUeezx4m0QuHTv2WtcCr0/io+QLa
OMs504kQs6VaqewgCjjA0vwhUU0yS5oryD+d+t4fEBHOLMB4zWhhf505eAVZLgqnc92lBzhU51Qm
P8/NLybYSwXGaAY0n6MfikoMNy4CdXnPxzawgt8CkvmFZv2Dwf9udmzCfqvmM/GTFG0zhq9w4GvW
q9xE1MqjomHshuCCEWMOlsqz1kfnSsq48HxeJA+wZykp1aRNBAqaoZd6yJOr8uo288QttavHhbdM
Z4uIrbLYwlFdBu00cCxuLDRoZyo7Z7lDp1KWnPi4hzFvbHBBvj7JwDhZhE224LmpzAAok8+sk2EF
kc5FTFkaDuKmHIFVzb/LJck6UJctRrYEGFr0GuaYAqofZR2utdck2q3A6sF4tUDiejRmZt9tHQY9
kvi5xvXcJwAJXA22z9yiytwAVg9nCDrktuuWWr/HuLeCXA/VDz+NsSZV+78jgRgXnxy1eNJOTZvv
GIZLS4C6hC7eQpXxD7MzTLZAuWQCk3y4czvDXmms2Lom3OU7fZzLy9WP6VOfZpIV8nDQYMGc8oJo
N2C8r0V+N8Oa7LPZlLIXdsWS19qZmYyyvBQFc9BIW4H10reMPqVli9sSAzz6g32H4EpSWEmtljl0
sVRYBtOalgvfmsSPDz+YNbQYr77MxrI8SEpaKJ2WphchT3Z3Nk4fDdECqlxHsUduQxzOEp5AXW6h
ZkfAukR0Zp/7/DwlZTJGYaJOtnPkGFnO74R4h/n/puWgSQsUKcBEa1GZjqq/dp3z5WHQQQMpkr/U
Y+XSqb5k9n0eyRkw03lsQiRafPJaQubL1eN9o1e5mD8ZFw1YA961PSM+G17d5QIvEqxMVlEq0Dbk
SxD5S+SGPYMY4tNBGbW5m9W/LgZC2HznDbKC4n1SduvBWgBTBN/uv/3BUUsP/8C2RPBbnjwupMTd
wY/VuiqHqgLYCdnIWFpNFrMkRxJo4KgOA5xmJM3IiCVhZJkS/CYprq8kzAaWWvG2ikdqhfpyEQYv
0IHsSMsLCT+npVf8VybRweOpAk7JWro5NMFy/rJiTySykoEyFWAJWavbw3ASTVYk5e0tOy/hj35E
VDCFjBg0VmwRr/MWSCz5mwsMWloQ14zXp/WXkES8Swc7ZbasKj1eWymPIudsSqYRcTLkf/GpRQnT
MgwoUjcp4m6/SaVElu869Gke0ll9ED/1EZJ/okFC4QBrEx5BBvBhLDq1DAqJoHZ3MxRf7xPB7ME4
6YLU8nbo93bwhtx0voFfq2VOvL/6K+/4MXKEAgUDcyOILm5ZWn1KE2ot0+BeTAKy+gx0ZIfuPpoT
bqZfTqYrbegXI49W4AOQRq1I5XmkObzvxdUku3U1pd8AiWvT/CwcpnlPTrQQeMKzoq5Jyd2ItxFl
aE4RiTiy3ktgezP0ACy2psTHAth+kDSYCc5/Nao2TQ0GEQji/7j/TAFCD/IAevG+TnRX6KtMgGhK
TCwoaiaWk9Ibwm1ZLSmgxYQZhFbBB63LSqKDuaLSzapja36Yu+T9xO854/nN0FQGu9TLIgiXSE2W
HVgHNoOPeevLCrSOaXpoge08hL3ncs3tY737vuPngA8T7f4Czw2y+/3uA84qXo/Ty7aYb5VuQQnE
v6Vj9KiQlHnubKhbTvSLNp75vDn9axA79Oh64R65kpHljGktxq/onwTBvqNkJDWXwXZ+YFwsjv4N
9kdAhmDmckc0mn6n6za/uSrutDv2nAKO3a+s4oi5LhHJZzMkYi3wRH5zGiERtydmuaYo7nUKTDXk
aS6Zqu6PrQF1Zx+TEeB2YHxTXZPdEXXCC81Zl/tUHveNkWiMMrAxY0M6i7k6NWNy60NCsmEerZIC
ioBu80hqsKoXs7IS3Bp/ChvELFzicqNYT70lizayO8HC6nSn/yRXIkCCRD7G+QmiinNUbOWN+1lR
UbfU8zUBjJe8y7SNei4zA93etYjVOnCS64YT6nQ2sypwEOhKwlvuLoZ4IrdjDhuH26fLRlJhaea+
Ou+az4Q//fPL+XwIwnd3xcO2RPc14gc70WUOewbBguiFbPhrjn3ugRe/UJMv79ePYNVcgIFrVd2P
HiGRadkdUFfrAi3E91L3zHIplmCbTtXUUCGI4gmv8+UEt1OeyNaV/TP/gZa4hKxvB/3+aklTUOFd
Obt+jZSddcvvzjCj2hLvStMFM7qIxku7BqUpQd2S7Rdlh+RJg8UqeZrHxZC6F3282yhjgF8MHcAM
8uYwHZ027NVWhmHeq/4PT8H9ox4Qk/XZ0WFtmTMquT8G2Gp9y+RYez2hfdZK30CDK4Ysx7iK+wS+
My9oqoitQUhRzu4BxgmzaEnencnEKUHd2QlMDIbGRHGFCHO+PqDHD4iVy8hmU03Qebu3pN/vmmqN
OKpnLFbGn7pnCtwbAj/j9hoPeCuHTL+RLGQYNSU7ifl4o64ZqSPAm7e4EcO+CSuHmSMKbgLpiWk8
fBlS0yullS/+iosNG4CRKUVAkRbdOzc8SevJm3DD5l8Yr+fsgU+k3YkN33iQdGyHBh8j+Mi5H80o
C0MB9drChuK/4VHadHdHo59tu1NQoLzUAXwUbl2EhYIKK921vrclVNB1HnS1rf3enJsWXSC8SvwX
/snzdMsOn+e0IXOXJXeueyeF4Q8LBwPXWkHRMrIuFT7a79193ag4USAEfhuYNNTstBFudnpsF/aQ
Hnq0DVZ8gJ1a0QX9QpYFuUOYg69vdU8UCbZofH/4SNttAoWIt/VIn2SnfgnpDmDyuWneRlObj0GK
mwyDt43YPJY3RcMUOXquDxmZnrFBJnuXfnsvM93YRQbf2sjHhmdVC3ltCe2YpRTGYNpnX/M//ADn
bTETbk9pOjr5KrKCNOXSm3sWJ4tWYlvAo5xT7KZ9sXQKqma51cIhLmsvIbZE+XoKoK1+0jPisMDd
2tzbZgIyk1hrQsmtygZ3N6LXTQywKjPQnMGUiidTPWc8bo//iZNp7KmGjwo+oL7ixGK1yg9FzyT3
wBGlWcfxWM4nk+0nVwTu56B3n8ND1VtIDnzyNfpoAmWzvKzChYg09owj8liauYP2cPQo3je2tXgl
e9EtXwjUWCfuDcreHjhYyAfwEiFr80lMXmeLsGbd2cs26YIcJvV0Nly5KdvYB2RUXQxsscJMpJRo
Op94IiAH41QDZIvNLTEouicwhO5V8FMH56dAc854+BBdfXo50lIy4qr4jXA5Paqs1dRCMM65p+yn
lZ4fJFWBVuzuH1Q9zE6jsZ12Uqm3CDWcEP9Bj6YeI0aTe/59JussnjD+zg7OoojuxG6TlNH63KhP
a8G/BYc36nYptVdgHIZ8Y02fDYqfQy88pl0IcSCKIP5vZGTduerCj1EvSOOZesIZLokycDhWE8TS
Gu3XvLSX/JRB+kI8D6+uZYCH7LuKoqk4xtl7hHqMYEtTd5XesQg/vSo2sbt378CQInNTNEcJfyuP
VRX9vN2y0zDz84dHc1p+25PXVgEN/Vuktb7uViF6BguqsFwlTbm7JpIgapA95Ylh3xpe6KRi6KfA
hfpAyNVhbFVUzBQ2yjVHaSHNPQBDfp7X8h8IwbqH1hvyGNrxp4xzRvcIIxVbe5fyMVwckfr54tcL
Z/kCh84PKSxZ8G2jOHkLhpT9SJ0RHn140PvrTjZ4nobJDO2ZJ9RWHeNmHSffXAHYcXkaFVuwZE07
m9ryXLiOKIa9blBRuC2/sk6c2bBwF4hS12qiuaZNRzEPlLgfj4sTdDQsnrxaoLPmnvSCv1Qub6Hz
LBZRHxYiJO4JfVQWvn7XNrAq4CYZ7l+z/tTa76/4FYkIAZ+aRFLd9X1oMEBbO+ugt4Q4ZX88e31K
+Vo05lPIl44nPjQaM9ckLXxOtqL1yFNnLErsdC77bV53lWxhPcuM6Njd3mw246tEHt/6GDlA/WDz
6Glc08x3k/kvf7hHaJfd8AhVud/Sz03ft4oxzL3xU76nRYGbMOsj36DAXKz9Hw5xRt+9zGwwVtNj
BA+RZw0oUjN2AAwNHwysG3bSPyOWfTnh/r/IaB5H7hFo6SJ1jdZNV6amhvL1ci2OBO4szpmJdQRd
SNKV4lQ0OPgvG81KGM6UCsWswdzJJZN8xO/0H2fJWIRjvdDw27rlgc0H/lLUuIgGuJirp1Lk1y+y
PHFsxnalEJpFcZz2Fz+Gh3LDOlWW+PTopr04iTcEfz01l3ZadnHrVXJYFQUq2TCAl42HgvXPkHbn
f7YUkaXhZ/9zo6igqtiutvFBh3w6ADYOW6+2fnH4jJ5AH7z3xz0ZY6Kr/Km5/T3ChWtAZJ+xdPX+
V9CX8O5qRnvmMu0sniXykOzjgSWeTNacLWKW2193Kof2ydpNeqqgNZ2iX6GwPppjpVn+JChR0qPU
BtgH4/gELAOoaKWJsUmwWNoGxmJLNuN9QGYVgR0syuahJjcrVvxl/R+SMOYJIOY2c5826oUA+aiJ
V2mbYP+nuvP7agLLMkZqIbxhBTD1cbfCMPGVicDC7Ib5XaSIWJ88O0XBIMa0kDILstwbmQ4pDhNP
wCiKvEjaJPhP81AEsqA1Sdn/pAhxsPmlN/xvZPvRDuMfdaUnNg8WyCEIVH/1RsdVLGiiSmXxjakh
zn+fBTqmPgo6COyCfMU3MqnzmDhhqLvqr+FH14YvMuj/xOHXUkug61pXYAZeQFFwT1Cw5yutnpMo
POP1E6UMeoiyqsbcO3XUItT8A/kzVhdMbAH9tPoex+JbufSBXDc+i5WaX5kAzbYLnhHS9zMgIVxa
uCGYOf1DfPbdZO5HFdBJPK+/zvj/PPIJAIxmDBe9sZv5EMJsClJI+lSbSDsrPbWvYgPmffGQknlM
XndvR8sWlylg+sEiEu7J13WojM/wgzhMRecvbgn9AY0S8T8HpoM0Na2BXQD9/DaMtN5uN+rsf9Dd
RFdxk8jIXmju156c0Ya0vzHgAsD5hAKNh7SBB/LP/cnvcQQ81lk7h2t9r3ojnMpva2h0/DrtI1Ge
PLXyawpFsP5UytRwnNENdfqarR8xInZ9ia+Z9ad546uxcnHiYkRMzQFXKtbzeSa7fmBylEYd5mDi
rwj5njB9rOo6dOH64qTZiJlFRPyK/ODScqGCGGOrNlG6w43gMJ5fZ9TsuzT/D4Ir0b9Zz+lZqlIQ
v1rpD+o78DXPyF9wq33rm/w+PjeBsP38b2jeCoAy3HtD1pw25+F0L09xD8YlStyLpp762ZQ1vhV8
rWM9wvkbcSf9B+5KgoksqzSuYyUot6YXhSJflGylcRbAt5xDJW5SseN+MtNWTdjB3vaZ0khWNYeA
RKgfV+0X47nazngVU7rwjpqpVxLhl2G4rxVAV3wvjwFQuulVzdNS1MQ7Fsw7uG+UnZOC/qcWqB5J
NBOmz7EkYVbthJII3ajRS0DZ03lt9SGC17q8+Kf5VOXDrCNTJcf8AJYndvMzMqK+x4blRNiwbjus
SdECe4hIlkYKSxRw2RX69BNsYEPyDUs4ct8C345oqh7MX0CQ6ld9c+x9Lgp4fqoCh9jidqg0CZVU
3+1qm+dsi2tVzuZDL6Of61tlyVOWcYxAVjHS09dleeH+RN6xGdHUMXLhtNIOVmg9dw+cS3aJXgDx
aKycf3KdpWrS85gyU7QZYuAYTirMSC+URuLmcrSDsiHVs0zx/xmA2fvVWcA4ZotowE8xYWNJFr6m
tGaYkIMvYZ6NfeygBYt4Ed+dYFlxManSlXt0R4UE+OMte4rHzw0hUIpQL23uso3gCEu3/f9tpY9E
+ElRXzJW700yz8MaPncrrZ+YXa5YqQ9N4y5+gKQMO2WNhOgfM5hyQLOhNXjRyhAplKvFFTCRKOBG
Apg9cUoRLVYv/OZHkIClb/2cgP8gmB/2i9kCY8pnPMgEtVahqE4QTKDXjvLrh2VzLcfKb5fLZCgc
paHCzcil1W4sGh46Ee9497acdTXW2fJR2n0IU4zmGoOWQplCLyqLZYtX1OpJKJn/wqGnprhi0cFc
5xnu9Rcdec6NgxRhPHjiItVUy+vXHkhJWNEdcneFCkzGqMzMG3cbYUKHzE7p90kIfH/423Jet3i3
FO6g7zjja6O+iveK6e0Ao1OUWdKkd84iNWWwUf7c0M8jG4y16/Sxph6QJYQm0Sl6I6rUljDrYXGr
ztYUsasFazspEZPST09yw2U+rtnxdXVVSdhOH+dURjCEa384D8hnzHFZfJ5vOL9jY6wjPTAMnWrq
xVt882uXdD+9SwFcG/1dAbdhgkcu57FXozgqgPMIXfiUhnXf9tVmQQgL5Mf9oPAjXSf21N91wtgx
/O+j2HLIwPTW/s9rSboHaKZYGFqbyGpFJYd0umEfO72u/tF90pbiU2WILPVsEFtOPHUfadzoeUT9
M+GhYdP8zLJXjMfh+/HYd1k/aMk1py61oR/LBf7ASUxS3Vl6NLIALsUHCo4mF5EAoaFHFSHzEKH+
DbXqqofQMVxbzk0BeWQUereuM0185p7G+Ql32I1s6hSbJTQJKZtoUXYhfTo9g1inrg7vgeW7Rhq7
7yoyUopEI/BJ5ueYUSy7KpesYkp96/QGriejK9rpBsOEpJgV7uFw4gqJArZ7rDNhdcHTZz8rd8Ql
Hf/DwJ0xlF4CJYvyaqeEc/hLxTqEPsHUqHLI8y5uoQWi35QRQX/aF9BiM9Fxxsezc4Liv5m42S6H
GinxgthBZKGEHBF+DrxHAnVPlpSuHhP9uzAqzyhuemqNdMQdYLXW9qVf1Rl5oAhC3BRLcHY9D/An
VBbBUGTie13m/g/qpuxzVaM3Munuqc+0ptEpeyiHCMXaoF55LPCZ2qQKbE/XaCVt4X/HidUzZy3E
KwRZp+0vhopoSj/ilLHO3lcRWSdpc0vU+7qHkOgYyz/bAvBT5jhV4HvfUY+HeL0y/0PuUSrIoMuJ
feASxo9TwxUuFHwtzeZ1nolonPzqaSuzUsp1kv8ZU/XP9bHayXL8Bv6vbAiqMpfb43SjuS1C5c3P
Ep3Wo7Y/aRuKvL2P91yXG39oq64av20SLW4VRO5dSunHYHEPfQbFh1/bMJsghhWRrMX9+kEsS4HT
rcPlJHUoqWRZX4QWCXKlWNrVbWDKX2G21BrXxuj+M79J6LGuwpsjsXoSpLyLALATJ2NAPIGEt2n+
2kEZEiMrRy1c179NbyUVrWU6z0jFKOjIJrYO2rJKdo+5luQJLsUCAoiSX4r7F8j/ORlaau4+3QLq
AMkfplN1lr5K+rNHnIuUmMdNFqs+lJQDGTbSEzma5pGOf51OTVxImvVZIe1hI0WTkLynk4OGOtQi
xcJ/fyAWilfm8sKWJF9Tpw6BgzcWEdJwOTBC3gNQvdzDE3t/vCSk3JTwEUb7ycrWvWSUFKUCbZ9f
LnpCzWJ2Oh/zojNwXLGVoYonunPMj043Oy5J4gLbaY3pFH4u7xTj+E3pE3Ul0V6AdoSOjpHnjhtl
ufORtPIzXm6NwxU1hgKfS5f7z1HzJwf7lO06Yr6ZgZHb3wzW2AGPMLQMvQ+UHuy9pNFtZn9hxD6I
7sRvwBIGxzLJ1cHF/apYuDFLgKzKEjSuF8KEerlYkhD35KiVFwZrtc5S5glhhLq0/dYAmkQyCgCS
AdZetdXa078nm4o2Z8mAD95n/MqdrR8UK+vyQtU23yRDCvu/qpIMp3G6YBBmNiV6Uc1gOJ2CGv8T
ZUb7fQjJFN4iRz7u2PdWblgD5KUWBybIan6mZWsrz1uGydt4fjXDnbTMt88U/BeRSvNQklSOv2cD
nxF5xX/0gSVEY236mFwngnncNv5sCo8hJq9s0o0Z+idqwsdj5Wsi9flZcvMFTirswPHAvIx+48lo
8V4AyeRdfg8udN3jtBlJDwCJ07z0Hdc3iPodj4MHTLvQHggrry0sAHy2o2vEA1CXgjQp4QdaaJAO
jqB2PR8VzlDIPTLt9xx6HqWIhl2ALhHwSITd6vNRoPXoGBwAsKmKrC0GkRTGvIRnHoLn/i1yrYaJ
RjwySB7qUxdqy/uvV4EeRccx204wmqThhi4YbNCvfHZZ6g3cW8Bg66ZcjifYWKW0lXXFktI6BCih
yz14TpXRWSbbECVSxjZhYSdGyjiEeGMARTilKsI/LRL6o06iieYqUeTrkskKYODMUenPxL0jKIRw
Uq0OzWFukM7WcelaDaHlIT1fhmasBbuuQBzwxFbGYG8B6x8yhy5GDB59vH7I1fGrZGiJakEPl5xw
rWKiRC2apWbUVpZ0ajmgvAujTAI5bmo+o04kFhkl7TFoiYR08Eb6Rh2ArYsaX/iHnThmoE3ipqsR
XJoLRVpIGJ4WkLP2W503BwMtPDrDEb4jK924buqwHztaBpFVwo0K2gunjcm0IKX1LT6v8lfPosb8
sEs7d4G+KTci/NSwsEAvcA5Ul8X1tUoCsGx6YHozsIR7MkfJlydkeG7DJ+igHktFImiBhe6V+8IQ
c0P4zY+ZtCQ6F/FeCYzfUW4G+fWNkmt61Xcv3fkjZXQ/c2rvsDZFIpUNkFfvs4sHkLJhvBsI21jj
ir5A0KL0katrIpNxrJMg6OHqiodMd9gHABIEzfYheL8iCm9Huyr4X4Vyh7Xm/ra7zu6y/a2I080l
1OEwevFOp4Zgi6oTFRNn5r2msO3h2DdXDZf/ReauY3Arq5fGxpMQsf5IpskxjasmNG2hWGi+MxfI
oU7DT7VAqeYnfYZcNGN563C3m1RbaaeM4I2o39+OQ+hRpbOn8hCgXZQNA9yBEtCabeDmApcjs4A/
KomlVaxrJCL4UqxiT9pq3gqv4PtEV9nc3u5t6xZFZSd4CnvzjDY0AhdScNILwKxUm1fFaoJrmeve
RoNi6qlbruzIvn/Mt3jq/PMIuwETPCnwUlV45c2AODlBET2XlavURqZafr8cjgFLw2fuB7LNBamM
6SGpvxTIgh0JRFrA5XqqV93OdGyM8ZHQstUspaCas5brzn31THxUgUXEiJ6R0gD1RVz4KEAbB+DV
DiIjqTVLnyLqvuo5/Uvb4GgCgLlj6uV8wKRAzNm+NH3ZHSO0iJwEnLK2SN12JUaDm2YAbSsXF+Q9
C/dGS+ehJKMn37zUA/VDLsbyNDCMXmD940bnleD84u9qvnEzNkrlzXz1Wu2zpi2OdhmSHdkzN8Vj
pa5FsuxjOoTsFfLKZ3yzGHv724i6kGyKjp0Maiw6kj4O5USwuUsdreQpByXt92oOcggB0WtBkKnK
FxXbEnlGlqjZ4TSirmW4xDehnUTABSIvngP/z63XorY+iaIZKqKB0LdfZi9EFT/yWP+ECWEmIwU1
GwQg2ZIZrxDackbNgLXFd+9e+bcjCZj9yYIK8eZp6TGcgdmItH+npf8KNcfJfOdTjOqk/QMgIfHZ
hAIpKwFQg9sn0NKnkZKasbFKhP0tJIBDamUOUvrFVVJt8IMx95HQ9VZkTVH/B/uA0avUq2Kpqrz5
2a8bHU/rgH7VKpazKzI/fCKOmwKsG+Tnv5Nq7jkS4LTMtWRODym5HUKybMJgcT6CVLX7xVCNCv62
TNIs7ZG1iZ6xZAEBWXIxIw5GVYYgJAP0RICDyFbwFOG9P5Yls8CMk/++pP0RaJp/VF2T2+J3TXIp
+vrTqQRW7q76Tm+8SWP961QLa5GNBEm2kcExZJ8nz0lon1E4FDptqHPgwcsHrLiak9rfHh/vqcQo
TfzeoOWJFkvQQtn0T6IXy3AgAQm30e0uqiSFCJ4gSl6FYDeDnKGgUrxtoYkeRCrgJYLHQG7N7jc8
crGscy8PqyUzhU8lLL9J3DTb6dh3Tihs58L87HFp611XcKj0VvmnyqyNT2XMVEk5PZNRM3gsaaXu
guS7vzZ4lF+85Jbcg92NtQFm3GWVit00+6VAzKVKqFm6g+aC44zD5UaH5fLkTCzV0hv8NrsnrMki
cUeKcLH2YXlzWDnyvEWp6b5VC/j+eggoqGr83r2lfH/hRwfrwOp4xRhjGCxsw3zZfusyjTmMW5Lu
ERRB1iGhwGxc3+ks6u1FGuEcj4N0aRBef6OxhWTGVj8zjPasmmCi88ReFN6MIN7pUZqIDdd2NtwU
YmZ3QGjKTH1BCJEW0p1n2TD6ESflI+orluNap1/JJFRuLvU8F92HKY7ZV1ekx70hwbtYDf8lToKp
95A0pbizcdpkNI3fisuBLGXvhzlXRuFd0xPMLdGdLnKM6XofBSEIgpPlWPh2sy+IJF5kg78+4yAx
UGt9Xv2tsAZOeJx/vZzMaFR1v9jIrvBz2rfOF/g2CgwyQJpy107U/1TMVXLc5cX7ZR2WMI5gMv0C
nRNKD30sP02oqszSWKy/jNo1WaKweP8lBOccLhfmKkymaWXhyT2keNuA1uUeULUsV6LXMNBpj50p
VxQgQnhe/CJPOnVQqWVFmCH0FLHZN5MjVvTY7GqJbKO4riEtl2Y6YDSSjvPJdlbJP0B8byaCYN0O
3m72kJUmtbCrHgYGijAhWz9aWkEA6Yve7Vp+IrY/MgqmZ6Cs7F/RiTKextXIFuW25kCS5O1e6fwz
EVRCtbHh0xO8PH09cXejhkXTXr1OjIR2AiI1MnSGUKyxJPbilJIybp66uAzfbG1lTWvezlh5CIHI
NFyOWQrRvhr+w8azMddLLtk1AO+R/B1vJ8xTsLNEjS5IAF4lVjKu3Ugt+/DUBIjaPm+Jhgo6eA06
ilxRZRZ74l27rqIvQPk8R45p/6+kyYEGsu6Kx9yfdiFxlv5xR1AR3Mq7t0SgMUiBcic5lJs1yWuA
DdCHzteLtUiAyjSrofuGzzqYYm383ySUYGFe4QwhySoxzzy3hFQeYYIpZzkStgEQ+cdF6GfaYIL3
3qgBZ0HsPqbuKBiowvRByBoI6+GVifMfEf5ODlpxqaEXCgo+hYLZwTJj/4XZL9VxK8mEstdn7bX+
65CJWri+Y6/qTY4Hxt8V/FDJYiJsptOF7hBV23N0FKTJDGp6lpG9xjDz+vRSq6D+N65VwOAOpyF2
8mBKnxjef8V2PbqVQiRI5jCEeG6hBEBtjzx9rBXRRgilIT32ikt9/nQA+c/iZ84CPbApoFoy9roe
6LeRJBtLJfReldvPUknWCcz33k5qtpC3Mm1HQsYZSLJiGXYX6B2QmveHAjnjPOHN+yGxndBPh3ob
KIBl42ChRJB4HIrktMnBQaLfXlck9CjOPe+6kzXYe7Toyb2scdbVpb/X45Tamxqp/XMrlsqeuXBR
H2qzDu6J6Jp148EWTS1qTDOfWEz5ctGVdpX3iTJ1CNDfAVdXQKMCLQky1AIZlO9lY3dRJmSGBZ93
ey/ycR63OaVhc1fbVpZiGmc8MoOfd6U//fbAKDgcAwfin03dx+b1WdfLpyaR3A6vCCOC+rbD0Eoz
Efpxb9NVQVjwFYbTW1h+NAIS63gTDfkzfYAzpdtws7TOn36up+gwsRYTYDyphLdQb0yI61Lme/vB
gMlWS1DR1omgtLSnnOErZJyYNM5a+CZ80FTTQkKjicMvb3C0ry8/Kf80toV7RzXupxQ4MzjFk7r0
sNaGUo0+wpZ8drjrf6ZauLYYfHeypybcsG/S8wSh525Sd30jQmPUzPMg+lxoKTp7TjnRb5cBA8Mn
2GOFQvMhKq5Hpxd5x//NXxWhkZv0Sf4LBPzzrmrGw0EbpQPNsNI2l3ZrXn2lyhG5wpp3fhBZkvqT
EuEq2E+1Go2So2CsOUN8kIGqDk/FY83/BhBFq3rLTuZqpBjQQqA8NPKnnpu/79rEcGO4ka14sIzS
xeC3tlYdmx7h/3SgrIehep6iRZBXG75rIkvv4NFHgpNwwHopBE7ZiRFRJ01KJyyJTL4V3KHmwFvY
dTS6zfefyXp9KV0MEJD4WIexXmk1BTc5fMq+0MB7N8DnDiUXhdC0Cl4LhQfZMTbtO0/SwUVz28aj
cHs7Bf26Xx7FNrh0IrFAjtQceyaiX3iJu5Wb4LVUZVI6HJz2+rdaeZbJQ4fjL8bqp43LKEn/6IPi
L/+nZ77Ytg8Bq+YkViyeqla+TdGyIV+ztaaREzHzhYqpAO+NvGjnsbzOqk9w5wr6zhgYDcFIreyb
NEilRqqTMYgX/SIHiVcCQvvcin9DWFoZomCk9p/DUIOFVxvVuZnaIBPbjFkzR3+Is4youQxKwm7W
eGd+p1RVbZL8UFJIdihBfQTournXqGR1NjZ2tVn3lIFFPM6RBwo6YL2gQlMY+5DW0CR0ilp3CIeb
LbP3cqDjBOpYZsvkzzW2Un3AUiF9bMNA9JeHd1kTiaYbidWQU+JA832mJi3WJ+bEdT+DvVHqn/sR
LKnr22wmyTlNZaTjtqgyHKIGghWizQ9OX87G3e0Y8yvcAXsN1BkmsaO2AalTw2CfaHUBiMF0Vcob
4Jf7vcWiWIGBGn0pVYWfQftYOALUTzAyEJmHX0FU3XGEgcOmoVLozAJfybl43AOcRkwqd/0yvdQ5
Kx/7k7yXm5JiocwGZvJaO0/Tx4kbhxuEU1L5qRBUKgzU2rnzNfT0HlXizOIfqN1OJ/P+89yAwUGQ
XC4TyTUQB7dQFM7bhAdGsitfemZFcehFIojvUfIMAZ+ha2We4AtX0JNIZH8dct+6bYWZ7J7vmeJ4
q8ifbbmA0wjyencYnRtisimq/jfBAA1zodMB98LZOXFkFDZaZW+PpIg3AarZ5YbvU0+m3KbUzKR3
4vvdk0nexVjNHMe1ov6mZf1Ypv0xix+2bs8ZbWsva8lOPO9zTnKt+nab4cfFoHC/QxZuejD2mY9E
v0hO6XvsYvgYXY8w/QdrrfvECpFJxMnSAOZAOIvGAi0t78P7xgvjVe+A3+sHr2igJl4/Fh6x7P5h
njlDf7VDywvZ9yvIY/hvEZLerY1LIpDajO0n+gxWl2Ij76q4IbPDAD6kC0FPHjKUpoi/b8MYE7cX
8G0Kzo7ml7Dg0qrD0G3qGXjbBR0IjtTOCOrtJNdB6wSdi7SDNUo3gJUcfCBT5Uck61ZQkjCJY8td
v4Wl68fgbYFahDqXmFEmwANY7NLhKcqpOdTk7MV9ahhl+5n3cVgngvC8mqvdxWdo0Px0Li3WVzov
cYKnhtfYDU7V38ZtKZZTUuY2CNGO4+W9WK1+4OW7Egt0k3NGl6cE1XOlYSTZ/iWFSqiMUpltKg0T
Jzc+DrD+ou0HfyrP4z0+Wl7ZrcqP5XOgkW9roMJJ3H9kr4LYzwgTK1jVs/wPtBySwyhmFONY99o4
BSR7hzy+4bOPMy4lSvLeg8p4il6gyF1vfQG4/jlhw0m7pWqwXpGLKYrI+w6n1S17RwMeBdPUZQjX
kN52BxaoYt9fyGBhZFqgtzMrR3x5+/pJ8Esgr7A2VscequxPy9ve0pRWqo7IIGGdZRwtT7MiKwgT
Xr8CJPCUJRY9DWaWTjC+d1G8ty6HzarVC7gNqiiWyzQA+mkl/rwEHrdzcUsO7YOC9VIgiXTL5VEO
bH1ocJYTNOIc7mYl0n7VIlLIHX/lxcd/U4MPIq7aQOwVEZOvCTW16/W/EJkZsjO0UcJPr/XKwkIm
dyHA3iGoz5hLhQ5AVyV7Re2ajwwvOa0iCS5lx9a7aCP6DA4H0pK0O4pNE0jVpTzRDwRb8Nu8dJzA
2Yp73HtYiLwwPb2UEEmcozm0NKrL0AEDA8+x2CLM+RMM0+wI/9omTPmYlXhb77Djm2pMzJwtSEc9
V/jauxXB2mid/zEAukdBdkjdQMlWpUpY+essSok+GMZTjr2TzqyBrZj3NbuZCXGEGnJqUgu7Jzdh
qh1h8KpyGYd9PtBQNtyf7YAch22ShJon4K+FhOUfdpNfijFY8iaKiKG+mrqJjQlNu1t/PxBJcC8Y
jE4dNCyl3LYHZ40voNa8OKswqxz+A1K/CCZz+JTV2jOO92KsCj1tGS88OdaxJ4sqhgi0x2+OXdWc
2TzGh9cYmCuRlItt4M0U41qhZLgWr3GP0IPGYFpcKKFowo3PCBUUNOzW6k4VkCwc+mdmN04oft2Y
9feSDhLbx6C4VaOVZ9peKv4H9yWpQw4+EoT4jJez9GyZwaaeFBpFrtV0H5QyN8odN3fR/vnTn6BH
muhZmhZd8RA9ODpYDlXNFK62xmATWWbH26qrlcE2ugW8OZGTWWoZvrXRDeqKaoHGRfQ0t1VYtJHC
/qAq9Ctjdq0M15BTMK319sdOYCoCH0nuL/awCEl4jw28Q3YxPAsDNKP6fEjdvnUNBkKZD50y73Jq
vbnAFaaRsF2bGFZ99YdNs+UeSZqHOVt5bUiHgMZ4yDs4vIF4U0d2Q3CFBeyX4g0N5iLpkbw0SiAe
TzfoKpVFDfONtd/KoW3JF4MR96qjVe1mygJ2nhgPBQy/fqXpkmhcF8rciuqhPn4SH8PPDhz/giSZ
L5DgO4zyHMlUipkw/VuVqah70EfcWGTHEpG/GIAzzYpY0brgHG2X1EmYV8oFQburPKBZ7ffUv0Qx
GqfaubHORMnPjJBn4avqVT3Bv62bdFHO+fhCZ/8ujbvfr0dKS1dUOhYWTpPbyQFD5aDL4K9PBvBd
jCO6Zo+xmqf7xOri6ACsgkMXH4rjvYvp/TugBg70tyBJh4SeweK3i9gBPmvyr7DuG4gKeWv4/KFh
2bCodreAAg7ZzBeMurUTdztq3jhGAQA+agksPFtYVQ3Opx9x/FxXWdaXbGCbthg16ogPkXVvHBfp
Zx5jnY3zl5bgcf+cKvxaZ/kJgtnUay608zcHLTQSodj/aU1XkUnLjfSMhkDnZ4ayS9VdsN21Hnze
6oC4nFDeeCp181C5j3QgawJ1rxXuUEpHyGsqYdnp9frK+6ElgOVzDfjEc8iR8vOkcutKR62LDvBQ
GedxlCKf9S6O18wycEePuK4azu/VOVrVfo9A8UdzvttFIzYImpTPzsGKyDtv6xhQof+gvLi9LYai
NHEhSilK2+VMqEj1hazMrTyfMKKzldRebxY9cPHTakLA+tlC42mUiNA+Vpo0BiPTV3RjBUSnW35l
0Nn+0gtdo2o3dfLZEixv03bn4fQ6C/3cIla+PSHxK3ryyffvYzrrfrIjYUP3/jQIWQlyvJ3TBFYE
itI2SsF+dCU1JIzT07Gvi3kCtFMBIp638U9NM/UzcmOgtZrRZiYxtQfNdpd/bHhH1v7jIC5tnIjJ
WSWB0BtelBEWIbwMe3UZz0x1kCYtRo0RJTE294JRHhd9oQNC9zDjZzu9ngOhxicqtEFvtdex2gLk
5JcoNZ1A/iEQuPZ9rPfyVS1XdBkX72Pav5zRdTLu2SiM9ug4Ewq60IhbuwzeLQgnhiSA761i9FuO
xZAcNpxdBrxX3yafuDh37RsmKHiFEH7GXk55Odhj6uRYZheAO+Vzz9Kk2PpuOqQ9jeZ85Ces/CTJ
78E6HQbFNS3H0qVNk597PuYiGadELaVvTOTc5SR6UzquQuzsH8Us93gK5q61g1YMFjwOcRj1Vt0C
4K5OZCHjwRrQ6n9IxQtKRkRYTV9cYMfBNQsi/qIhtwIHwbr7SenZ5jTwwF8+NhnWIWDf2VKWHVi4
RDOa9HyasNGzg5f02r4BsXwFkBcgGgkT79xgo9fk5OBvmrwdvbCvq7NDmIpQeeZ+SZDUkOV4KjcS
VoQR1Zp7XUEozoXFpA9FdppP6AXicuU57pZyZvNAAxk0defOyQjnP97B1NEh/+4jVkCAfspnEn7O
B3/6Leejtmmou3NjB0tfFCwMH8KDZ6MCKh3pD6RM1+rkloLdQs+aA4LqjlEdRTbgX1itVtDQ6fdI
iKXZ26zYpj7T2ouXK6JepCG2QsLvfDuGwtNRsJcsoCeWULllRBzNqFaiJHkCI8uHiK/zssjHOjnJ
TwIxHfEgShqSF4B1Acqg47PAc2h/E5GXy0PFf5yw/Z2+vZTFnznonmpjAYOlY1r9DWlwt6BqnEw3
wVJ3A9dYvslkjsStGzAGBX2sYayHUmLp03srU0bxfsBwtE6QskyOcO6wjoY+k2bwyCOanuFbSdNc
vglQTUz6NRLg33SF8rzS+J78sf07KszGQtRs1I+Kt16WJnpgPC5BZD7ZVjiEPr4sxARvr2d+W+Ne
fAjp83/NaDFZZF/F3yjE8AKigyq0J3DkmMw9CD9tHFjWc2Ukj7nHlieL99XaUS2a4MJGzAO9FKqY
sY3AevPw2p3iHRr7uKJ9CRbscO8LyLNcbGfqvFRHeDwHwjY5YoMg24vyQqMWN3qmGrhB2/y5q4Nj
B3QVLN1R12GpL0G6+RQbYbMdM8KdPUM/MtPHhRK88hMCvI6pNbyaOaeUHUxd3m4YIjtfHn9x00eC
SDToHO1xahzYRwuP8jLLjA8a02o/A5ukBMyo8yKFIrXgb0k/FG1oCoPLXHWSZhkGoGcYmQIPwfLa
PurKppQUOnc693tukx82pQlDLlO7udO0oMewjM9ywXMPrE3WVQyPQ0Jwpdh2uaxs+fACFX2FC0iu
YF6q1yGMSUED5gJ67MsYtdY98+vFgQ6vpcxE5iajpmmg4UGDbI9wgRsfsBZHnYKRozwkcPfww4Nd
QA+jn3b2N54RvDmHxeYNXbGSB8ZPyKzzTNp3z8UbP37K/4rPZhgZJ8HMbLASLpiGrNciNUYyWZ2p
WvaVugaF/wAbmkybkz+d3bqeuJSVUVa/47pDmltkqm/D1eonx0Q8jw4jrx1+Cs4xOyXxjb+9/BR0
7ywTKkjSCN6yxfoVermyAsWXK0OkZgEL0UEQ7D6JgasxpTZweEAbMBTqLzWlMWqaYhKpmvhwaQPC
zjZgvUZwgwR73j5neOn9V5xKmPTH9p9Q8uSfmfSMWrKtO8TCzqWIoT6VER44mr9/LzsdABUbXdJN
33ARUNsAGC0jTF6xetIWCqCq5wMOmnFhy++8Eh/BMZxRkcl/8X9Hga0cIdzGjc4jcjpLecJKb1SR
pP3+66LD/gsI2hv103y/yvnngaAr1zQqGf0onkr5EGCdhnVpHM2FjDBcNC7cP1SPC+Xg+qJXjIxn
AuA//RoemlhvQeRHN8WZaJELA/GUJaB/VglJ1E91iZGdLqC6uzTxM+f8cjA9AJHQOniD89w5Ddjl
u80hWWdYR4/ISadN62gAuszM3PgsZWxtJ7W5cCFkKNnzN+pH3ZtENmfhBHMzBzw70lSjBN2NzMtn
zVXFlmeDoP12SfwhfhlNRiyW4QLTXnEb9zqTXVgXyb/UbKuQNYkeRrvBfmp6WiPPwrIGXJHfWS5y
fAYanODvR2gYEEUwaNEZQXP+VBirzPBLj0hNtQXZT+fMQR5JYEK4nmDtb4BV90IP3i2/yHPc3ip+
VDBTAjH/7zqg1MaXEBhuyjUF4HmfwkLHvYvB36AHH/0UBjI97tYjaHmzoaCtikTeXyxtd73bTLCv
cCe6s0cb2aropIgRJQn100jaiwO9MsP0K4zUpt7ra0PewGFm3YP7P77nysX8eLuz7MHdozcupaxl
n+yuh/azOHgw9rDBgQizLI43pRGWIOt0TZzwa08yUXbEBWDw/2cXI6SE/j+iGvrXMlHb0Nk6asRJ
j+t6wGQMjtmQAD+9NHar7oAUP0unDXvROZVO80NvQKrTYozRxGYxnPawj0v0Dy9IECXCr6Vf4QKs
w2Z8UvGfGMJkc+JCPBHxEOoAONSZGto2lFS4UmcTDvnAE77LPz/0xbXu+W72JI5LV0vEuMaSg986
s0WBDtbYTtT7AmeodOegvFlvClSZ+SnLR/O0dcYHbpAYAkL8oc6AQNeGduul3sWMcPRG8G0XMIx+
m7byfNmkYi6PSzw9iUa0E4ivOuCf+0PRay5R/L5urJp3bUvN+hnrH5V6mT/6GSVj+oVKY8lIOFSz
NPTE5Gq/3ZlXExVHDBEF8tUrvwTHUKV/EafaTNc0cg/wZHu+yucOfRaZJ+FnU9OeJtMLKkRUo7xh
QBksYEd1nkwasBTYs6q5eZ2tLdEBzi+daN+aT7Zgf/6SroNTc83Ev0Ifiyv8FBVlPCI54SfUiyEM
Zu572AZHHVIUXROwTA2t8d8AnIx+asMVhKB5Sb3JuzYL96+UQZcYXUZfPOjGh6CAsqYqgRfHZZvs
yBR1IUJ4RQaNJe+q8vqBirqSHhha0vkLrFmu3I1yUMwYJOPxw6mbaedhWUT01q1YHY/7wEZGuxAi
uqt4MXQCevP31zRoofuZL5U+BoBaBuKoxeVj2WecwNUOMzI3qXwCIo6ppOj22oSLVzESXkmgU4jH
B7oZ2ulTPd/8a9YT0ZFsZprR9Ln1RfKCQpHC0jN48RwdRehzcBklM0CTHBWzceZU8lJv9fAhP2B6
RciQEzEtpkB9+UrPGFiMqehPM7RDSe0irCPxa8x0KPmJ/hZYox/pMc/ymF0aIRtUOZTH68OegPsV
UMyRJa1TXm+glNOQv0UGKYAdJ1ZKmZJqRDEBO2wcYHFI/UPpoYHKtR8fpzCxujFATyl1DRMFz7Jr
LZE7x2/zFy2NEL14pp5rpSxfxgPRGfZh+ZMzem5CZRWWR0AlwUdeATqMFAdkBrt5w2tHDPxk2pA0
v3cMFNwRiFBj/J7LRXkMc7TN9taxzUxeDGfOu866NB5rWTN9qGlL5KrOQfGrYQMLpgCjBXN57ty0
1A4+aJYP8M+GAi8gxtyNuV5g40fw+g/qBIR338ekaisIWWWctpR0CULYjdJxtgjq5Akq0Z2rTgSJ
WBN0GJi7VoYjFypCjwFwhDBGvVvvKAcuvmclsQyUd1zyTz2SmpP5TyAM9FQpg4mCjlcNLAx8z6ZO
i8A4y5TmyuT3vZibe3n+5f9GD6oB6+x2IiDV8VdWRl+Lk4vZ8mDvJUSsS+hQRbb9UqWdWQjVvLQ3
fyZdPapjk1ktFnVqnMRkwoUGq8vBMNG8xAS8CJnANOHO+kyR1rA3xRvWtdblGn8aNQsC18u2mmIW
DXMxz56KKdt5S/5PK7Hw+SWo727LBkINNU5i/EuE/Icfe/wjFc2uRPI4ZPo+Sz7EN6nzg9UjUqji
iPFkiz3hOwR+dpHNUeZiPIY+lklOQA9xEALjZ3ipSm+1HQMYaXvBWyIu6oFOEjmA/rj8jJ7TzQKb
6RjGSTZqLNvuBESu2WMd29KubAHpCvLiRY35ng6DZrBPrxvZtjhvml+e3cy/VdYvBPUUOTpdbodi
RWMapftD8QpyuCwBQ7vrzhk/aROD7PyXnlk7kySAEzcx7y5pPR3ES3MMHRzsmoIBWYwMgrLzOs73
D7IJ4CMlqNQCnCahFumg0A9Ic3To3xQnuqTdEOzUX9VRp64agnUExsQq+AN8IeBBN67Y4sutZlZK
+eqGZdainIW/b81QH0WAm6PFhW42o2ZZZTqzTHxSCZCaJjyb+vIZpOOx391RshRPWJ/16hSJbcog
yf7EjpQZjdf1fT1nvAGtce1MXUseBTRx7gnR4UMvkXVr2f1CN037sxE58W/idpEGjdp80LdPJJBq
2kgUlB5FNG1FB3ldFTKsP7ULD+QvOKIE/iVB1zn8uTOE3VLqN5RuinobzzHlUwXcI0xcZtPzzo88
Ro7qLGUH3V1KzsHLICROjmObeAqVQ2ZrKZxERAi4osq+Zjjcd4YcsNEkmycjcV5/PjoEEdCrTykr
8pudALbWzuVGqVgPAhd5cz+sJBI6ei8zTypjSkBklADfa5AryCzXTYlXUhY6SLiko0GA5vp15iyI
ZsuvNFE4896iGaRqU/Xcb2yqsoj6dAtdrSxRrd2zk2dHnuAI3PVzZkulE676+sBbk7QKwyFgd/eb
bd0B+HsXqlc/yxi6RijXfYTFVKkMbu2c7EKyhFDEQKIrEwRZ7eXgkN4zb1HeLDG6vWeW4e3t2U/X
Q3wZ4yrnb4WwH63ULzF0CkAo6Que+pdoYU6jBlKTm984OO3NOre69Sujqn9cz9StZwBWRu3UJOxt
uV6k+Guda94cYDAIj+YI+5qiNqt8QACEDiObOuqs5OGJWQDgyq5k5YBxMw/SpXflrpM9A4/HEyxK
iNPFA1e/ecADl/43M75G8iFH00N7GM7Gh2h9F0d+1XOvRXd+MsNMeZpRRQrl9U6pFPuYIWm2OWkm
xvfVkurZfHDmKPb0wzxJ/C7GzhLEUGMWqQVlgqtSMwJpS8sCY1G9pUlOzYoQlRcHIVOvvMoTx0YM
PBOKM4l3kobj365sTs5hPstL/pCdwUV1/occ07TBDTcgBTTowD00ADOVgo+1SCNo6M/5gakGdvfJ
97VNER+BZINbCVYSLJkizU3c/J0HXgXoSv5uTd/5oxZdZ2ZQsKJzzw3nAfskkniABCmPZ4FxJi59
3NKBurXGGXZWoWw920ZheN917Kn4avHm3kYDRt1Lap6upANlzFTGAmX3yWqBXhKsV4gO5NuBW0eT
tXevgDFZ2lhd8QUjdhA3UpU7PsfrwXLOaXnjFOU8dr7jf19bpbjBTk/ruM/Xs/ui7e2kGPCn9suC
nRy401pcPBAVNR0H/BiITz8fcv3FlfL13np6H/yo4+eZbaGl8bmA2b832ip2Vi+/dWpiNHhZ8ibN
d1lVQ2lsq3PePEDT0EkEJc+lF6Lsg7ZQiVzrWgV24rdpjBKPqd/yFKJnzokAbGmOBhSXcZ/insv7
rtVOogy23SUTRddCIWmC/DpE9CT6+zLT2HLDjv+rTWr3IN3jBfRZgU5uwXUE3rimxQnLPVlQ/9Qo
gTlt3eFy8t8LChm4awhEJlRhI+VFoujanMwvyHXJz7tBYXHZWNb88FOXkkHB+KJ6n6ZemhiTOm6b
IxqeB9wqC+DY6/DJE6OuFMnrQ8glVV03i/Z5wDpawKg8EaXQn4eC6Q1+WwqWpAvSR+QoWuX53QZ2
8dXkhIF7r8LvgQiv6gpRxB+VBCulYyrmhav1L5aIsXmSv9n7d7EMOsqfghadmdQkmwkBKU0mvw1X
1gxJZWEJKuk7NwixAGUOPQpkuVmb4obaWNaLXLyHINhFNrub0F8IYKLkuj+yejz+TElgijT0LWvR
WciMoSVgBhSETyc2hQ5muGjtvWZdEXiVl4PQUHtWtInjbNONle6NfmgE14nWCCcwZEHfVGYBMaG3
Ml/zUtkYKVSnzF+YAWqTDzTEaqyDYyFcNglc36a5XCbo1Hv1naXevBjWhgU3yUxAgfTfxpFKn68D
CDbpLdKyolLgGC5IS3TVk2w/J2Qzq6VCEAvNp025XYicGB31VPeDcxh1SbXtEQJXesHRM7GDCPH3
e3ZPwLLE7kHkSZqI2EuD/pvh+4Gl1uMe8HZMWHb3MsAKOWwfIbTiorvWarFf9fG41Fr8O0HA4hfQ
alMYK5KseoKXmhv20aZxTs2x0VOr20shLfUjbwMakeHC6IrtLL/MXyzNri84uDo2ehx4NlLejROg
EPw41aUwbHo00b0iS+AF/35XSycx5tQ3liJF6664USk7yD8+81hW+H5bDB6KD3Q5A8ixS87nXnLl
BcTsAR2/rqXl6dUVIau05+rZ3eH37lGZe3DiHtrlrrXC2AJLc4rjRceI+JQu7ZREadRNOXQAVCvz
3Wy5pBt7md4fb6DNUfkJQwt9J6F1vaF6poyeocCxdIGC2s6WPgQUWt4Q3X68jC8+DgEU39Fk5axr
s5/l/Xk1qyaJ9NbHXokv5VXi8PDT3GO+jeJeet/yxopAjMIi7w8VMOB6NbBTutDcHxeW49I5Y3hR
sCNukzgxeJ3Ni5S/S1/8BdFS2pUPETcGkonNHlMI80R3K//d3dAePpqZFVB4wfeKsIA2KzVpmLvw
ghT1c3fHNwzyIvD0YA3rWkz6647iyP3GQRum7jGbDNa8o3S1Xv+edB729g1LinPx0RxKQNBeVh/I
VJVMu2j3EM1i9ZKMPyxPuS7yOfgIU0opsodL53jTAphoZV11GRSqgDoTDvxYreLaHSzRXq2nkwYC
KytPkQYYyiUycNMWlNEAub9vCPcZSwIH+4EYB/f7VfpdQETwycR/Q4ttyL0y0TpG1l4FY0onTaBe
M5rA/zTasfrVVMBHXTu5nmU5ZI8On2FYxHLwQGKs0+8DxseErmquQvohkknHRLJTUz8JkyTrXcR6
3Yq/1zeDX6s65oSAjlKiOHxDqswUyKXfaJtYkl4W7VS7wD02Z0+/tGzuTbM2F6fh5wzSGuxAneuh
6Pwo7G7lUVUDBORm3m7ITI1CGkqBWtV9hUL/UDo3/NUrGF0X7eoBk3oxMEVG7c80zLJj7sxJt1Ue
7hq1Lyzvv31bVZsln5ZOdNNSwifXDsH8C81VR/TgJAISX6p8+O7FJldsBRcfvU7v2/rDd2h15CVQ
yWtLUPlsSOA3P1BE2MjKYBnxkfBQ/LlDPVWTzH/RR0i9+vfU4Zi+t/KZE/yuoOSUp3SrQP9IitXp
dyfsqCaDtcwMPs2yS9sFOkV0z7JyacDK/7tgpeqJr5/1/nkC807/KgvQhMb/LDPowqsd2rlnHYAB
OvKC0ouwJD0qhw14QPPFtipl9IrWDX4dI4StJFcUyC4oMnS2TzBFGe1Y1SmDCVKxy2OGBlHBsM4U
htMGF/NwBOoCL5iVmmpggNwM+xhwlbcZEstfS0Pq9pxuZ43imxqiDU+PkMs+qtJtg22Tq8ed327G
6QH8/q6+54JvbgxuApM8/i3O3k/vii4zvEjZV08Faz+lNZ+WJ4xoNEjO1RM8xAvlqPxLBJDZwjZ9
PfkcbWcdISiqs8aUSdUT+CQg/dWV9K7pjXtDzV8zxyW+uG2VwhSKFe0en9sbeoI2WvZ5cjAPSnWd
Aeho3EaRiOuYi4vqiODlef7L22M2FybsSpBGUJtNCrrCtTnHvDvpYZMpxkbhT6ahRaihtfugN0+0
scWqJYnPBKTU+FybKu8LubFkiWRpzyTp59ilqPVcdBGEYY4w6YLkkFu/f/z9W3mQ0i9bFeYWbIbh
nV4XuExjqA7SqoEz9Kk8AbQtPNTfV5uhIWyYlnl3O6a/6KYkAskrvQ4/ELUl+cOh4g4y6UoDuCxk
D0YxOQUXZ5YGce29Z/eXMSGmg8NO+o+5pvkYWCZQc1IvQMg1bZkDmB6OYPhNQnTovcG3pj3E56S5
iw3Q8oSNOJ4Slj/UrklxiMZm9ATEJeOOdMLMB3D7aGB3k+nNonzkwh9ZWL7gkvQ/SLMl36rdEIna
wpLbukunIiN80uvs5Yoz4JlmNlqQFPCtc5jjZcqPXerBa2Ugb07K13p4eUcn0QayGIR7C6+DTbp6
Fh0caUKOTaQETXJCNnJeyIJjUN2NUkBe0u3ZVqgkaUyI6SZMkynXDeYv2XzGnk6oZMJjc5TLaAPC
Ylfbcq1qZL+TtB+8MMb85Ng3xrQ5hSq6meYXLfX0B//uOVtLyf2agEvrFrLVYf/B4SDoVmoVU/DG
J72oxnu7HDr3yAplA97UslBE5WrvzVEtjQmH4Q86w+jTcBxAG+bYfnFNXlnanm3EUasPVh2DUZs7
Ju/Wj0NyAIW5IvDWZ0CIqZJlA7xetzDVtOfMnOEnCJ8JflPVWiIZ/LyR3oFPLjEEFXN6j3TwEBcj
OYhyz9TXZSl6llSV3kQElGesgId7a+rMnZJpu1ODPyFZxCEZXg2fGxqBTAnhE9JGwyUH8qi0ora6
v6MXPl5Bif8/hRyoLku42j5UqMuXFswzSAWRoNxecBuW0onNncZoLdTNs77IOne4xhdv6xpB8Vpi
QAebsjMFsh59oJMToa6Iyvmlz5XhwbmZmbZhb9IuxBtWmLcTcRXwUi/4rzWU6rQPgKv3aaNAUvVK
pVZx3dqmXRgomhM39UK3jEN9D0OT95p1AiyS3pSqLYfjnHyMrk5djoNzCCNLdfYYX9bHFi/Sr7ML
wa1H4S1bCXJS7j1K3lVgtp/5+SoIFsIVZ1j2mcIWSQ335q/12GxSnUFE0cIgFNeDKwIGDO48xM/9
yKTs1yRx8axhgaFo/pNNV+3ljLqwWOrWpT8OxDS+TWiI4Fpw1z2up7Y3kdHHGbysekA7p4K+CWyP
+aP3YrTr/qFkgXJPXOJwMykG72/X+T+nqlEUkQ1UP1BDtB81Lbr+5QbjB2V1wxf7fToIg2ZoLfgf
mnB1VXK47jsaf+xNPPIKV8K/MD4q5rZ9WYzTtBqGBbP+S9jyNSQIlRDEmGet7MKXrj6Tn/ek9XJj
0sPsFDSFr+Lp2O+74og5UCsQCT15LVWybbcxOulP/yXWj/k4lTDf44/tarYXAmn2dTW11M4EUczI
Y61j5KpMjf3jpJy7NfwGi9dW9thx9dOBByShVZV4WdIIHmy8QxizsBt61QZFpWB6wY3oyzMV3XUg
tDJRYfYT2QiKOLQzrEdQH5PxAPM3eamXGxX1uOvJZiCB26IpWwycWck7tzGqW9eSxF7Ep+gADoJX
HIYR9iDN7D1ER2ATZpoRuuOhxVqK7fk2zGO3Jc/THyx/+XNGLNKVlkf87XvuG2qVs680vJRT8m3J
rKrzN+6D3nQlr0x7NDOGiqbNMjKPwbSfSQ5NZ8CyQrlGg/Ljm2arMMgoH3Odkx7MZdTYrLuKWGX0
3u1IcGQlnTb8GExasLz2r215RV5dKgfNI2z6Y10sjmJuAvrKyFdAjy9JU/j8xP4ei5JZ6/Jb4TZ0
Z8PZM06IVNmVhwCJRPMxGxvG9kzKWgoe5rWG4CUvVaN7x0f/oHu2OqjL2TanOqz8SsE2M0maOwJ5
aOGLq3Nuz8cJN8XFnd76DOcujQIGzj291Tve8R1gCC8F81XJ868VGy3Q36KcTpoLiz1uJ2M7crOU
t/OlwJRN5UwHO8t5nC2Lv2e0xLjTRB3ocWgDec+3+BgcnrolQb0cwATQGB8XHt063GpN4kA9sXoy
0Ct8/0/5QkVnlfI1WvOyfwOceKFE8PEPrQNfdod8nr9+fl3FMZ6QNkbZ83S0TDEOjlzA9NVz9T6Z
eO31T3o6/o5AbMNASRLNp9s6DpbrmxSvWvzoPM5gABoZ7LfxyfMh5H3/jBfpHTugvHeHSf+EqwLQ
4wFDNTtrdFA09S0n+VMuAw0MSugyVWGB3lNhhBHqG5BlFpoSGPZKHunohGMoZogbpeH6Q12EMRtF
NrzRNLdjvvPz49/DaPONU0kkkxPRd/qZRtI1808LcOBe41RdW985PJR3DqoC/Ongb8iOHHfA9hcL
c6vZuzSJex0AleoSIWp1146oG53uDmMr1ACxqQhlhdj8OSenI0JqBqH9ZXC/+VnscDG+w1Vf769H
x1CWefHfQcb3J5+04x9l16AYjemDmDmIdkW6HMEeFGm9wfK4ojQi88wi0+KfcgOPl/0KYhbQ8jL0
6xZoySXXW16NxFSP2U7Ij0ditlpqtqOH4HDrrakOrDu9IeVl5ixC3FnrEzETz4y/H8RbFIhNfp4l
R03a1kudwqau/AxnYy2m9N2ooJeSCkTPk9v/8fbCS4aFN0am3ySjxKkbQqrlP5DvjMeOaMzniGm7
wfTRO2Pvx9C/PznSzFcgDTF3EymLChgsnSY2eYB1/VaHey+xzpEFL5ToxfZtJFgrJ9PLoEMEKbLQ
2s+OzP3js3TUPTFiejH5n80EUaKYtYmvfrq9K2/5DXuhPW34xHEPWpPNhzbLTn/wCR8AgCDfqgE0
SRL17fdJjR4FDq/a+1h7MVkXWCSlLSN34GFbRsxJfBaatfRY5f7PByldz50X8BA2cS/tBroK0lZx
45m30HSBYgEq7vjBZHrc+6LzYkQRWz3dqUGA+Y5GiSzmQOxWpgPB57JvNybJle9DPn8tRNclAK03
GlrEvmqgBjD6opeNEZZbIbnxkd+jXjhHBib084q2AJ7pHt1Pvgd/zOqtJ2sUI5LTpjzBiX6ERGxQ
zwIOdZF4DnTzl8+Rn11at0KeS6+3bTQQYp9AFqgEx3ocQ9oA8jgnBeLRhPWHEu4yOp1m2sH6ZBPP
Q0ltKIE9Hw9ihCh8SdDrU3m5SKSa0ETa1flmSH+rV7wEh7Wf0sYfeFAAll4T54DkYrETH9m9JDa2
DLCB/Ud+SaS2ZyMvQiZrvqtbEtZxQQvQn7nR+7LFyOHH2ZJtDDVk1ILlx+fKgEPQoNA4LVo2KxKA
3m06rLAx0msFXJ3VxIYQbwnAjd8Re1efWLhZVu0lzT8QSzrGzBwKBkx4aGkuRj8zvy+hrgCT+EVw
cF7dXNOkX3hBn7DB9ofNrYs+UMOHNaId4/1yAruq1F4LAfOsf+YKrEsRCpCleiflqqU1U1WpCqjW
f+7tGotYMA9yWrQL68T6K3ojRujgunGwF1C983P3S2a6tNK1c8AEb2AupFLtDtr7t+EDEiRiiLkM
QLrGlrfBOpSkyh5G5PVVludAjShpyw2c/OKv+wLA59DnaauYX6V4AtN0QojIDgAuXim79FY6E2kp
6VqTPslQJhpuBXYA6IcOxJkPyDaCBxNpOAY2DoA0xRIhbWzFZl7Hmn/sZyUy1/1EUJ4YpIZIegeE
9yryUp8fs3EoEVEL9d8uEDqcNvO4cuf6Mzc3GVZmqQ7UhVDClqjmXUlpNZkrRJbALpYnL6riv321
B48GUb44JWHz+//VV5grFfi3IYeHoceTZaV8v7ozkID+Zk0lfBEJReVXMZCmWWvW2Dse6FlF0KQa
KAotKao91fBGBeNzLKwdFxEgWj6jJszr3hgZv/mqF20qqgDKmF8JXiHupviDBPVSqS5hde0rkZ/l
jLs4wlvp1QddiEa/MpVwDUzQ8K7Er4wRN2710uTqlOX1vlmSE+htGZQqlMbMqAi5+8unDm56eraz
ntZxelb9QlZMk0EA/FEUETyRt3gBy/KMpVBE/9nthEtD4L9BR1B8J4NeuAEqb/zHeK80Wh4PA/w/
5A4MBKgDwnfnea2xvjQ7RTRCmGCHVRA7lSiC7HD1bpKMAcvWl/NXaqMiEPAwexqAZcF4h7uTdEq4
BYJnrOWDXSKXMLGjR4PauqOvvnPQ7M/biA0yZGaQ6h3wRtvRCcuFDLI2yp15qA2wduTGbUpUAmlQ
5IwldeaQzKW6K6f9bFallqDOvYyRUG3UUEOeS0Divs8FpB5+cFvl/l6oCMgoH6NO3c+QiU9Zufed
VBZi4XBKDv12upa+00V6bSJCQf6EB5ztdlpFkTI0Xo9U893H49DKtkBEkjsHbXbRsdu4bMKyWcq2
0cu8P4NQhZvgsIzjCdIiICLahUowCKxw6S1wPAL2XXd6Z+QOT0ufDy1HSP5oDkbSlVLYUFsxoXUT
BdlgvpUgHTtjc4ohFacfe3nHN4VAwz6GZXRjidqyyWJ+/ibAC5uxUcvIS4fuxGcwYI8eXNh+U9SI
xzpNf+ODIj6KproA2p0dX+c73DSvAfT/SovaY8pNLtEr3NOC1cBNorb6+fbyBCph3y0T3n9+/gU4
kgPlVGvRh+UvTw5A22muuo/PYuoYAm9F+RkuyGucVQVsC1NKelHlJchMxv5aWQ0SORteu9esdbXr
tW/AQ73EhUMzXbDq6j0ict+VmdiMb0TYe8z47gxC+8P2Mj4tS6C7IQdGdipsVvTC745cCxWw4WGQ
PbfKN7M87KOy+W14MQLZKxcyS87/kfq/9CwKabBw7JeRWEeNXwbL0vdoNOQm7tQhFOV7oJdhv4Ny
VBNL0OhomJLvxQZxwmQHK8+tlBdlU7sUkHxFitVsQzHOFLcU+S8Mi6z+9hn5SuEUgFluoy+7EhJ9
tEwl3z6zylhEEIZoLxZhvDk4oxCPD5XEsFNL3z4gByk3p3O7+EsUKPB17zF3nj+h27q6QehKn8Y+
fRHtS1HsZkAoIiPZtQbhWdSiiRkfcMQUFHMF5u1qpLRArijaEF/yFqWRBsHEXIXTvMZ8pu8wLeOM
U6NLaL9Y79r2vnpHgVHSIs2xd/IUnbaVArtOiizoMkdVpJ16Bt3aMoMZjq/sYZZH3d9UFrl5P9CZ
zFkeaMPfABsdJ+DglXM4QzvuB9as43o5EDs63hJNROUqr6SlQ7KzFcZIUdFk6e0ZhPnL0AsTvo8P
fjQxM1UsQn6ojtygztQ6caBN8BRH8GQmK/31FkqHNdWQkDHGryWCoIcDRR+Eghcm+ekEADcasDrE
tvn5rGFSqgVeVjXNKHsnnfQmnqezEK6HBExW4UKH7Ii4uClGjUCDItS5Kjb3jN92yLYAo/Dqgfw+
63jEWdurdkW4P070MTl2Xx9uLj6EbqnFBZInxOjzoqKW5OskC8b+/pWgPv+Aq0KMwTUFdyZhEHru
HMz9MpyVP5sJGkq3zdbretmj+4qPs6WUuOdAWvJfr1IWi61zXzb+8s9/7naX5Z2xqrYMBMj+BDvC
mdeu0JShimrFuJU3SqXAv204kFtQ+m/Lyh9VicL6OMCjJzXqAXNVCC9zyZHCUKBIxgDnun78Icdh
Y07Nq7AOCUr3zE+j/IKEgPZrqdqgOC+Y75yM6ntfqBgsBnRBFYDaBc24LhwFQokiOwVK2zyhfe4z
8H+GdTiY4g3VTwH9QFmMzsC3NOs82gqPY0oJ9H15gYCM0epQi57SQ8RDIKhmGqhjuG+l0J0Yjok1
EoqoceViSDBlVX/AyFx/Q8lx0TnTfm2YwqFI4vXiQFdMFODr5hmH5zitF7ZqVPOl/B42+uNfnFNT
bb/W+MtOA2KaymXgx3BB+D2/R2AfH8yyNsIcbd76dd9hXq/ZsQBoPDWmSoZgypsyCYJUb4FPQNvZ
ZNUO97hlQieNAU0Qm/PHvRRdHVfrleuiLF8deBP9AbtJb+cDf2qwRtajHg9I0cmoBkkd4r4oR0eL
IHJsPkwuar5T4dOQEvLYAdnf+JUF6j4BhNrlcaFqShVK48E3uEWsoj6Vkj/dFIFHTyiz6Xofhz4S
/n3DQmSGlMxK9CJNEmp1PBNoRy1pR1rfsfDz1p5rKC7e1Fwe+DBzqDLvcWqIRlIaPLIwABWVep5h
8Q5v2LEBfXrlPPfvs+NenMfe6NcTZzNxXtWtJgzvHVga1OrwUDS+I5tW5hbsy+lM8gIGkzCJTF9G
a8yDyzx3Kg9AEYeK/ynAclqehr12I+g4zJM8g+YFLX/AD7KktTT3keYyxO89BFKotKX40Lh8cPDo
GfBvYR1l6KDNckj2XS2nUtUbP6asEUmDMfkEmrzexcclMMhtRe5I5HGsjFH/Q36BojBxqedhkOEv
r57+eO+oQMbqiExnFSjwdX1sBvxavzWwsHNeMMxePw0WJ1jNzSLLcWWmNdBRXCouGL7CM7XWziOo
PpKDH6K5QPC/NsvBngNMwqZtv1EnBiYPX3k8s8Vx8hiVqtE5PIVGFkrfjFx6DszqsW8vFe8o+Xt3
LCjdmqtesWDwhIpKu4BSY9bakn8OfRhlu3DCRSa05FmaOWNJa5ODbyb5v34C2Dj8QkwJ1HDHOezX
kC6qB4+9mSn1Ot0sTq+QgbjJYoDHaIEe862ZFuagTVEFfOnICMZdYFMtJErOzw90h7cVzR05r0V1
frfmqEzattf0WiSpGRsc9ywcATUKJw0SAtZlLpQO6sxKUStsVz/tFeqeRI/Oa6srFKOk413D2Alr
OthGgO+fpa1jlhSThqObsQZINuc3bYCeHCvf4OLYD6g4/ZVBNAhv8uwOC6hTNovDKwOi5M+YRQZW
e1OGNQhF4MJnLk7tAzIairRpoIbhR5RUp1lM+7ZFM99+1e0Tq5TO8YXlW3nJ13X95sLYEyplMeqa
/lDW0hyQATiq+H/PVNSSbvm1CavZaigbsYNJoocGpowfNYlOKg5RD3GiBcCFh5SX9t1KXUAOsxDj
Ow0gwMed3f7/sBob5DM8t1EUL27kKbhJZANWgV+zbcl/YNcpzTQO3tIGSnHnkS1cuuzGyVN5LbSv
MnNLDyKjAOU9y4WS1ZRv0OfStgmnDW1Z8k/6T07Ry1M8oAtq6tiTemmOTXqV4EfRpS0K774qNoB9
IpYlk+4vqfwd5fWCxU5QUmuVjbQlsfaooZbEno79MjsRbg84fDjRSrbIEsl9ITmDY3bfQGKotdN+
OAaXZenLCQSw9q5dPeDLjCeOALJWj87H5lvQ6zLrxVXk0W+aCUgS7pINNXfKw+mkBqZZEZqAujAH
44qPQNZUgepNyBRQd1hgp4IPW8INPDAvK7+Sy6a8bY4Hj0tW6y2qbCc4J5S+mAPqOfvgPpVeK9Av
xYdvdnyzX/EB5sXq/6H2JyTO4dvZ+8RF3FnsQ2YZJRgI38YW10UpIGrrwXX93sFZ7Mdj33h2pbac
D9qB6x7t97l9daI/hzFgeu9U1hVMxMjO4RX5/7cAGODJou5Nc0rHTjpTG0QMC3xVrJ2g+WefvJJo
xh8tCLI7u9Y6lIvif/lA90g3dg6BgjAhz0uQ0bLHfewXIcbdmz8Z4SqscLtLYt1/NxC+KZwJ2fyw
uNtCesVfu8PbaFyjOKE0iWVphFDGSq27M5vc5GyVSn4ERseyXL5DDoPlQMQ+g/8yyEBIIIgvtAcF
SM+E/WpZmHs2obH6rzmH6KjkfJSzh6rlp6dx7G88baSW8eGBdKL871AxeumOpSegYTJEUive7J0x
Kc0Ky2R1qIIcykQ4KUDZiyT0Xx3GMo+WvtOnsXZ5Q1fVtjwSs9mFn1jx3/Dq75w5kO+2fZSEShNS
xKLYaQkXQSjcQqkDL5Mg7b9/KuDmmrApfz3pdJmCCypJnev1Z5kaViMDMxcZgjPue1eDbCR234ud
96XRxSrT/nqWvb5SeIIz8Ybqz776pM8rws4Z5gEGIlrkfikvz8whgD0VDj25yz6fxtaidWr3jBC2
RisYNw3jtwn5co77WTu8M/5b8O6SX4w0E8yFHbGTSNi/W9BjTHPb72r8u2ofWT5rDG8DhvmCn2Zh
G95n74OkdmB9urDu4Pu6WJikirBF0Pw6B10dT+TfBtW+eWvorK/pdijlZgaf/9rmwpNR9aI/32bx
IVpLL8Dc5LbFuvtTsHEP2IJWjjRul8IneowGHP9hTAbduKnCL7+PcqefQOaZP2o3QZu8PsPs6eQh
21V2yGxPdEqI7DiF2RkB8iV4rse4sXcfv+fzdqLBb1h4Z9c41KRd3hWELI2y1Zh5v6vp2Ph5qKyu
U3bcjK/F4tR0btBiy6ELp6aOIexhf9wKSEqPhBjEfRih7UudOqjJfQjUX2A8+tFUY8E/cDZbegJX
VDrL1JTDdmZe7j/wzs4gXShXI7sm+XDURkOoP3Ivw2xlEALWV4vIiWCRbuNKK7UwRQEgtFKEYFQG
2QVP8BRVb18SfgQOy+tpMcUT0KHOxBl/i8fGKlRflvGDbYB7xR0SuxRlLtvZ28QJ+HqxllTEkC09
2UpasIevkshGLOvqmBj++JfMl3kvG9tUVUaovGco1CJ+Vg6PJSWm1GWhThCNGWnlY6+Ahpoj/bLo
UXMkIBUJXTCvm9bwuBeKOXj7wKe8LeLBA61La81sFy5t/s0JyPg2sCAIwWlZ4VUPP1i6C1yqHebX
UHcWhwxZTSJtXA2N3eoEaGl30hwCdS40XgpAWE92mn7DvgZ4wTTB5yncBP7DXw4dG57ykzT2wGbA
8O/3Zjw+Cva0OJw+X1/To8A9yBDwFZT8E1gTcN0869lVmB/ZKHe4T8HUTgYrSG62JGNODoxg6MMt
8APMyG3Lvfj6H5L3g3X3YPpsEQwrsbU1HFHAbEZmiX3Lmuu4zrnhmy/IPIyErae3XB9WGGO654Nc
ZeaxA2XSMy0I9L3qqoJwIjpjxr9yUmgxdw8Q9oDpxLTIZCYUuHnkFOkne3eczRp9bPLpx3j+n27P
VyuADkntSnKM55PxCU9JI8FXkOJY/73A28/azjCbnRVp9ro+EDJqYr9ofK/Y8N9ljPFOQ5VrsOAZ
OHtDy5iy4UFdGSW0PQOyFm62r/bNAXe76AMrFj2W27BNw+h8uDWOz03ggslaIUwNGDFpopRxyuCp
lWbe2TaZgG7ijuA/QVb+/E2JH/UhiuJSCKTmnejSYU0uUS6kFuk8zo5a3qUmEA0wB96jvEYDSNXx
GCaR2TD45+JQMqKPDXyDH6ECDi1kmndlNq4o+wJmnbDAFlzl6ZnxDentWu82OoITunT4Y7Xm6by2
S0dXKJ2BC1K069pXHPgRc7wBDVmKnNwwx6Zu6H+ReOcUaR8lvq/AUoEVhyaCr8Bn651BWNsxq70K
AOofMkZyI6zIEcy2YIfDtM7BezTXprMEtQRFlOL29Ig6lfaNf0zTQ6vBBvpv4lM88Bxu45CjJo9i
bbc1vQ6VMRc0WV1hlbg3g6+3LTnIhA6CjCFCWtEas5AGRFZp2Nr0Xu0jI9X5c+rSysJQDzxJfEor
SahezUKj/X9X1YbMxRgaD57okacfrBTADmf2eiLr+AslvcwFMI7uMfiYmSPa09F1lUgz5N8K15iP
QtECaIUNbluPAE9tLKaCPciTNqaasg8t8XD1nfGD1IkQV5mwfy0o8GNlhl4gxRriAyZ/r0qqm7ej
RXnATSCUjF0IFrTuMyVMKbIsfcbOEw+Z/h+P6yIp+HvlfQWamTGHxDIfdffmHd2cCjQIclrzyRC2
FV86wyCBtepI3I1LjtHHpdmS0pYLOpWn1/Rs3tuX1u8T8PUBfEFMaY3m4oCltQnxAjoJGFbUCDEZ
CKAEdu3JsYH5HVHzZ/2MsBXhnkVjKi+klYbsRemJH+ciksQNZDFy1+QzdVB72W4i5+nhg68f9S1F
lhuVCtNiCmDJC2cZAlxwaRaPx4bVqsG2zkqXPzvntdbb4aZjPNOerAUQd60zWg7kFFVBMLjh7eXv
Wfh62kMiMxDP/RFiSSCe8iWXugj1ixjA/DeKwBd5TMkXsmxe2OjlPtUVUWiiHxGP7/g3KVPDTiFx
G1VRbfSa9tf5euEBSioc3HEvmVH/7FYOE8cgL87wzkZwOmlxMpbgzzw0r7Qn7BmKMqKc41vdTLVt
CmKRANDckaYTjyaRaOwfeQExhg6OQYYHeyKo7xuv5p1kWIf7YLqCn4IvY6RB7P7gSlqLqPJBubEY
QCQxbAJWn6Y0cL1Zlc54wig4PLle1Gn2rcb8mEB8pw7kSBrXoV12UB1rkhBJUrhBBb90Umdad85X
uCnqf0wCH1bpv7HjdTWgP3lBj2j1uDXcZjkHAqGrfYKYGAnI85VZ4ymOjFNVR7JzKhiiADMvOwpl
6tr01Z5a2xRjG9jZI4nkXCYkfNrtIF5RnA4aW+BgIeCujCX2LMy4HcpWFgYE6tk2byVFmoYGCzJN
uumxrubEOPXJ0UvhiqkQX7NNmhoJ9PSwtYJi/by5uGGijKusHame5/1AmFStaHNTNWsPxshCQJcz
drapC4bNo+xSdVsmSWf83wdunR9AuCNs6n/bFr91VQp0bsnGEfVe1ITpCLTd3Koi9GAr6EE2Q/JY
FtxbQV7yxWGV1u4X6RRu8PKeY0q64v/VhjCj8VYAlXroq8QVCD7q0YETpso0oKf2W/hfEEEYS/eD
u+8pnL/paPMv4sFpXH2EHnELelY2j4wXnb8p7pbxclLMOKGB1aZZDr9qsjlZPhQgucY/vXCY6fur
kAz86lgRBXEm2f5XLuzRm66XjU5WQzja8LTUyULCy0pvgawfyPIn6aXXg7FSVpKvwUC1PPslj9Hg
knsshxhMFipv/66WSTeMy8wo1eMr/OIyiI56s2YzXZNl6CgFgw/RHmdl/G53clHxWa7pInW1209p
Yw7Nh9PNVSkVfWm1HvuDGGdT3+E8tDa/tH2Neoqz62q5GaBCgpGFYyTrpauAyYtBfRsOFvMtIgQU
r9ChX6+4i3wAZ+I88epRQzTHfFioMfoNbU4yHQGFhMyGnpZ5PHrB99NNShbKa+SxP+HXgMRxWOAu
axdUm3l0gW7Dxfzmrl/8c+kOZKvuzAzi35Zdv85nhMIqb7uwviRn97NKS7eerOiP8OES4+HCkum/
eo8hLMiZOk8NuRoqdDGSApqVVXm7ksvopTd79pWD5mCf3oC1zAPzHJxNAb3nYg2bWJwu/66jajQS
Q+fzmjPOUA9c/jgA6vlK6eOubdp+oO/lhTj6G5OEDIAqADdq9ylK4ls1ucKSStavPct0C2e4zwfL
x2uU71edGsXRrm1rppToFzLb12BoYXYftLxWJCOW6w+fjbu+3F9gfFCGXK2D+Qr0xXqxlIlG59oS
Ou8n1tnHfzHBED4wRrpt/rrxGn2iasvCRmW5Q6ePvC+oLHp0DTXNMsNpYIHhk860iyj62y4YOyod
WdWBc5MGlZ/EN2O3Ec/LB4gEQfapCx9K+IgRtHrHmIqZ/zUBQ5CGPEszsHe0qoGaGG8Yom/lPvOg
nZf5MRNQ/VD1Pf5vQyWBGVI5d/Wl1xtN1GxUrJlQbdgdSbXp8UH1rxEzzw0cv89N75Uena8HghbR
AYKdDc/XZ1n9wY10jcOfKrCaIjd74+vnWTq4JugQgd0dkRKc0EFcCI2fUFoL67FZoCgaBqn/n4DI
Nv5wiXFsuA2iqaSx0nHLw8nJEoKyawnmrWT4/4vHHYABd80yfWV7rbahqCA40LcpPYzPQ6pomg30
HDcmhetWEo7R5jA5Q9zr8zWfTPfVpE7o0c7UvTpLUnngIZF84QhKCtvvE7Ogja6N5+fbPAiKuGB2
Ygfab7dwV8vUd1QghHxcvyPKPNupMxQkQP2MiY9CGiEiQbsHpoC8ebWSEOgoQNV+spzIcq0cOetD
dzK5KreCdx9a94F9TH+cTf8Gg2fGkKjr1lDQe1ewR/VOhLXdDnh2n2yNjImoFh1yfx0WErvBuwdC
FsaG/kFZR4Z9vqD7uqkY1qkw7/2dxziuD9paw5mpymTb9ktTYXLgRPhjNWyJFz5owA2tNtTnoPiJ
ZLAcpTtaPxonErJABhU0d7PZb8AH/JR4FLeH3OVt8i96QNV4CW9pU63+f5KOpbnIZ1Ss7l61J2RW
vYdn2Mia3vAThojCr1tX1SZoQWSCGoHWc37xqsJFtlMm0QkFuDESNyPuL75kMrPTJqgF38h8tUCB
L6XAZCbZAPT6dgX6txy91UFY1+/fzcVJXe5g82sgjMdD/xx9b1z/9FMkNLSanF3GpDQbQtEZFOHm
lFCSTLUF5NvARTKcgauu1d88YAOFAmm9kA9YymcqnV4Fi+tv/12UrEgYYrXqJoAzHhRpWPEAOUeo
4m7IKVY9N8B4L1ymxBSwTxSrzTwqUtvyJcev5/3HKp+CwzqWH+p9W5iUWJcFCAxgfcVvhC5vrUnd
bIAhQUzckSGboZV82dY99dEpgh5gtQN+vGX+dBf0MDDm76pzD50tsCXUUJUDQhS356U+nlSnwDfi
j/DHzeZU20/TLwbe/2dyr/94GTGCXFeRXlL86XE7FQX9wVu47q3n9urrp49PaJOyYpOqOiasXDSE
lH7y21XajDNZOqGqajIEsBK16qzAL0B3Bfup3FPiIZs0oWncaJvDZuZnrsLn+uKFMeclBYhYmlTI
TgODniA6NoCYlvvnqrl1G/wliHDabUVgaFpTyQQ9PAIZzm23OYIQp35j9M9CI8vzIofmeKtZc2s9
C7zgK5aia3XctWkN8DG+qxaYwHZ9Nuf7/dCg8kabDlC0gy6U4Ze6dwc4NaI1ngUkSqGWmt4ck0WA
3gHe3MiD+0x5mCpyndeQcWpISIIoNqxvRDY6u8vWZPB1tqEC7wsSLDRj3/Qwb7LwEpYQgb0YO92Q
AfVzW6l9ZYn1mDkRSDK9n04aZX7Tx0kxPiW3z759D4T8VI8Byx09Y3PyjAo91Yx11Cnq6hK0ir8d
Y97mXfzDeZaX/2XOsM0+lpCG3gAeILgii8s8Le+6aiTYS4EBSMXF5ZCUJdwoCDhVhTEFMBbdnega
tA2sFMf4idtneCTM4bHTJXjwcXJ/Rt/rbdif1PFxYk5v+mixRoDr1/a45vOAnbFkv/6C75cX0kJS
6kUakVODo3OzMMMQz9IUmH7EAevZD28mqTQIcRXO5QCMMYfsNAyLFPrHm0mpOGjz0toRkE6F5ex8
/U45/EYOcF3p+aQto79jvd/2dOf6Bjmqn+C0BthhEJda9wn8gar7x5SaZeDe8MRgSiKfXYpnGWvd
wWvfIYpG156jVDKUTnZseWEJ2z3yftTL8ruJs4SO7QSxuyXe8Cts/ZZqnH9aRf0TLrZMudvYpU9A
pp2V1tuzQMkOog+nN3fz3/mvYWKyOpjUMlbOLQIcHJgK4LUIhsft0QXH6MxP14Mu5oc3h1XUrAAB
OL/rZncXjgqo5nlBgAjktRQLiWw50au5lOVt/VJjPuhqMzItCSyqfGq/e8B8fR/d10z2ZqNKTb9y
/4ShN2J7dYJ361yvfkDY4H5+AxybDSXdhTmbW3TVBXkPeCOjIgYZsECTTlZ6jjwCSRMmSqJP5kIC
eHYSKyTNNW3w9TIh+Z0hKmAckg8KVDH6nfw1GiIwltaJL9w5G/npZapzHKtUDwbSWLcT8UWTuvbe
xvIg/RQMj4K1uiofT7XZ1wY//XR5/QGtiNGusWe3+v3rZBkch3TDHyVvPR9k4EyKBf01f14MHixU
XjbF6Y7YOiKDzShwLo6Yvgdmh8MnUL/MdtjzQ64spjnG541YIouu3WuaHBlrCxmtY0NUG4o9vJUR
s6VreM/oQbNWjgGd/rMJUVzxssjDpRJDWs7EsA2BrVOzlH5E1Z2+AZDm6d8ZDiQSPDiBHLm7ZDrr
+WrjpGB0ltOwGOGwvgbeDVBor4COUbQwRNQ/cCTh9g3HqXpHd565XVkeC2e8eS3c2+m93Z2yZuQl
cTZN6lrCR8hifXTupqCeDyBHmGIuOv1eGy2b+s0fPe3wIfDruZvKyWTVa6Q6zjywsW4vZew4VjTZ
Pnf+s2t9rlgo7uIyGWwp2TgykE7VwkMXrGqmwkvhpz7M82w5MaxLexVxfJqOxUvaAGsdQ+2h8Tko
zjoKfpAoqqVmGEnjxL02v+8QCdN8pCQFqoDO1b7nqivc59QSWMNvFYUJTl+/gnrdvqCfyck9s1eo
WS3Zxoyx3NFFpjZzdoK/QE+QG08aKbjerOC9P4LZG4ZE3EPxEt4F21ue9/L3npuJw5T43bplQ5AP
MMeHDesOkFc7+lFh1tFpGTdZ58CE3+R7mfT/k5zRdbg31hrBrqxpvhDVOjXoy8Jk0dqjQHuZaUzS
VjWPIlfUBzTmrgtraQHkYO7a/anse/nxIAf8nrfjxPoNaJ+U2T+u77SW30f7nEJ/Nzj/uf6JJq2l
k7fdj5qRxEIsiOOVZgXqrXg57i/2O8zA8wgWRg3QHiqRtjxfAHnIfFe/j9zK3PUnrpmVuLoiI2j5
r1CzodDD00H3ZiElLSSSuyfxTkeEC9xnykktM+2t2BxLYd4GcgKT1Wv7zUdbfSwiF4U2Txb3Ao4f
szD2ydUC4dhT4rOf2y7xstR6f+mIzVo0SUE3IOHMsEcBUjwBI61Vor15Lybw1keodlpGyH+k6O/w
BFpCD5qnhhpSlTmPeK0LEE5fsyDoqL5oQg+nDjiyhFrgFAmPs9S+3LyZ5RNL4XiD7f7CC5UWMk2S
4ucVxHso7q+QvzctPvfkwqAZYLpachRwZZU4yudDVXJAXXptdIxH9JTTPRiOfNecHS89u5dM26ou
OPToLRnaeD9PIuyXBoPrI+XWlEZTQe4MLHfKcmHVdBMpW4G/uS5sOIplmYy/u+hADFF2AX2XHMdu
8kOFt/93GSaMynRWf6FwV2t/K8Uvzb6G7xlOIuNkGXZbX3LBw07PPjR3Hete2Dr+Y6w19thr1T+q
8EtFuA7knzWpyO4d6FqDM9LWn3zzAiYxnPV843YFwFfnWyhV2AqBGxsC1U4xmsxBPTZ4kckVYv9A
DoajxYI98Mk5e2OIV7Y5v9Hn9IfLS99bhWNFLjbxMpVHLAfiNDbY0ztFk3wM8FzshPBc6kzOYNUm
A2XTrQaWAfCCW+7q/ghzDCcYkzBZTy8qGXaOvmNsDI89z1LystOGhUGhntMmhhke8Vn/U6V8JBE5
k4RYuklvvqnKH9D8RtzdcGLGrafa3b6kgf7laSOYHX4OfgoNilGhMogldz7ZH2dEmMO72lgOCjtC
b10J62thh8N+4WU2cui/62YE6nKOLKqqtNPWKETvdERsfIn/5zCq7SKGLX0xOTElp6kO01qGqLsS
BJq3z2MSNmnFV5OWpGUoOaGr57w/NAWOD1rg+KLGoArtI9KHnmuFH6OpdPBsuRPzpvQvK/OOEoiy
CJMRjlz7H+LqfrUGiT8GmG0HlAm4or2LeQ6W1U69LzsDbJ3GqUH26gliOWNkX2Y1CJAZ7vHlpe2/
pJ0J6zWvT5zVPFywwIlerb5oKpJfNwhfGlHrJKKESpxIFKWBwvvTIoVRbcj6qJiRqUojl460yAzb
lphnlFZPbOdoAryO6kYZHBNAO1gZ+S4STLJ81GTGwpVCdMDThF7UfJEsObY5Jq1tsvfNgF0V48PT
jyRNTHmNgHJELrAqIlm2+bimfYsLGw115Lv/dHk2MIEC2ni1aIXO5KorkU7bN3FElqGHhyeHlVcW
4udwNv0IRvxPTGWFiWKnm8gna4XiflmdgmLQ4ON6gm+J4pSBdiHJGtmKpEswRIyslJMkk+lVXbjM
jaHlPIkbtPBxJFNCaDSQQkwV1mbOZqgrHcmdBZKj/QYvtKc4c9nBzs+7+Uw4fyN5gQy1cmdFhi0t
avCY3Nuoi1Wz4CqrQUzjUqhYcRFHqRjD35v6MqpH0C/gmwjETUykrgPL/22nqE0fWIosJy4+ucSG
UG4yMhycVgEyYIulXEDiec6vZ15GCwvY+L4qrCaXkJAvWldM/t+2WAnZp5vke3gtHpQjvotGOMtf
+Ii8H64jVM1W+6f6k2obyDJRa806YrNrr5Kng0uhhSTYL06+2lZOSxi2OxFSbhNBQjf467wf9uiR
qIvt/wXqV/bkiL0NC/LWKIO3T1Nwtm9ridIeERtAuKBiQStUQ1m7iJsJ6DlY4n8VQGbIwJ6f5XcP
zM2t+/ge6/DlQ6fwV4WG/sDuCN0XFYSYlbWICJyfV9qtCk0VAh7Ae3KbaCXjLbq462GiTtoNOOll
m2esq1I8mPP1MpcE14UZRIdQkHvi03x0gSDFtUc5LuXrvPrpflrwhbDhryQY15Wxw4Z2c1HWfN1/
gH6TUg99US/b6AgQ68rmuJbdTumYThwuY9B4ONY3dVa/PlmhmGnkIOs4BO2W8LJ3m3p+QV0ilAMH
xrnYdkfSf02MipDo/AX3ShuShgn+9j2QdKfpNgAOoHy1gAkTolrVHY0MGsAfxryOfZHZz7+trz+3
PdlU+ZUwNfBDFcGOk0NAedlm2xamGj4t8QsdhfQEcSd84pcCbRdJFG+yMUJv5aUaByNxQ5MGHR+7
kaN2Kg50ra8FKml9vkS0LWAJEJNbmXx+l5d0R5R3wRw++/sYraCd3mq5zWJ7/n4MhYPC8xCGe6SY
KwZxTyigGUB/AYhBL7m7jnXd6xm6i4m3702B0DgVcRf46b3cY3UXjy0RGNd72nMzhYNRMllDeBtk
0ZnV4aE42Tt0qmrNUi08UpuXENM1PQGN7jKv8m59j4u8Ywyay+DRvPB8V/JqKk4y7RMdNuFTyg5F
QyoF0+YiUtFL/KSKjf2vSuXLb7/P2My6cZspeOKWHZaMFWoFA3r6C9FHaf8Q3wIor/n7FABndyVy
AtOoJ5RS4DUZCtCIBeQMZ/yF9dHT5XHPhZQa592qiv6sQ+QparybGQAHocCCzzUoHHl20cJc0Cl/
rHlDN3Hcz6kg/ddLaVjTqavLAx61Dq+MrI+C23NoI4WwmY+rZYeZpHlY9IZWdY5VNr4RA9smo9y5
k7hiuf1Vvq1d99mpRqEX3qXquq9NwZ+ikT7Ex/YKOO1PwVQ2l8Zwsl2Ds8j+IfoI2WoDE/E5o2ww
6/UtjLnagm5mTu2cE7PVVPalpR3rVoZtuZqSk/ZJXSzkRNW1fYKXQC1iO6AgFUGoY9V1+a/kI/AX
TXQDTXYEMOiWAuV0Xh/SRD18G1NBPDizYPZwE9OQpaO28KfNnD4y41odbBjJJuJOrI8n0IpovKBn
3lU1Smy3bP05N1RSeno9jgBApUl/f1WdJ7JXsaIolWXhaSrHZyJXZQBZlp1hVY8c00Blo2BfbkVk
KBc122ewjxWX17sxXcndBTkky/kQ6ycwey3fIwBDUBV+qRcVlE4z71/jC0j/VpGuvBbf0/Gc3pJD
AlNwACklrYjTgv1pJpd2gTONlNq7X5PAK4CaMoa2B+jrhKecAA+KSaB4oYugZIlhdotdrRSAgxwN
nPfwsMpsoYBSkigM9DuuX1LUjkCKV7BoIlW/dmV0FHwRDyA6gQ2HYi1Xf+Lq9yaEieG2v7kOMx96
itb/hc23AQKWogpQJ/sCSslnEkcuRq2CTyzouBBWd09YPkcBCqgHpyX82LlIgTcB6RaA4ULu91mS
LBOuPALjO2krS/9QN3SLF2mFRrGY/EcAww5Ko1wotD0u0RvsIFnfCFZ82oS+IesI0KjdHhjoiSC/
kpdqx7OWwvQkOzn7uW27xdJ3OsGmkIJTFVR+8Mxus3csDiDR7Enx5CT+Ddam0P9FJB9ndAvI7CkD
s69EYGe2TlGQ0AdoUyHHt9mSQ9rhrHJrkFs0wbFwj75FEauX2zsd0++6Qhy5UKd/cXFYwNM7AC0e
R/Hq8VebI4HnYGqUrn2rOi7CGea+qzaw0Tpy9p+MDktU/BXFYqukl+LoXIUUT9sEkWkEkrAMbb1u
r9Q9s0HC1L6g3QTSRtbo3IIxpIr2nhOOTijcZd5sffqVWQVPkRCmvPCWXBxCAM37dW1INiQNle0c
LX6sCc/GFb2R5LXKZFP+fE06tNHxsgnOOTFRCLGtWRDkd0K7abs7h4xprmwO8ECnmCaXA4UWxhI/
IIucPhpbd3T94AnRGFBlNK+A//MNOwUE1x6O3gae+wCcgyAfN0T2AuniEiKb44441k6a8ZEAUjQa
lp2pBozjTc2StSD3yAbYUKAIt2aLvPbCQj/8OFiGNv9J/5ghUKESmrBvKp66lmQ8iQuojUc3IIBO
9zOe/4KcK2PwDRMHCRlkVKd4btISwnxR2S8p7R3dlT4kots5yQauXXrd+KlSz5x8R74+zLG8ZTqC
ctjyCebtpdKmnyKS/oaSwISEow69TuippjIR1Gs8dk0Pyd6QbVo5iKFvLbjs/deuaVKF02jygxn6
YZUum81VygUP81X2qLgyo0DTTPWgSzERsBW31O02j0m/jF+nb+e/R8kpkPpa4fSVJFnippUUmFAz
C6b3+ea+p+SuvuiaNi1xI//SGH8gphMWr3vqbJRliSjtj5edmbXrwKMqEKlkNWUY94+XlJoUWxBO
YVnD+Bz4jpCCa9ylcyOdIwabSok8qHnxv8Cc8Gt2KRB04OM1mqhKqemWXdCgJ4oTMfAWuGCap/Be
Q5Vb6z5upsxwdBCYAmFI2UeW4jGfGzx7CdoRQye5+M5hQUbiyYhW1wrxz6MuUN2T1r/3MTvN62JL
B+CvrKp11XQIuZBawyQk4do/g+HbEwgI3v8lMCQiYMh1BCD05QlbqNwBZH5xoQa9UQGTNT9D8PHs
c07GJV/heMl2L2tRgL8PlSFWxHH4AZgdIUt915bqCYC8r98Q0BpsnyqWD4jk5zSI+9PmgMfs2TLB
CHq33wvSel1AvZ0Zs5mV0QmSNLLH5ggl79Z4NFvKOqBr9b6Hk8S/oub7Jfqk5JMOlhO7Qz+LSTUZ
2FmfjRvRfkaEDyY+KNTWt5gtdJ+xSpnuUsYMMY0iFa3MAbbrm5rA9D997pyR6amJL5sdWG3iAuQI
FdC3uk/Z6L+IGilm/4JIxmqh1VqyFTvi1T+xJoS6bHHIRBQQXrOs/IolQY+qlFtkhFMTs/KXAbND
5wzHXoPbhcm7XcqOfcVZ6Z3xZ0Nx+3h/0hQCw5Ayuqs8J7jt5cr/HXNONVF5qv8yzlbFlF3K+YFQ
d2i9OeXz/VMJr/sUOx4gvFMNlOvUxtb1qEKu62R9yON0ivblHzzLVk5LQ4mgE+Z+szLPPo36TR3H
rMGKqAqJrRf1qcrj/FGUvbR+u+C0XMeZANUcuoQFXs6R+kCKqjnnrkpZVU1cHgRjCgtDExNmfIIh
uhcuEgti0YziqNpc8YJj2wzo0FZe7SL1BIhrzuShA+HdaAmuFccdrKenrQ4sOOUQSW8aGQcNQwNc
4cZpNOnLlZ0T14EH9/FVHOYKWgZdm+a9YWY8Tx25WSOAZO2++HFe32QAk/QXM20ir6hF1A04A9KP
VYCNzl8oL3zfhDY3b/4E30CagyqVaabdGeTFp9G2FPacR9Iy9tOHt5aIcVnzwVK+KpXq3Ub4hGqP
ix/rxHWCaOtVRZIZvM0HWcAyZZvmYQsS6LJj8QH1Ljc/gJ8FShJzN44Sg2f6/Xb19k+qRA8fT6/7
weJ1lzpuYuylTRXqpzq1bL35yLK67fY0IfC6RTzhsKBX5l5LX6NcosxK4vN2SvOfo6H3JqfCcLR0
zDUG1KAT3wdQzbJT33Wpu2jM+2c+SGw6mTV2pYlebnqqHiWJP3vaatXWlFTj8udpScfz3uQKu5wa
6D12M7c/zxUx+525ecW1BPaVcrvezhwu1xnm+eg0o3Fx8Gdm8om4/KMWJ4XMUCHffP/nMJO0E3ik
8StryHWTvcPfPs122q/gY5rU8KLLLICaLgEPHVAc0eIZr2zYH11s5gaUAYdWjkw5ym4onYABk2fU
c+LTixbXG6Q5QUGZeZ63I+x3qxUv71X6hgqCytT5tABDj8m/DhkHRBfR0EN8sGfpKIykTebx16R0
kumLizpUcyYMSAbovi0RxIPD8Gf32JUuSZ4Yp0Cfo22vFxmlcV05aIWhTJelyX3Ewxbzek9dxvQ6
CzaVPmI4ZYpbgsf//GMNx/P99R6pgnmUJ1AaqRXP5veyQZ2IUNWADIhkUEKHBfuLcATdmPfVlA0D
KyEEth1Eix7+vlgcMIm21wLe8FOBeUXy5GzBKoj1TjJ9yvXlG1i1BzlVjzGS3rik8tqvwmyzfyMn
FCx04zucEakCB7F01TjPNbahl0xw62PYxnQPyne31G6AqbeB5AE3uMdR3WQt5JuBsDhHegnVyp1z
MraUqByVgGiZoPLEk8CCMWz4D07dajQtZXNv08jaOwQTDDd6nDZp22UJvj07npqdFMHRvt6XSN00
JMRzXK0IsOSVWBdOYtJF5O0RW1P1cwljTeLLk6ovH9T9TEUHVIAslPxB8LelziMEsVgA0ziYCiSD
rVghmhsm/pY4cNWYfs4bUjIFe2dz/ahguIsHNcyXyvNdYxm1xzkdggpXRkcj09E2UWJ6vdEX5htR
b+Jk4IceygkzIYvsV1Qz9Jm+pqlWSbcLTw4EO/b6ypjN1UGUUqRPOqWiVjb5vth5s2FHpqNFqD35
v4ql5KaYDcQxzYUMT4t7XS2FpIP83Gn9hAWwzK8cNQskwkdHpP30nzMf6HriZlhjuT83GHAEyeFi
/NwnQUuagiGifiDT9h+ki52ojaoU5h6l3V7At/6vczAqMiIfPjEpOo+NWiL+7gPS/nmk8mQnrBG9
LYksi/xgJVU2j6xX+faUvXOnwqdfUpMF0/OMonHAfqEi97TlS4YONZmYbXRbtTDdAyasrHzvHuGv
/L66CeDdcweh+uC6ZB2bqZPgZxzswyajQG3DamsrekiQNGkEa/v6BXBx/7XWuuWbxSmjfeCaG3kC
YLCrTHM/vtVcHxs4L7hYGz659Tc6prIKfiTuO7OZPVB+F7mU+c8ZHZrrm1DGL6A54PIU9fOZfmGd
ef7E8VkA8hk0uluILFcaY+0flA/0L8BHbJ0eDGbs19FElSDAFRv2JO6fzqAMev5WYBtHOJro5nad
gwBoiLx9KrVBUZyWkXLlpqAjbXhpFvcTwUEXIY0WXy7iEmmwkHwrdoOUDHRHfvM2LlKrNHIaMmt2
xpPacIgx1XXNyqWdNQWuWRZSygEHlcYLlHRU3dYPdM5UiNFQHEX86x34bn2ivSrPY5jZiDcgT6Ze
cQaNbrkovSyoHLwEROikXYjs4KNu8ukYTYsgRYYTOGGvXS9kJe7S0+nVYJHY7W5HoTsL3wFBC0hq
2VS2b4V8F+MreUfR/UjRX0HWVJVlAikCD/5W4mBOekB8q6WQKiT+Du37f7byoawE96PugI5UED5x
5l5j0XbaUu1QLn0yDPLei7FGuzKJsl4OKUDjBroux9UIUiHx+Ya66C4vE2OakdaJJYCOHy9qFAxa
rFW7gNFGw8ji824yMQTkfYGfTE3irEs5yw9NjskBlwJqU2YIBLep0fVHRELVx0lxUNJ36WWfwNjW
anzO5Vgc4BibYMhXUmhFIZkY2L34ulWt/HjQqxlZ0Te2ZnCNpszu3SoTdUBjgfCM/5G5+v+r8i1m
SQ+0nKVHoupT5SPHXzxnRjBmoafnwRSaaHZfgU0x9pn6IrS/fzvvJBOrYKGf4IIR7uni8IX8iTyo
/zyoFS4yEbYewJxItPx8QRxBmq+COtJmSDnFw0j6pW01U8AbwlMsc7UckKAyj866ZjVd8EzFe5g9
4gieiFYra4vWktZcdj3UAbyiNW/wthjc6S0/mhUW+wE9QX8Dyic/hBWfznM5LehEKOFyTyEb8Lim
dJdweY3FUSRAJg8mSdZbvBbo/nOF1YpNDxQo1Z56U8gaueWtB8Dsw3kb66UpFJnd4aGzrM886enX
O1udSmDRuADxr7hZWUn4I8uyKc14T6Uh++xf/yn8poo2Q+huuIISEp+Crct74d5n74AXIKRGyDCE
ju/DJ+Qc1dX6A/vlyliwSsICAZz7SbX4KHWLwGvLiyok1Fbmso2L4Hb+5iKVwQAGvbEm6sOctH+O
GPAu7d1lOmWe7tB/YSCSrrFE1SuGBza87DZ5yD0SuNtVPN6POhGldJLBSm9tBREigUpdBhyrA3Y5
mUZfRTpkZGgQtO4XYQ3rhl9DHvjSwhU3/03uB8Dt/X3oL7X7m6zyucFZ8ED42lyMf7n3GJ4LtFZt
qWyYwWO4QUWsp99AWYs+/XJkL7Jj8z1mDU4kzEqWQ3nuQLpV9XOCkcCn77MVMweU9NcnqTsS8N3k
WuIGWpQrZysjPb0iGsBI/rH8v3+lwdV0g+KxnA6A1kJ/v4cmdhJRTp7v0zitm+DR18HX1X+La0oQ
nx6ZckI8QyeaY73c9zrCA78ZiTGdofxuoxwldipLBB8t/rUfVGXSZUzTF7sgQIRXW4E6T14ELQ1f
0VSoOfzQrWbLT4A+msj+qsOe4lOtskOcdByw6OqZhsF2AYSykky19LDyGfhpX5znXF7QVsH41YIK
wWLLiSBEi/b1Ff9rBxZ5NM8NFjWn8ctf8p6CXYRPhfubaD5lV0G7aYAv+roW3OriP4MPDyzMjq5P
kn7FFsaXXJOy08/MC4mXf+FQeSWNp8jvt1p5kmrq5beWG8e6sc5gJsFOJYdJ6+e+kfba6xpoMt0i
DdnnXML83HwIy1J1EQM7i2YpV3Kmwug8Sww0Rwo+5Ps592dhbDdswQQ35O3mrhxfObnP/XwbzJ/s
f/xioGALVUicbA3QuDSkTHX4XOi8kP0TUtb3hkM7wiW817644fT10NchDRdIiedRUlQ6YmsDd0OP
uhyOpveboF03MTmWZutzWp/uw5dv5YHhWU4SZDWOBtrLOuG7I+hj1Vo/PdmDXn7InA2ZRYYxUehn
M0G/rbmk4tnlGl4VkM5zktX6BJ7mTzbwBPcj8WOWh2+fVbT9Aru0oszOdckJjH7Mt2FHi4Big11y
kLn7M3M6SnZUEfpxFZ70ig1nfy9GbsfzVzCVj59RofTAhGYOwlpv1T6VoPqCqKfv81PwmkeWfCky
rSXZdefJyBN9z5PyEaW3zhlUoJm9ouVMLJyqmunBS2MqCCDdCl4Kl7AWt0K4XltJu4UApgkCrnqC
9Dig9BCxdl2sy3u9XBfGTCIQnXGWbL8d/wwfiw1k1VD61WLFHlYmfAUM1dMPod7iwvz5HOp55LLU
Zw8SITQ69kAu5OPTFL/URGvaiYvUUotIm0RSSvfiORuN47P06+1eCDuChMiBTShohcZ0A5qeVyXZ
UevMlqIXruZZBic4tGx8GODKcdkQzbTX4ulYXsI2/FBbubJ5NpXKC3Nveu1dOCEAloFzDcbTnxnd
hKPBNcNWn/GjjP3btOURlXHkGzE4VsZJOwlDtRAGRl+Io/J430p+8hmFxdl6IW4z5xK8XS+YWCYs
RLj50Vw+MA5F3+YXpXGDHiRRuxyxoEd5uoUHkGzAeZPMTmETbrJaDtBGkspN36OCjeb/qntO++Bw
qkhQdXzX5uxGcH6aZKsfAHboHSTGZfRVFoGiaAZLenL6IbiYlaF92+tGxg1lhgjkJPEGVCIFa+4x
24rNM1MddALcS/v786hgJngo2meiX4zkhvvyt0HkUW841N5blqwH2UAd5TabNIaqwvdplNEZ2McZ
kWw0PXvQrk24Snrux26e0U8amJgxxE9Gcc/N46Us+9Vvv+4DdJZP2NHBKDZvUVZE7maw4aZ0f1No
TrE9ZZ08R4CcBsvdq9FplPiZoqTFmkHkQrL9cxnmi5RR5kl9Kd8PceXn0hQmQ7UD0UfuzsmREeIq
c6P6b9OjYYm7i7HFiacOuHub9s4GBguokxjgaKoAgrqBk58ZtaSuOALRSE6qdzitVHsQ4brpvIGL
pIvkBfLa9VqnvJMO/Y+3sj0HrExuGMKuYTeXtmpz//MDezPCbdGZCrUsosR6puNRky2QC12Hs9AM
lHSdgwJJX+nesQMJlHgDRBj36P2pZNiwNvysNB9f0CQz2+d2PaAwfHLHWZULr//c+uLBELNqT2AC
GLIrnVTEwMz4Tz5lPMCaNHzq7gjE5zEg0QRpChnnefD5QakEyeAe0F1KURbOu1NhFo20ARIguIP2
d5jT1hlpPe9F1FuSE10shKI0s8lJPJIljNbAG3Ogah0emjxN6N5bwd6Pu/PfWxs0X8Gz1jaIu7oQ
UW3MbVUSO+il+FmaIt2v0lLnLu37n7x2k72u8pXWdvjXPOqTNql6JzUfY8wb2cvFYNH1Kg1Hi2Q+
WPYnPqEAiOs+r81+0iwCwGllmXdY4npLoXrwYGLRkIjQgfj1WZiNOs5ce1xM3LL3dRkB7bnlzZBk
/B2JUXY2D+ZAjSBcy1j2ATRjelplIOB74LYTh2ZNXTOvibcGDovtD2k7DB8NKFopy9I+P38HGwwc
p0FL3R8rPi6h/GFDSAIDGZLSYrE0xF7Gym79aM7MzCJXEoh4nUZi8MrgWANbQWTKh/ZUkP06P4LJ
RS8OlbZluBYanf8tkJlu/1MSZRVxi0ClQAl1v7/WFASS7UaWh+CCBDF1iRAqUwrDotzyhI3GQ0ad
QwSkr9utArMzizK9cutOW4VQ17bGp82TzTRufJlDBXpjX/Jo3+9B0/G+ek5Ko50/TMFA5SV3QdF2
iGaj6ZKSmK6mPdJf/UXbC8gwB52+yEhKFsWF6i/7kqnnly/zlG21wfkD18UkIMOebuES2+CzvoaP
LFqZsAbKGngaZkbjeK4KqyfGzg4wtMa7KAd7eVfTM6acnk+pUHAKyXgwAWHjDyOb9hKp3R3PE7GF
2jU39jMGlqEOENrfCFgZNRwOfxL2v9t8zrlENt6yM7Psp0hS72pCQ0b6IFNCYULSLUWoDn/66A9N
hBXn+u3gtzCscWWlSsFC21Xt9+q5+wsEWhjQJD+Rk5MvnbyRZV6pB8UfUigc3LkT6EwoO384p8bD
xeFFnq9tB9VfZcDqzZSzZ9jOPXr7+pW2Y7SVkd4/4ccUTUQpRw9cRoUsl1xLIzzPyYuiSrTE9ld9
+TqblMf1BRtpAtxO9Lm7Q0Yb+STx1NsWX8mKq2IbFDJCpHUnrpUx7KPYYdTQz02tO5Cy9SpPHUk1
McMeM+YZj6AET96KiOFmuaqICTGSxoWqMwVcjnUzdjCkeIf7eM0i+bTrBseLWY4a9xtyNi8kMFcA
IaOFBQv6kWbw1DFL+yFDcZ1B9qPXoG9o3I3se4vHmU9aIV/PKWWBX/I6OHaSvPxjz79D7+3GAcA+
4fHjw3FSBUwx5o4nSErbhw3h98gaXljTIRKR6fNQKaGWazQUk43AyZ5n0UnSDxLbNHdxADrE+TFz
wuZc1DPzHYJi9lBZUxGAU+w20IMzHCmT3LrOcsKK/SBzv9HjYC8Xa6GoXaxAZ7G7uj/rUhkdTQQj
2GRdl15la9pw3n1tfT/WrRlRnT9fggCC7+EJkp29bAS9PxPNxko/pPrKqYEzflI4RqRAtmzQp9FI
YDCPk9mh2aLxZNPEbuDZyaPIWXCBgabzIfPRlquEAfCbODDky/gX80G7xPrzaiKc8BBhoOQxstK1
3mj0X4qvhKz89d901rW57qrAGZ41y1/k8+Zp1q1dfoIMKAZ8pgN+UKK1UwryQVunS/hGAy7+72JV
9kvuoqgrXafBRhHlKdSq7+kHxaUC3APvyt27mf3p8FZ4RDLxp6nawtKSpZO0h/paVjOjEFeYkuQ0
JhB3YuUeow28j94e6JlmzJxOqtImEIYzbKKwE2uTz03CKlURWBXHlEUZJQNpjaO7jUDhVvLNLfLr
KNgRRLwa5mkeyXX3Ho39v18OSgRt4D/TBD1hesmaA2BmYWyS+7QX+2C4BXuTmKHVqvDQRD/8xdFB
OI1Ao/1/8yiDUITs0bIcE4t/4pzp4uyGl0M/cVzFifJEMHng8SuX0tHwvKZ099SRjJzMb2Hrhjtv
b+f7fLOgeRj41QCX0R2IuDbtc/kWihD3XkUD1XuSbzYYFARniyeDkwIS/eAMisAKURZn95uJWBE4
MLGzxFpViIyUhVaYrdpif3AS4FMrqW5xVSJk0A1ekAek8Zwx07QIuuzQAZZOtFA8tDKfdRmmxM54
Z8uro3LIP7fe4dGcRD35YFD0ByiSTZxTe7wRxI/E9hNqPFpoqds+P4NDikfkZ9Fn62tZZohLpNNm
v9QQBGMwd2mkTihSvcsRUzk+aGfJVSmdNLMuFUnEgaEI0bAi8RLxJAHjxhHFcFuVGr4QnqS5mib0
zDhCv6PRjcOo2GeCygfQoMAGWNiPJegMWNQmbjZK67M8S1azW3h3iGV50EOdFduWjSNubtUV+qmA
Kvs8sQaCxGgqBAU3nw+cP2SO86VzcpaDcGzN6nP7EJJByatVB8xypBpbfQTKH2cUjsWNciZVt4oX
2pfyoW0CHTDEhN4jNs6VCnnTftNjmjfCSeCSg0zhq0yDS7RQKrO0/Z4fGfvbJW869Tz/88Sim3/g
smb/6yB8bXuFt5kpT7+Kc1ClUvvwJkiCJXB49EyljjGXod9yXO6+9uYZjGhyuriVXdHgFNxuCVv/
8xzcZ2xDcmORWoYxzcQ5kQJzPRJlU4QQCmOnMqf3syoMzBKKzuu0+zxdkfHDE0Wrez+fwU1WJlSa
uOSqREm2tDf5k462mYgGxvwhFFzQjPdyjWW05brv43d4yHLsudkv5JQClk5jVJnrqZbIyI0aDVmb
AEg6eVtexfyTGcOZhqqrcvQwQ7uEItH2ealj2eTMN1oeM2VlueNnQfd3g1pPN3JfTA+okxpjvEAr
af/BuMc17VPjdFVDF3szFCZlKjOKloIBhSQUDPAQGLMo2eBFJl86gi18Eys+G52jyp2XsIu1rcCd
Vs07ERfOwn2OgPik76+I8ShFcl44H3YzJpR1sHTGHdsmDaixahSbHgwm8QrPkkEm+Us4+5Zoj9uU
tTyY1NpJsuxYKu1Fkk2oGIW1od6NjJwVj0yssgOzE4sBuC/Ew1bTcEinKxhDnnsE21Io+Dh8yht2
jtxsLBOisTMbXL8wr4vRIXFDBb6RI+bfYTUDays7QDPRHspXCdi+ceL5t1RZgVgV6+TkBxYYqPVQ
mMsYOI7F7mQolFkXaX85llT9S3jF+nXLm47+oG2DeYHL55PT1KlGjky1IsxQIsFYj288wexKJPmO
EyfbY58IIztvoir2vvcsaPBT5CQ3eW/LD+/E9Txm8ayhc21wXtQVgiPkjlG/Hjj9dYGoLETeq4Pj
K0vHRsn7xMYkVCtloTKkbu7uwwfLrEN3bOnS9TYxLpeQj2ZT/2b71aSGhUIMHscncYr7Lj2zE89U
YKDPRF6i6ebD2GBKC9lOtGM462umh7CFkddNQsCrXYJ8Yg9rrxDhR3Pupm5elPO9GPyJEklGMIai
SEOjGnMvZg+SR448kbIjCXVIa61EGphSJz2WRZ44SGD1pLHIOnzjF8etgd74JpatfydqUg0b5gpv
PlyO0pgjZL8lBj8lYZw2g+742rN7nkS7CgyYOKlixiD/aBGs8YEl8dQvFcq7Xb0HPkpjjXpWRM90
2Vu9nYxk5VoAou7hF2+EXDYWStonhK6m13vYfBfz4oyQKK99U5U49J8cC2XAQLu1f0onOgzITLP8
gqZe68AeInLLL2b0fQV2z9yVQ6qGI7pCpxhaTTSXgyvL2ZKGTFLlYZwZNGaw9+X8bbLh7Tn7pVa0
yvd0srs3HvFXkHoJGNud1WDo/knztwSDms+rcPjOin0YQ2abrIJCD/Hse9/Yp4fCEEAfOKVNApNr
9vCVURmud7qAMkXJ2y5lfJAvjHbn0oxoVDQaYXt6mNo3TbohkSclA4BeZixzSvOxy7ABWhci+1JB
fuKqQ+X6lwChCNqvCEDJwdgmirjjMemDT0hiHl5ID0KmgunE9cwtzf2hnH1nfNiW5MB7XtIz8cSq
CtoFhMQLEXvCDU05Jypzsyl1E4QeLr5Etpi7L+9t9KXwRpEv6SoZZ8BVcyQHviHQ/gvn4SdA2zVo
GK8NRzgAEV5yNmqbwnJCFobO+VF3LOmIRj+fD7bpFUhyrffXLp7HnHzF2N59mru+0ld4VGZzRqup
5z1aW7kf5+zEvi+pnZZICxyNO3hj6wju+LuV7LQN1tDhHYBlK4Md50XHsnbNzdGGd6YJCXgdk6P3
rO9AWIUyGVqic8mP0BYg2XKha8Fpo0P6NuA+OxO2nmlaM5eqwd47RRxvM1sjC/ir+Hj0ohzSOrFf
HRJp/8lxJXcco0lvTFybZp6f+PKCgiam6OSWouaKs9tmqV1JF9FqxXTnFmxGKaN5hgiKGlVxT5d5
mhvqQGYj4GHX4chvzAFJPg3PNInk4A6mFPWvdH61OoeCrhS8ks3NBy0NTmthcAoiM4t6QvmXJZNI
4UGS4gYzShT0G1r6jGNTzqNDb2+Uc0TZVopCcyNXXn9pNCfoyLTr7Rh+Uk0foAdLcbIbt4sKxCnD
jsmArS4QbIHBLPqkliAYUZweGrvGyacrMws5FwW06jD1vik3Hqo5Xqab76Lu5pb8fvZeK/WaIBX9
zdl3YiHud1ODGZI1FYL3zOJl8m+i9RsasZj2CIPwx0ceCACNZiXz2cr5IZZSjVoFlY9V0tWdkg4z
w7qTPrxOi0Ei2yZtMAhYPY9YxOy9Uw1OXYJG9ay6E5N9L1rcCAOPk+bOeQh8RuotOyiaGyDU5xuF
sYWKuMV06jNQ15YgcKxKGI2yMVr8ZtuSbomV9n42UjeyZ1Mmq7sDU9hY6A4g0n0qS4fk4wrgBWrD
QLnuRD+rTHdW6nwvOXc72x+Rss85LZPGazDFKglGEAheqyF1z4TIi5okgkaKk4KoaHI+TEL/9NDa
UmODgSQ7VbBEQ6NmfyHCZzCZue9EEbJFY1X4jZLwic9Ee88to8LB8CmmkkQBWh1VczpUj8UtHjc3
a/83eTZnkHIF2NQ7V3aAlicA9n6qGz+F91/biDn2XiM4hqRSuJmGiBQY27IUBmlhl5dgrRXnG7f6
z01fm/C5WLDOQhiSeoWeQaF4yta3yPgGpyQA+xTCAIliB0537B/Cc66EdTmQYeV2zawOc+Iy+BHp
P4O9BOT9l9OCqmFUNP/zv/ejpNz0gTeoLGmJKtwPsixWoYEBDCxr2udjYlNXgEWDB/ApDI202LMC
HSn3sp8cZ20Hzj4gxgE/78lMXr7QP0VwzvK/ox1KHmnc4RBtVEpUtW4WEKZNDotu7kuTcJWdGQLr
0FYYWKgVOMHerHQ6FzK2KELqr4MUGmuOXZ/DvGiaLmFXvyZSHYHI0g87yck6NQvQvIoQY/e5pP7c
w2GduTqMXmzql1zSyITy3eKL9ZD4dIEfhG/ExTK+En0V8gCgBd737o2bljKHXaJ5Hmqwr163aZcH
b0qTMpEkBhj7zkLpKFh+q1NJANuEhA71xKxSmauuf1wA1riLWfaFi+4lsXEkCmBbhbz+nHoSZHKw
1CG9Mnzo2oRb8CET2Fxm/Kt4BMPQJ8j4vQc6WK+NmLDXxwB2vvuHocyPCEYG1mxuhSD/lK0XIe+P
RskcfLnw27658pVQTQ/2YGj5H0AAqbsbM8vCk4TYbMylSEhxPdrWxGHE5O/xMW2tUGyLuRWbToL3
R1qnCCVF3lHroVBF2xdH+aUv/dSwTSiMqgIlOSDn7ZLZm6vfIGbpOw2xDdVaV7+BdBd/gkxfIaXX
oZXfDkNzE7WLh2/k5P5afSOUbRKdWNzLAKvJUTL0N/H0MspPSQHgUDKFeUHqaFLZBeT0zqCr9zo9
B3K5EUfF9jJMiU6LxgLkgbFjZNashDtsnAN1c3yIqo9QhIi0Oe5pfuCdQOd/dzrwHMYFP0tN2+Ss
GZewvG1R9M4L51e6iA8Dhy+cSmUpPKv/ECSBydD+W9l9UdEnDUJrRnWtC968fUsGMFQFiAR1u61p
zoS9xMtCPZ92OsK8bLFTZ1ux1qw91CWBks2ygD6gzq3LzQrG7owAyaHkr9xnxBppCBneVtNvtQ4X
apx8wq6TX/tClLUyY0J/jDXHXgoIWJvDn6y2njXGLBI75HjUIKoWfTxNHOVmwbYjiOmDnfUhryNH
ldHLse7FJls9ig0YQSi95wG5jguMC2UCOS5Z+dwFIQ7gA+ePGCvq9IeCg/NeWNJjuQYCPCVehxtc
HqlclgpFjJkqe8FmW4Sy4pVT9vWrgRqpN6h8lLcTBsmg5zoadnRN3t2PavWZOLcnxutNM76xpzAd
ioID62/ymIap4h2IH/vyw1ly0H0eGggp/jo69FibfyDR/GDq6mkEBS9y0R9nWF80tFaIcYYjpv9s
plsQa+z7ipaldJAbiCYhX1VGEmF9BfvW3oicPffwkAH2k5uVawFnExOeMY9U/+Z7QE626tjIyd4u
kuXeXlv/tfPnQFzf7pqDhTJsl/8zPpbjQUkAWGvcxgUj+tkfnPmVLB5HNmLev7b3IKdq1uBSVIqD
GzS5x2f5kG+bP1nbVrr7AzA355OzrabfXfCWTmNTmyhVswkUUrmjWFqEhuAL++xhgmSQIG55PcSN
V10SVtoTuH1bMQXYe8NRJix3w+hoXRpEm9OhnBhMDhsmUvU2fHQ1FeyYub5orflwv64kZJt7RyNq
0odCOB0Rit+Bij8SsjQGD8JEWn9zuuHDlbqL7tNrv5mA2S+maNfO/iUxR37y+vH5FeYV8sowvm9W
XL/D5GJKZR4gVcEac00TozLIFWAOxQceetmiCSyj2ouql8PFubZogd0MEercmp1oKzDGm8Wwh7SM
mhVR/GUiYcKdpDV0XbLw0j7g+rJas7jYWi698POzxHT3DttEW0ww8IDUHBlgxjh4AjtqjF1UKu5/
QsfxbQNtTUDv/gVTPWDq6+FZoVAiERUXDZ0sJisJLb7SaMS5+9WXw7KAbD7ONuR5nhLWoOaYL8DC
b0nny2ku0l06UwS+uvd2SpJNN2gDk5oA4EaVXq+nawR0bvvqJfwFZGlQlX9mnOtT0ay4lvMr7QeN
gR+hPvyoplzHc9MefyWHXsk8/RVgvoSdM4uSFeQQ40PZcUig8kEIj6fZG2rfea/p5PzvJukUVam5
F/2y/80do5/sUIXer1QM4TL6ZuQkYrA9c8SGiXW5myKmFE1x5m9Rq+IqxrFWJlslJYPxyknB79ra
2oXiOtHhiSPCoIAdD/DIPA7w1HJ6JO4/VVqFivP7CyAQJ6NTWLG+j0g9dsLcCwQPn2IgwiT9bifS
MBSWKlh6JePP9fDDqdtWiqd5xzkKMfOYchQAtVAY1DqcjpqaBu/CvshTgY6VI3R22idaGKT5lsdX
sgOjj043aBX3YhDcA+sNeH0dmG1lopEEFphYnCb9s6iCwaTtDiyNVDdHwvEACHvQEKmfXezcDEjy
VGM8d64wG/k8/aC2eKnbSVS6BUH9T8DrYi3cNazPfMqzp/klVeJjsI3OtHo1C3xyaC11qgtC/vhV
sYNrnO/drv7Gm4j2EBlVe/qxbVDWX2312C7lbrHWSn1Uv9iLy3QstS0KJSuuF2QLJDiw3sv8TqZZ
1Y3tJcK0Rz8o/2utIy9kTROXt6jgmhmFWe/R1KB5/pLJlJyjfxaP79UUda6SmFYnqIs/Cd5PNqvL
4r8RhTxYSft6AEy8vBt1kcC8/anVKuDzZydR5xZkEadiDPtDW9zVVFe+F8RrZ3oDwwQfZ+t4LBgb
z3LuhARJuF3Cp/7tX+EVm0tNne06OeLIGTWQRGbd4Vuut5aIqLClXP5Kzkp+HCuDwH86H/Xspk7Q
2Ii73I58bG/zyljtzZRyGtgldfbKj0fXQYI4QaXjHkjKbIxAIt8uKwwGLVqIsaNuR7bBoKhrrq3P
5pF17V48raNnUAi/h+bRHWXALTG6rw2l3/t9Q0k61ZN+Hfdcad9AIDu/fhOv4pXa+F0abaRZNxyK
9E8skdfsbbbSpgqmxE8gwZ/U941ytgq5Kl5O5KnYdlJv7BipkJA34le2CeAJJc8UxLq9RqzXffNk
scayYSi1McyWlTCNs6Rkqdg08siX8KZhXlPeJfqrDkeALIgMxG1jn0vt85jtXa89DuKS+hAt8hAc
P24mdV68DFtDZnrej3pmrxMf4rL+v48Lzi7botCbGjlJ+vJXMty8Bf1gjp0zQE66CDrtRGuRNTBp
1G5hIh/+nLULRE3v493R6f2BSXHfFAdBI1GpN6Q0F0sXq/nyUKoKDYvcfHGxwahi4Odw7GblKivY
R2xtJOKeq1SkX9kWRlDpAvkUdkoW4WVF/9DWwT3z3U8RlRom43gX+uWIdlqntQpSEyyPohALz3Ys
1CfHsfY8jVmOCTMeZL33l44cWn01afWso767hyuboYK/m6hnCnGZ9oNUgP4sjnBCX7IL/iJs46vU
YsHlgHa8KFJlClIsFaI7WzjDKsnynCpZ3G2GCCApOYQrNC2xl/zs0xkzujxDdQyhYTtfZmDy/aUV
zVd1i6mFFhqCICEVasxBaX9y8srveZk2qj+XbSai5OYPO3bIcKCPEOfXFoUdMpkaRGB5OnurairR
EM/WYj5u/bo5DoxS5DfDPLpUSm9PCbNSI8eTK8H6iItgZhSoSCrvhhfYV3s97d48dVhT55ngK6vO
SW4zOrEI10XIMryL/yk+4wDovEm9DbtWO93vHCaoohOpWG1KdtaXABmBFpDfHu5QtlHZlKHFgdtK
silJEXnNk6JkaaJdH2bQfr4OeVr2lNKMoRNXy7GTFa5WOng/UKf+dlxVW9xoyNxl+KPaf0Tw5jo7
UoJWJ8aIAeYDLtV29TEslsnWeSMmDYGcJyE1HkGByy2Oi+s9DuzTpPeW3VrdtPANpHc/3cIMRSyW
bMaU0mf4rtOtV/lO4hw3zg6YxCPtY9bgOf0qJLN90p65Hce1gBMp/Rvpg6e4HNYoP8q7wSv1SMb+
4dTWDnVP8K120RAi0tHDe1Idm/Knb2sPGlRs8wzCrAojcbk1suDX8XG7xz0x5I9l6lgVeBiKLXp9
mLx8n3D/PIpE1+JX/Wn45xgfSR9ACM83+ttAD5E9DVWYXeQJvNlad4fgWMblyu52HPVvoW+QTkXt
+25BLiPZDod9ErHXTg9DLOrCeHwP9MI2OYp5peX+Cl5ZelLkg9TUb2ToTxRpDJaV3mO+Vvryj0Gz
FDPOZwJwpuNCq8ircpO4d8e+4xMfpsihrE5eP0qGz6cPIi7tPMVcGmGhLEuILCZcT2+laIEaSB2U
8RRdhD0cDHVeE7h6SlSBmXQSGdmO4ZKa5yWXDoKECkizNsLRUoR0xToT29+Mo4tvk3zfmrtN4e62
mVY4zJTSvzovaa3CdPPUnFlXZxqrr9x41nuyVvT+5yRdJcMzuUracqYUGd4hLsKLOKddDxLYLTI0
7S9XWQhFuvTKWyF4sCsX1lqFgQDrWoKL+BwYatAAt1Ik/8sWJdHv4Pmo770Ise8b9o8lbWgLUkav
f+sjDZgODzSXfCK6DSbB5MdD6PPf5RVLtr00LWgYa5Ig0XAJSMWxwZDTO/CtQdIfweA2nuo7aiMU
jTrZRveFH9UMufbNw+IyuPHKEHVXB66EDRPBDxFMSKK+f5OnXHF5x0B3OUQspT1cO9c2N4ryyYQj
WPfuWbZ+A4eKEw/CwTfz+K9uSgNXLIRj9OhnTLmJG/De0dgQG5RsFtWtHwR4/UW0JolY1XBMzgFE
Sq8wmOCiOIfvsB1f8+uIl9BEjPd4GRACEjFS6VuvabxqkLUxnuuXjud9wdw52a93ejm9DDwmbn2W
TQkhrBVUPwt8PXcjJpdT9426oji85v+mUErMXhvklVu18ju0stlKPUyzKbOElqi11k99fNPBOvkp
NeEPRj3n+C6GhC3FWnZx0X+SdVKn0hXncU5vTESeyPn97UrwjNYgQMAusZaGiqiIY06HMlZK0zJ7
xjFPpPGLv+kvsXt+UIgIdvDoxcoOPGxl368SrTU9S7hW3oQxG5c8A+kc7bcaRQL5idQMIcygli9P
X6d1n+bS7uFGQBgVGw6U4cRgohpfQ1YgBnhN4HsDiCSeBFSAVFC/5ad2+5U2r0GK1+DVHQQe/Ytq
D3vcdWIc+s6JSC2keobsNwDl8G24RPZHaneCGrC/yLAbhiP+XZyclslUC25tfONhDkeD4nhD/Hc3
0g9MYYndjvHQMd0c3geUvT7jwIGsWvBhm1v8KMF3bn1Y/KGXQyZxGyDYhGKf9atuqE0mO46fNkmo
EAEuKlRLCtTkFC1bcAeWPnf4o9oNN5ERtV+A2rI9Qf0JCXVS5OSagPpuu6VL9+owo1+bJmY5+Jf4
qcael9bZTtgSsCiCGH14Hd7qkLU1KWkiT0wFWniL/SttxvTyXXP56OI36WKZbcVaSV2SVCn5EkVD
prh6WYVq+O1EUIEW0Zb9IP7BbY8gXPVf8xYG4GmvoKEoFyfCj74m8EPdUfqhKT6wxD32S22H/0Ro
pHWQwLAZmYM5rIKDMSvoEZfcwdGfXGEaT1PftV5P+c+PMWgydHwopNwv7fN40X+HoL+V6yS+ntJv
7SAM9GoExPCAQCHq8n+kfhtfqYjI+mEVjsiq4BabTADA5gokTVHOtOTPEG5XCNGVLp4qKs+jqnPd
Xh1V8I6Uc+w759mJRc7dfEFIm7tYhbGUpUOi1RNasXwyj3zGBPT+b5loS2lT/CS8YYPAS6AOYTv5
z0EdBtqWAmE5GSp5v/C1NSxqVFaRjO9hRfhgRV3a0LBJ0vUUmLcm2JqW5prchIY6bVnq+OmBVPDH
UjEXcnu0RFMTHDTwIBCLHOfD2Y3JET8bekhaEMnR0e31/fzysU6U+/LX9rH7mm3hYL1iWvolMhx5
y6nFNUk8KOJFVXacROtn0oNH39ZKfQ6Nz39nZJ+j78P1p1vPePKey3OUkzxyB1xEI5PJArrEKloA
lEoNKfOS74vWlkXldyfLHG6Cti6HzbQKRRoO8+Bi/lj+CWQJ7q8JwU1ry/rts7DnEa32riu2TEF6
cRq/kdNTujzw9dwIp6TjtV04Uc3xKCGHLlTN/oef5Fs6luFQwM15WJsRqgdvObOoUkd7h9ZEce2s
+AITQw9fi1tU1iOkN+MoGThnzrTOz6rg4c3tS/M5hcNXRrJfnQ8byciFtZTiCbNoffrHitdYS+1G
criavR7LuM28ZConYU5ggh8SPpjKJadzg3kkJUoCna0cTUVf3KNBkyAG6I12tlHJMTO91si9cX9X
+kXyw0RHpsuB2hf+Gr+uKMQhu1ZHvrUGQFImwHD9TtODz14zPwEyCu3vSCho7BcfTcSssWHPoTEA
dBoRojau5pa5sYJeTUiEyyYU5gApUHDzUTCHJZJcRPwH/BOT9x7lkMXqraY4ZKtFNB8uaVUoxpjS
JZpf/3Yja652j+PucltUT3DM37LTYUC+gTZX8+EyvkGfyxE7DmLELp1bYEbocE1mpHGvuvj7OYTR
JilW7RuiSwwsZhywIAR0Sh7jhxL4mcnQpVqRGQd93R801r+4ljD/7lA8mnV2Hrl14hWCD84DzLtz
owJHXq1VAXFNHJtrEl2h91lWk1SEV7vYUiUe1OOeG1PmcjQE20ngJ4c/mbp0BUQIlxjMcr8IyF+A
rssVPLQPAtItUDUGJbrPIJZwAqKlO0P8VnWBZunarzWALWpcKkUbu2img7A7Aun3VcqwTnLslpPO
nn7sPSq/eaqhA3LNYLam9oR/wSbbvUY1W4PrEl7UsGTjDoycEb+i9i+OJ1yuRp04uYOsRJ0Vg6/E
SLiKIMAeDEFO+nVo/xsYs3UZ7PS/AFWa7gKs0Cevvnz585aOF5c7WZayLCyEa+4UWixlSuqHCQ8c
oQoFA5sZWrkQGbU/ZKXQjslkVcMfWRZDlLdneFpM/9A3maYC5m4q9ndN14bTsavaaj56/B+Qo57a
YPdYkq4iAJYGlXm+alTyiU7SOnoU2brrQLspmiy2chAxFgmCVCcN18Y/qacjSblqgQnn6tVv7A+K
8ctjn+KGfmB+1/iPtmnWiXAZi2lXUZrfPWWtIWD3enmhcoCEQiOW5k+D7/i1o3EXzlbcwwYxEzAt
hwRbBiR562K77Y1u3VovYlW4e48XBadOEhYIyv9ufG0xiWaGS+OptsDqeZiIDqs226cq5SEhjKQf
urs54WdvEF2rjdVZsDnA6EbCT407l+IHjCUmrv+9ZpDpXRmtorMejvE1yRDwizmGkCmlgPyIkG8w
FHxy1cisNJuyoRIUD+tI/BRDn5FdmMSXP/XikhrgUbkdldklC2VhQi7RHe/SDNvSkIEpx73FJe+d
ew/jyMjoSHAqC2UW2NDnN/cUvZ6EItSTgJTYW608zx9hxZcS5UTZN1FQEyxI0cKvYlQ/TeT6C798
m3osYtgYrtGQtLMfMniTFgTdrYQ+qOCTmwNRqVTeQKpYQ0PEe2sjxyZeRSdM1hZqAZz/iqCwcNeo
QKj+xn9T7ZtU5zI/rbUZKPbNkqNa5mpZUzFEFfQvBBP9Q+8YN+ll5MyVHuSrLfU9ybF+wqo98g4U
Dh5ybe7yr7Hq/b6iWM8oEl7ImCUqDVUOdEjjt2k+Dl7wdBI7LnyvQB753sLXWKjyEcd+TbYTPLUs
PsMEhZ01tGSYNLjT2yR82HL8YOXy1rUqtRNd+HjnonPkWTQLYLYyUPyW5bm7LxbUvcw+au3TDVPS
Ga6y8yisbLunJI1q5Saik7TAGFJN/dhnUsCjlUjgK6dx9m1rBCa04NH/3VDh8Uf3JQBhe4I8UWO0
R2R7RJoy4TEf+eu1oE4XWSWUqx6wGBSdenveOeHCWVAm00GaUfxAZ9ym3wXcXq5gjHsb9/CYb3q0
yjNqS67Fg87xvPz5LlQmjOwyT6DYqhkDPpwiaktRMkLRQrQkYBhioXi53LeS42v96gcU1ZynQCn3
V4P0Z0s+EEFwGCFO1Wi339E5J6l7AYgJ7bu5cfhNcGpLhJXxI5pa3zLPjmiNiOaWZg0FWcLjsJzE
F3m+JZeJ4q72ixk8be9bC2JRwj4RFvPM/RIVhnLc92Hl9SPyizhpSm3J7fo+6iPW1P4KHxDMOr7e
y6r25no5Y0zPc0CPSd/hLVrlTmT52hr6+NtBzHrUUpX+gIhrFpVkwtH47tg6zksIA1zyYQDudbXo
ouqnqgV62oTgsuq9g6FXCoVOOqBEpIjC3FKMsGj0EhZabmymv9aIWcctan8Ojs1pyyejXDDO8o+l
msXDih425RSlV/vVRzcnH/5OG/BkAL2GlQMFazdDa4Q476Zyyi5sdOywNvc7Z7o+nJQ6yMx0kh4q
DgUKdFSRPw+pNOxYRMu3RkhEJwpyv+xkHvFh9QfuX0rj9GK2K0J/Zg8OvjR0wB1PQAYQN5FhVy1c
AVcS3kYr35kq0lkKhVHtHT6/GLmWvuZb8wTWqC2c2OL0j0MbrC6HXNgZcvBpiG12ohCoqM89s+Il
F5Tt8BE6KGyFKvvrRAnwBemwTJGsH0z2FcMrTNkg8RZ86boOXPNaNobUCqOnA99ERmR1+/E3twdL
Js6cClpNM8Y2pleBJoWbJv6G7QjpieXIR++AsZkrUqwPMjaRSHCo60sWjejdkFv8jMx9DuNipM5c
uu73bpErYBFR+IxsWOa3cedGUcePcwkiEq0WpU029B+ftDXhBBdj6lb1cE7XP08PBkNmRU2jkCjz
nJ6H4yBVdiILgQxdPywMFHplZvJtFv5U5W/RYCpeuKoDEl74JWWRUj5TZQljObklzKziks788k2F
+mY8Hdh1fJHohf5vdgCm/dH9pqq3mE4qi43LaLwCSBt6gTMBhcwg7PnW+0p32FUTh3iGTr6lpWKO
kXu8JwudnKjROrdkYYfwpcMXqJXzFOCr3FPhVNUaFX015LvbLleY8+qq5jJjes8EO4nk3N5MdOJH
bWNN8tiwitP5gwzRogxKKnfohpW4UqiXkk3Jdf4SoAaXUvPnFqnFm9E9+VfGuF7W14DXB2CTt13y
sYHcVk3gAhGFj6x2UL2v4fgKyURLdRJZSmSGhEqqlsqn7FQK1GYk5f2LJY8mkkDGR+KQVRCJKzmb
HjS6AADE/b7CVJJhOY5cbTnW+cOKnHWciP2j5FoEo7vnJMCtog7mAv6lFkSxx6q3FuxYahVDB/se
3be1S6a7iJDTTMc+y2ReWsOsOv1PhxtFR70vsNyNvMx3msT6cFho5VYe+Qxl3GEQiv2CRctweLwx
MGJbTX7iffHO9GEDTlnLyMBaqCMTGl57lE/UX11efwuPyESc1wMeAMJ+VDuUYuaPXWutTrlC6a/1
I5KjUs0T/wf7ZIvsaucfpwhHaWu3GR0i5xpv8pghpw/N9PmqeZXqg5cwEW3bEGbn+FCvaDs2wKW/
S3iCg4eh6IoHkZnDHxnHS97EcIDsxR08m+IPV8W1yho1bM6HfA6ziJNRLTWBIQmjEQAC+sePCpT7
WImPOp/kz995E82K6r6jRPmr0w5lqSQFalwWdpGrdwRQXMBa0XnDbUvXNKTQFEhcFaR17WiNUu6H
Hi2zNzRDtKFRVKoiTMwxNjwOHEfgBsHhVehUuCi9e2CydUKUFk62bDW34+85cPxDJmok9xkwf0a+
fQqCSd0lOygfHISa+uWWQT2RVRnd9gOEvXkAVehi7+CIfH9qdi3+vlrcYpwrr9X/Q6UXqhR3fmSC
lf9kKkDSlQTSKn9Y01J80ymLcQ2011lMUQy3lHz9F+RcuzJR62sRLj3+tmyWi6ltdeyjl2k88p8g
ZE8Dil8liSQGNTLsEBKSISEXyhAkO5SWjPXHfrL2BjT30t3yuYs34RN1rV47AJ+/gfyvrYnfRtYi
j7crw0z8ElWJ0IpIuXy6pdF2RL+jstzjJw9sf8+t3kwXksBtxxSq5s4CaZP9gMR5VA8sDxzQ9pXL
LFhUVlfsSHSigr5p1LZiAh1viG8gQ0PLB1aKSXISzA5BAKPrZEHx9mz3N5u0iZ6GHstr3bqFYjSi
qFtNVSTXZJ0TN1q7d+y99pmdiAu1RwIVnmxx17MrBJgqaGzco6wjMOGtBh+F0qXlZ5rQJyF7qvoA
9onRAidQR6DqmYZbPjjj8NPGyL4qRADPZsfaoVZXIOEdjSW50m9BEX86QATcNVoUadtNz2V0Irh2
6YeVswfiHX+I1atVyYkxZnwppjkzck55jkacd8IWKUaumd88bdOSRN64ya+sNNCoQjxfMBK2kw5u
TOJyXUwJqDcl4FVjyZb2GHowCZMh9pKaIiYZ6T14mSdls/ppTIxMOCZTTZiOILyS5Rh+opoxnowG
xgEVquVBMJng4MQYQ/E8mgMqLblCQ9ivgVVthlNU3nXqP0vQAxzvJY+kjcyNhGS8vvJwW6lh1shv
6GBP/LJVgW1ksQdgQS1cVKY1iZp4esgkfhbPKJNkqnqU4rz5+PFY9b5NJPqgYTkl9jhtFzunrh7P
ebuOP7E0NCl/7tveTyhiRMOVKp3U8BRMGuj9o4aFPHhT18zJ8euoZFvkJXRsMRyPKY8UDVGWLZSd
oeZ51zLdAKvGT/2ildsCra7hiMZFhSvUe7Q9BRdew+ozapDyX/0JZPt6jc4uQdLYPRwjqwpC3vDH
ACDwCpPQY+0Wb54O8QR5oCTuN5Ad/+eo/AAXA4BsKnaeopBssr+ulCTNLLz4o1ENb/SAL5G3aSIq
v657oV0IMIY24ESMVfWDyioBzvcZgz22MxGhJuWWaSvM27hjdTGn+XDjT/Ea1Fa9UOXOC1q/5F12
817EsK7aT3nybF2UbCxnoGGflD2zS2UjbS3wP1/BMQvkCKyGRlbIQHqySfHQBaAsJLMGVg9kAsgA
4op+66I65t9LkBf1aK0LMVnGRg6i1wLBFMIRi+NmKeQMKZYMLFo8U1UdbT8liNpT4q11JuHV0f4l
2FcFzd1YxcqY1xAck5xfT4vZ0J9Kxp3ShbaCOOdYfv3uR3oZxrD6vZY3bI3ARQGp66DEJ8CfUseh
IjwqfYdN0N0JqG6j8Bxeo2DnWZQjyV1WD5WIVF8ZzsZjizjNzfO2bAwMecwY2SlIA5jS/7uI4ECD
dw9d9c0oW/wV1wbAQn4/IuyAATjZ57yj+wqK5NpLdfHQ5UBDYAXz3docyG1i0RnRuS965Xq6VX0B
CqWt7tubFb5Z2iGmw5MQjMnyJrBiGlHrYsG3XvldI8IhPN3VGG2/FM/uGPBAXguTudDokWDcgcv2
7YexQ1B4MPJ9/JQjOpWHohY55Ugz5QS5UQWiaePbwT4FBkhHqkTqJ9NKxzqS2lSrN2woK3YjVg/H
TcnZ77IkSalCDqjMMLUtcwbf9b/Soct59WxhHuM7DNRLtYr0r68fv1oIIciYFwE678E5tXea7/83
EK7lPtu7DFj9WJEdjyWm513PnJmn6BULpamyPQowePsFO89Mq0NUCs9OH1f7SQuv2sILi2mdckkB
xUSuPLo+nzQcFEydJfWIJapUSSBePqvrZ+/YxkXWvmGxcNgqgPeVOsu9hLDt8M0XKP2ZmfG4WEKF
/AknjTtY99vyfnNPH0pVdXgHGKAKx8BlLQmqayN7RJJFr2GdTaD0QHAtJUwG957N8GuCMfXDMoaX
GKm59TVIOQpWnc+jdgKKPZdxfZgigvPHJphK1EFctlMQNs6wQA3Vie0utEU5LBsdGBAIOOUSIZtj
VHsRKE5Qoa4xP2dxyATIMUq+Os2Walpvx7QiHbN0Tw+2Osn+jLEiYw2YqDeUItp4mVpQzZ3Q67b2
4IcvjEt79wI01lu90TCwE/aQS+1JWuTyDGI0eBizBAe1zAf+Re2QhI/uwHPKuL6J3Iz7RKcvEZiQ
2/PMddYTj1u2twoImbITN04mcRoyJNhHUW0CmUAapAQxvDWA+iKHQnNYmzVBrUADMwuyUqTeR5us
qUo0ryhnG0h2J2Ub0LnZ5wcRkcQK+IFSQsfIw3VtU43iviL3tB8qdxRITSpjfnuv4Wj7B1z66JU2
9eWV8w0+felzGolpzZ6NDLac8bOY61i1+xg268yqCeg2F6QhxUrjukuDJ38xr/gMBC9ApHY8+5Vw
56Q/JMQasRe6MV3eNQe+oUqRo9cjRQdZQyVXph9F+UAbumX2Sr+yy93M0acZ/WWzEDqbs1eC5wLl
H4hnMV2mokTW0DEdhHmDaum+dSiwoBAwX1JdntStbdF/pAOZm73X60Ns3P4PHKO1QE2wccWuqb4V
iR1oK3NLVreSzDc0RTL0p/f02VNQi0uENmrTnyNOOa2tG3okegns5B897m4KjVVi64PkTJkS7xNd
NvGg2dmSuD3la4biolA//PjuoQ/JGy6hzgZiDEUaRZldDqitTmzaAaq1XuHd+PP4VAZjCo7p8cnz
KVbmMCH0JxZqLvQRMhplGMQRMUaA1wx2LKSlVCokdDP4wK9ZmwuejXN0bJM2tvPSndxGvYCCFp6E
EwCHdpiRdgxXAHMDhoLLjMVgqfqn5mnrJebOjeAF7wDcVkfYa1PPghvb6brxeuCsMBAWeOZFPML6
MzUePqS7s/qwb+i5GbuQqVmX7IEOOFI5gVugqCAy9YygxD2CAY+SQbW9TAm3JVLxXw1ad3O42nMs
joEHPkVkaSj0qOXrPjFFAB/XTh8uaUflEAVBJUwJBHwgwy9CtDxbWvIqH58J7/e1p2niZ1o4uV52
FARAFuCDyJIJvdeyz1G2UjyorTou5rhK6sFLk2no+ntx++8Zp3vM1FJPpQfxnvSbCnnk0E2hfB+6
rp6ALiIo39jSU3/2Mv2r5gJX9fzKzsuBf9cQWdaXR4zI/WjB9sGMlIwAZE9jVxK55FgiqQXVJteO
kFz7xo52oTbrs2/DhTBg7uLNPjT91WYNA0mJ/Sg3+NvPtuNGXmupazCNW3V94aXLd2I7S1Hf0Mdj
sZotUdkT7j7wVXFlDqDyKkLmtkN951TV0Z69mS0ZXPuUCyiCWJC0UhJ3us0AMMCwhDjJZ3L5AZj5
W85gnktxTJsZwWvnRLddY9eU1wlVLveQFB3EuvmhZiyvBUyp1El6XzDx2dGyj8T9IL7FJ/1tPmBb
vdlODB/IkI7OmVuWsRzeu9J72pzfWDkN/HMpz/ITn9lOmrLRlUcvoH/CKrjIk33tPrcLsjc04eDM
/iGNlpAzKd8lPvYkat8/uzsuP3EscGDSNJCzgesC78eHXuO1CbOSFKMpGcf1PozPSVcZmd1LCS/0
3vdMPn2VQ0tCa8lB23dU1dqRba5Rc6dXdsQIwoHIWtZbmEfnenhzkO0pjNH5CMSbr5cXPIBBx4kZ
4CbrrE3ALs1S2oc955bvB9z6CaK7nBgvtzq2x+u5XENMue9VnIWD69FPx+TBRBFxqWTOfv/J2t+b
Hanx0UWtlkJiqhtu8+v3hkaY3HJdXFegkrJmAPEy8bn3OQ43cZhEADVDwkJhvCGZYyYXi7b2ztfr
P5lxOPCjmYBj7TCCWfFo27nwQufwE0P4/jHdiBcLYNrM60CMVakFDBC1+bvAVG9BO3vT1zHoxCfW
hyxwV0Gdr4y1t4FXHyP+SpytrFl3i1kdbrov3i1t2UDFoYCz6XOZ9NY+u5hwhuH+O76bXQE6IYxP
SoECG1WxbL9PdyYC0340vyGLKQaVh3F0PL3cdCtUpk6SP2ovk4gsceQ9Y5A7TVxllAkZZmvXIZ85
SzDH7bcvz7P4UCiib7qmtPSgm5xjqomSetviQmfRVgPd9+tfCFwdvX8fA0b/PTTiXsEG/XU2wUL+
J+gSkoEyV4UNHJbfkFlQesjagsvX/qqf8462/f2rOEg/co8te9BUDB6QAsvBznsXo9He0YeWTIVv
ZukHjJuY4UmiwVIaOjjzQDr/4eGU8vU5x9XrMU58jAj45HmUbgHJBXqA0jSd/i9TlTC8iGqXm7tp
TwGMvoc7T8rSB5DaPWdEyBkbbuh9crUJ75bHIzRE/m4eAorYCZjIcqjq+HBqxGMIoLgodKiYZwHE
IymcR2OrMiezRMBw58EKb5NYouXbDSqYlbHgH48MV/vzFvIFKs7xD1Ka8Xwlu3Qasf1x9l4XvIaw
3RT5KNtokJuuqBRW/5jmG70puedQe3sykTaJh8e5/q0VuUzSqwGiE2ABmPe+3+gOyAJPiUToYjrv
T8a2rrTw7IBJgILwCaA1FbCor32fe9ARE/BCiHG5EaS8yiHUdxZmlDnvsE0156rjdJ2LmKVRLhVv
D8i1pt41Xlo4YdJa5klzF4ppIGRbGI5tyG+2Vc1/ivTudgrefqvj08cVJ2AfZWimgoMJ5x0hs7pE
LBmEllauOA1y96c31S/3QBf4HPgIbiAP7RNggUtETop1+2vZl7IoE+ElEJa6bs0q5t+HmwZXJuMz
8GGRfRlbxnp6jZZIhCLzo7nKLyOy9GO00/Usku27jS9QqdTbcVm8NXsP3UfkEi3+6B97X7yUI901
Uq1bGMz0aGYfibR+vHwciZtKCrcID+HMysDHbeW4YXrbvQB4/ilC3quAJ42yhgWRqc8p9BiwitmX
ZGtU8+Jt+3i2EA+StyxWv4Aeta2efsTnsvUMKw0maL11OgCrf2pwXsSTSLJY7W9Qj7qQBpr36Sxs
EWQ93s/bl5jSX3qwJiNAFKnKjgEbQTJZ7WPV4J/u8jWNynq8Et9yGIwJkydfFkzCiWJB+mGEa5nT
ydp+kLjUIlzQzxD+jpMzBwqTtpblaihx/iVd7OyrTEKnJcL1qUupubyJW3p0JuAaoWQot7DJbqwz
rsZDCO8a0uoFbDL7By/2K3ZmcR040fy9oSOTb5EmSKHx7a1FQ2fsoB1T3mgey+plK5kjS7TiTPZE
aBjypPCUzIGgzzXl2CgYVOzAcoHgkRcD6MFjEjXsNeVkHpO2fF1DCFxMgEPVZ/EzmA988bqWapD/
1Ig83tmY3atFvfY7+V2zh6bEnQ8TWSIFVu4hl8M7wl1z5sPdnPs0o4wpqHV58ojn7ZDfQsa9e7se
QFOpwMxQHu1nMEwTcR2FbfD2gw+wabUb7yPS3MuUc2X+zJfvauxaZiFWbNz0TYxpFj2+C6v31586
QTLDD/lPb3PCLQ1CqvaVr2PoxyxNgoVQ6SRxS9QD8gm0cnG4IwFT8BWBA0xd+l3mUmN95nIHTkXs
Oxy1MZ42T26Ph7WG9NOcoymmtQNqFhEcc/UIaF2bkYgTQkBu0S5WUhSWqNIG3sn8XCMFYmGYGRfL
Vqi0JDPyLe80BgrCeHU4o9SEqCtkBR7unZc/f2b2VxyhhzArHaU71Di7bBoR7b2RTtv4zobGxFM8
CK8Sg3SMtDNJ20dVeAdoC1SCDU3izVgYSGeCG1sZxUypZ/gQpvOaA1rsMdGT8YHdEggYq57dO2Sh
qxOVAiorWieQZFPHxBNIizvFyX0V0RifOavcvjN7GHr9LTdWObf1AQ4JzPaf9q/i1CmOzlBPXc6z
D+HCkABgK1aIdcI79tzuXpvaX9qPI/iEQ08bQbirw38/+8pueIc/njwrm9pQQ52rZ3w5XoEWfAXJ
hkqN7ok0RNeqeCJ4fkoVn3EB1ggkCB4Spca94mWVWTdDlyve09IQXEh+R8GX4iPN65i5im5j2qKY
TsAQHiAYgvHgSU12GmtQ95N1zBuRSrRzD3TOOJowzLd5Z3tATR05WgCaZHWyD4mBGdrSanKizFjq
nTdKwX6JJWP8AVfqUXPlc0rZQOcRvdFQ328WoPWP0Gg+iup9APa/g38g8RZVJLFluzK1J5rDj0gn
EGW5fvdRNxs0rEPQoYEDtTTKnFX2w8lTskN8oQMJ0J9LZt5U/5lTwzRtvRoP+Sssy1KuxZgsXJoi
439ZTVM/zgcP4aPufPWwCf6N/kBtsjbKaecV9d7Zub07CXdqYSp4P60mP6JWx61SjEYwpSxREe8N
B14VUNT8VVyMteB3B75QdJv8QF1ViMdlnCjXCMQAbC6mR3/LMKgNEQoFJZBkCCg6872eGTINn7pn
0OdTBTCqS15jnLKqjwxrmWF5A01GJyXuMLvO3crd0u4NbYiwwlIDj2khFX5qX2TzGdGFi9RGtZYu
yxZj/B+wRv6DzqB+sDN4Tq2XO7GbLOTujcXQL6RKJOT++CpQ0UO1eqbWY/YAQdrPnjBc3oKhPL5A
DA33lqBFPQ14Ch1FDG26eLwE1Ei1zzKRR2665wpsNexugdr4YGsyUCPXjgeL3vIe9de4rGgwvI4N
npf13kihIJXSuGUp5kllRZQZj7KVL6+pk0g5xr+Ea02JlG+GiJb9uWFd+xTjQZL0Fj0nihS9osbL
gw9XLCDBFdbnfO/yFtwBL1c+oAIa2kVnOCyE7DNCYfQDmv/45WyFNeEpaTQfroN6SeDsMpJcybza
RnftqiyDGQj7M86uGcVdWBhgw6L5hmh9pOnqdQeh2OK4SU1jgQdpPCl7GqWA4Fz8+xLu0sG1oUcG
d57y+dpaMRYhY4fokj5PphwhaskP40DJ/wsQ/hSmX4p/3ORetqoDT+PFlAV9g6pCaL5Ps0efzHFO
qMc6fPfht8xDZ5AH5aKPj4KgYLGYX0n9cYsr2Oc8F8ySmx4WXXlQ00ZcQOFFxpLsH9TYagV+DShC
VhJklzSX0n71q0DhVp8FOMT/78a3c0VrSYLRIYoGeS0vkpw0ljGXFNxkAQm3c83MIt6VbdQG/V7q
kRwEsKAaYs1XHP1vZBY55AXMmA72Md3EAdK/4FCs6MK9+F83wMfXJKQNVMdFJGRLRfO93pyMZBzD
SeDts88HpGXAvIaQ618SbgNEAUF/lSmyB68+6ThhrYqudAx47pPTsk1Itvit2mZfU/jT9P663wi4
eIhC8dmjM16z0HeMg1+6GrLlE1HzrBoipYQmqIT6T8p3ZY//mnzAujHQP7rKXEchMxDowDKlamD5
2m2OB87IYCPj4VFe7OUp/W908GKdr6x2hXxGCNjoFhcxrckrZ5V1BnytdjsS2kiOWZ5YMvwd9lAO
8egd/3LOVa271mVDMN+U2/ZZG2xUcFPsNVkhp1j26xwCoHk9Smpp9csFvJUisXFuN7LJPZHcrbog
0SQI+bfD4fZw6PIRT3cGWBWzCEWTVlzPScacG8D9PK+SW1PGA3FCwRXcJld1vp3VGUgTn/fCoctN
8qoCSOXEKkYBlon3BGMDN9ETuU5MTjU7pqz9roiMhOPUZVxVoWrEVJui5iwxxtP2nEqBv5BpBIlj
ZrnAH+MLstaQmY/2GnPP14klbUCQE3KblLrFl/jmVzXIYIyKWusmUgfG9q85e9shBVVkWZFtnkTs
RAuqoXAlEFKgkE0sdGgEx52WDU+LMMX4kzGuVTqwjjrgJ/HzJxC8JHTvkeIV3fl3XqCwW/lw0HTJ
9aTxPGJqdK17b7+qWw5iu4NJJvUOD0XgI00pt5GB4w/b3IMR53o3jbm5/kIc0lYoVaMu6C4a6XKM
bj6Hj6AaVHnBdd/DW4Bz4wgPzW4HDLbLULaRIqDNAkb2qUcZA+GOw1fS8EfGLTlC5wBjNylqYurQ
ZNMYgfGWhL3Te7DKanNAyj4muze7XcCOx8CB3c23B3C8zV2QJyK4JorAsshzNCCbIRvNWRSX5asQ
3fhUJNlEC2srIUcGqIOfTB1WQo91a0HH8LK66Gv+iLkSM5gCVRpxCqSdxg7oy/z4cviXTbPWxFEB
QXJ/0hf6s0C/YhYHyHyX6vsUJy5PR7mQ4hWX+0d931pfUbEWKnKHakgyvjYfkcVBfYOeA6jIzFqT
7xH86urvIksJ8Nf0F+lQgreY0HUSAsxrpRhbpOjhmvHVZg8bFM4FTNs1pk3nTXrK4ybVq+myKtE6
jzWmJV91QnM/o//YY4xh+T6W/Xc8QPFdHlgTuO3MHHAFhibyIe2w4HtOfWVkZdXwWRtfYuSxJB27
bdowsarcKmEbaWMBX0xKycFvdLH9jDyJW83cqGTG4siZZf/j+v3t0dj1+2q0w8m57l8rHZqKb7+L
EaMcFeblnVHWPelQP3yri9B3TwmJrdawfyQfzJ5p0H2LgNDxwfABH8JHJDjiOtuEy3s2aoPPWjvo
2QarMcTQKLy7ierB55B0K0LmwscZA8ICWaESkWUx4t4mOP6ZU4BlxhBcRiPvcHIo69Lu6xJjtc3g
Kk4V00qZiLybaIKFty3LAUbCPaL05nsNAsmXs/RIEJ+YjRvpGc/ryh0qpoLQX6pddJF3FZ/vgFo+
6UkpTGp6/GcpeEmyVOoEliJeSSzSe+hg/N0gl6Cy4nVxflR/SmHRIWB/dzhspGG414+gThwk/rBv
WqHBiUCP1oR27VNk5ECzvn5/YJizrWifngkeE01OgcZR0xleV24W5hq1J/zWnb/NEVxpw+cPHLbN
qeM0VF479pVTi2DdcU6eRebQLlwD0ZjQet129vm26FJlc4lgE0iDDOnpNbXot12zK7SuJAYhAkQY
i9QMyjHsLbMM6LNwq7opvy+cP/EUjDYLAhOQ8CYhDOkq+2vzn4vtBPJsWG27M3b0c2p9+AtnvupE
xOQQX/OtD6mZffxPEbcVI1TO6eUEIXTR28ttMRbayDDJP1Oi3OPY7JpR6FQeGBLb4uHvE7C+KCDa
7pm24u7d3p5P/yynehvWYRHnTK+CM7ao3gwAHy2Isqdl//M+4J2g9HD78XFfMl+9sLAkYu+Jw8rG
p61fBOOCNIQeni9W3Zq7AigkW1aTVgg/r5qThXxA5AiwdwPsfpg16+32SNC4OSEX6VOkr5bwfJnL
vFC7ep8K5coIjQ/pno0V48V1AEP9zNodn1iYT8xF4Je9lwq8xRZHPGKqthXpwxxJcfJ/XPXtzF2u
K3EFxAaoMn3ef9zc4wvhwC2bxq4rHRX8yPebAwh7ubaxLc5mmCFBPZ8aVf1j08Aa0U6+ecJBJGNf
Y/TafQgHFvmqGQfW+FNeeD71ASYOM/kc7SrVReAF2OafAEMSLoouwVyvqbF+MRuy2FSNi3hPJn8p
r8KmvXv4kZOPg3b6WKyttCs/pEOjfwpm1JNgAmC6fqrDIq9EPjDCjYgpXxNyY+f2xCa4fcmDTsr8
AiiJQ0DhKFXX82NqjjiWI0ZCCKxUvg34wVAiFA91XemkIrfiYcuAZ3a0yl2moFE9ofMa2dbiSGDK
T9YiUGFB2/HnSNA2FA+gOvCFmLfMDz9dxPIUSNif7Q14AguEWyllAtw2k1olDqUL220BgRgze9Sw
jhzOHaoH6ARizvXyKHyu3cg3o4OL3Cd8EacKFJRPU5a1iQnw3NmQUYTFhPl7s2Th84KQzwp6uqfJ
Op6Z9NrUHB6V5OuMdTtpBU663xE1HTT/HBH/RrH/hrpbJm47vSgW8Jf/leRljXDMOQ0Q8UwN/6Dr
kthuQWlT6IeF238YuUfXVc7+o3G9dC3aQrKMbqdX/QnXYzAxtgZN9qwSebX6YPzdoiY18pFDhf/Y
W3AnRIoVx54m/x+6bVBLccGDOfLA6sKj/juS67B5gYYG4gl7VSQu1J87UGbEWbQaFoOgAbR5thBP
IXS2dawmumWmB3pIXb+CKlPuoFTVJ9VXpOWZ3tKlZ1mzt+lIU5dWj3Ex2aRYg5IF4vOegkKkDl7l
wcoJ2r+ycQ+1esuqpjxGd4eKRLVCgHpx2Fp1OdstghWT/Y953cNn3tv7HeOucc3iWZCAWr9Yj+3r
a+ZnLrddcplRrSeC2fEYv8QzFX+Y96h9vXvJ80uKFz+mC9/d6CqXuNUoRgqcLeuskUycb1c08rIx
HsEkU1N1A/LKc3OxKWm1K+15PiYipTQYWFF6JFKcCg2Y6jx4uWEpwLkeLDODmYZJuwNh1+RwV1AT
+1mUXczJg5R7HsXOC174Ye7XpJaywP6zbbkrnHG22WF1WLLQsHvTWmVIjE07Xp+4TnlufB0Icgf+
AHW2CzeZzBOLhcCaftsZYY9Xfyu2Jz0UP3HfczRcjDRdV/b/bP+EEWXNxeBrNX0iwsoaAbcdrljy
WKw4Ppy5+3nQigTo+yIa7jgU1p7Kmzq57C/aWvcAdrYWvcSSU5caXUlsfb2fsZiHJE4I50c62K4o
umDJxM6hLx5oo5od37DWYafKzOTEktwu3t57bMHGDdqfeV3ZSowZEZp1wHYMUBLRcMjMER5NB1CU
ZVF4UNbTXq5nf/LxcVNrYQXUt1pkX9SvzknMleCm7LfeSqJaWs6e9IaWgDJDcCeHa/xGUENlLQcX
tRgfhy94uzgwSaLW6kLbdzasedMk1L1HUv9Zngep5iP5lsNtzCZEEZdt4kBscMvkfNMipvx3tGK1
Oqg0UXas3MP3InWJCmXUUu3jxJ710gcxA1EyLErau8ldGWV7rSLwSTMA4Jhj6WMGlQytXRZ3t6GE
3sAJGFxBWL++3mOtHG5vNlUaUUX/GBlBvsTDa32vECIHHm/DKWggNIQxjZspTDoXjpDTrDZdYnsv
ZD7n4lWiv3lNDZO6jb3xD6bGh1ulh66/Zgc6SLPNqNPl2pqQnwPxH1nFfdasl7DDDIuOnp5+pdpM
C+8AqvY66fNeAQoRapu2uRl6x3EaVzIhLgZ5LOgEJFIJyOspQ1BYePdmfDG3CkKSLBwSb4EmADrp
p/LNDUtzSvypPO508UgXCB6phDQZQb8RyA0gj3fv+39sSp4lWKCaVOBe91Wim8EGCbpx4bmisaDV
zSkxGcbVKGCrxHfOSf5KMolCeLsPjjWcgWXFTXGSF2jhomKmPyIrPXAXHGq6IhR6jfGXLyt3y0M1
JCWY/9Ko22ucd89V+/v+Xtiv42dL1zH3jRPDNCPekK80OP7wQ4qoSM9NGEJP3k/zUjwn2PEGUfKS
FWzFc3DKQCAzGBajDqkGQMTiZ9HcShujpAklUvpjJWDy5qaBHGLhY6BohnX/JCcZ4bCHbVzv9my0
WhV51GDKC75Ydil5F74uSJsnbtOZ36RH8kkXLjzmBKEtkehuql19YiWhv8G7JJkmJ/HTUWROjW8m
yAY7d5kJ/vJvGJweBiMVxcAaIszgCofXAVuU+dwhu0/GM+PGEuwo5s/ga47pfNgcZC0xBrUZyHmn
qjZPTPS6J7ZwRSZN4rSNRa53bynzX5VVXQc5zu4GrGrlS3Hm7ZIdTE/G06vr2muuzp0AJCdQZdc/
aTTkFAeoogJSmJRg2+vEsXBzttL5oEqQ7lBt2SfP4LpUGZTgrW4VWzrlqr35TDZBekL3tR0WsX5h
f5nH/0q6vsVk8/eoQJR3xyd5J6vOv0ClfYw1Z6Ro7q4HSgpCCVnnFFZEuJzrCrixJmanZoxjewma
5zInuyn4HYrNgM0eTX0PqZ69350bmtj3wu6Xibie8ssgJ1Fw7HM9stXElYgBLiZkHafzPFVT854B
5ibKTtvRp203s5Z7qWz/4NbtzBRcD62TEPz3lxvstYqPxiTk8nUa1t7i1TrXt+5d8jz6aR23wDbU
nXXXxl8ugR0enem4pUngNo7EME5nUa+XwY5dDnsB1xFXDF8AyeKX2P77E5a88FpMQH5tkioXsUHX
m8FT7393x2Y//TxhFodqH4/15MkEwXCZmWEVLP3gc99rWgOiVBs/g5P4uPdJEoTvUxyEkLl/ZEKl
05BroOTQ0xjJ8cMez/g5X7Bc7FdBgLdjGeNA65A8W3zkQrOpNDoSOlRd4+psbjWXMcU8yGj7UY1e
sKcYRZLk9U3ie8MitE5i23wf50jbrVeaPzq91SwkoOr4OWKdZSkf0WRBX7NhqMhxcmZmFhCg5uI1
+seZbhAXTwhECn4rafONMXH/pMrV/B13/Y2D07XZQr52UoAmvqmsQoD1MuC423Fuf9D4gx3k1m7G
K98WaFE0ZPZ77+cia4L0GuZBAYecR8vHS9i1i1jD5bQsZtR0a1q4rGW3+glXytwlqm/u/uUVgfGE
0Jhu7V5r3AilCTaH18gN95G9R9FiB+Cc9B+K+G6jozj3s1byYpE3fR02vi9UDlD7W0yjVuPmhoGt
OXHWrrVQIPqOQHte7WNBqH3GU1EZKBGVk0SwoRRYluGgMxhno09Wtj7/Hc2PMWoSpM5SQIjZV1gj
H/mc5H9BG/4hoLboJhTDjUcQKi/rjXsyXvk028g1SSItHkFqeHCUk+D1Ro8PXC3fufdZXWAjQy2x
0J4emNw7BxwnZmyyx7yOt7uaAN3Khe0lCay+l8uW6K5vtBRidq9FrJnGqI/VVRS8oSJ/RDt+wrpX
xN7ih6PofCnzP78fK4JqnZCvrzMHG6cvWhMlLje3bdnltQXnx4W9bg8zl7aQGjPxOja355nnj3Tg
co6BJZ2nxjnGQWvhelwAPQ8eymXYAypG0076ZkLtD/3ApIUDOzwdYApjKp5p6yaQQqZcsigY5Y54
uLXxZkOTvxop9EbFjHjvxfFCfdGHM1XT0RjAsyywU9GHhIYMt+PcvmZcqYV5j83qh9j6erCi7xQH
MgWZasU4WF5NvK+OAq/sN6aYQlv1UQTfZrdR22S+1inc9jnn4z3M4lwGG6+PmDU3cXzdPSUZgUzY
vGl1/eUnsBMzox4cAETI8jrGVyQGE/Iww3R2eGddqWLpRTCN0TLzc75nDvwOnHLE6GdDlGLqAndq
3PUd4xyF9AbJSuNwJ4UFiJsIJz5gbiKKyGFq2iaOJGjzTEybwXpsk1HLiGQW3uvUov6bp+rO/Eya
/n5dAxeJrkI6221ZiXGfsjVN/Dnu9cBIEZo/qkOPlfQzzeMzH7INs+JnNlL4q1KyYXlir8loBybZ
TCqb9GQSkVOk9x8xAgBqFVzCunBRSFsY+Tgjw7SOL3+qlcwS2mwd8QJiWggg4XpOvgx+BGYlOJC2
XaVwcB/4KKZy3FIUEtxiwPLTCW3Slz4W7mpcz0sL/teRuLFbC4waUN8VbTtLGgR018EA/Guu5v6t
2is5gpkYTorAz46opi6V7UXnDLc4bpwKVstl1Utbq8Rldv/nU4Mr6waT7cGu+EZ0kFKEmPVeDQ0V
SwcC1HY3O7jIUlc9z88cBh86qhDXtGevLmNBkI/Kk/ocj/itHs1W2DbxIBYZyVG3shKZnF9jMIu7
Pkn4y3L+OYEi+W3dNyDaK9V1ZZ+bfXqImX47N3ts3rdRn6x6WKudgf56hqHquGky+i32+TuCnLWz
P9XAd6yYqW+swQl3QjeJ9RfJVBckhcF+mbModfWY/GLqY5n9XUHIjmWnOhh+0Q6SHxOJ6gGg/bmY
2hgK/Dpc11AbgiHDxLHtOZz4AwluLWiRQRdRAc47l1mRQC6Ug2a5ds8D91RkRmRcCEedhqVTy5xb
D/M6C9DvkS2HMSjWRGYJTOlIIrXzkSsqn+yhwsqhJGccAdwM8GecwTo4HYKUlWnHRAjKubrkqh/R
lfm/m6sqlHacb98MbP+JF558PjCry1ecpOOt3Bm5Do7fvDFH+Oie4qYDhkIl3VtC7mNVC+YqqN8n
l9ziKb5fxHH5i5Jy48GOk3D6Wy0ggLkkWeGWLoC/zt9zKO9Cx/hHdw1vtOK6J8yPsS82a2H9Fgkt
r3yExgwaZpfwt+7sLtx/AT1h6kOd+qrJLTQjiD++1KR/pB26F+JH96l/8DaExu0RPXf19KgxLewA
jU1vNnTrv4RTQILzOXfNN+MQ7abdzOX6PH1AwV9J4gpuNHDtqxctN7LFW662POispkguv4zDSMxa
+09YqauJfxl4nujRP4NduflB4Yr5btg5Iqxr6VbMmSH6nG3UHaIweOBJRNGA1av63vYy2EVDxN4b
PqfSJ+ChTC8kV/ucXXd1pktSj5P8fqkbbZCWbDvyXiLe3R+OEaK5MSyBSIp1teaVrVbXGj2+mJhn
Phscwj8YmnE0LBsAJyrJoQqM/J5S97z2uMEeoDK8kvaTfigdq06YYxSskDGJ8KaU5ylJ2Fjp5s6l
ZjelFGnJXswq2NV9C3cy1+m0Yaql0yVnoJmeV+39g+GT86T0rwRa4ICSpm0SZ7UGX0DvROhDXm95
8Rxhc6pnTjI5eC+fwx7Eu7jC6s8MEUYHZrDRSKqXRRm+eKp3Ytyb330akghoxKKiwM8GVfpf1/Ub
iq5wmJxahBLEH2RfoTkW1cvkaBC3RF/0ykBYrnpts+WfP834ODEmMCRUCrIMbyqeWFacexfL6GGg
84CuRUSwdV4baNDTI/+zOP3UZYrkLbq3BlVFZDmlZjmlx9ROs5TcrpTcErqN/8nxa9JG9fcfUAvR
bcmPdnYilef0ja2EfL3QZJLjzd43Cvk4i4Sq4qUx4t7Z8fB+khVtGcKNoD3BJJ48EQl0PmbHkP1x
Sm+rMYJTOGGmKb4XaONHy7KV6jk1cKkHLEO7HUiiArCz+XLgMrkjd5JEu/EdcmxVlrcevettEFqk
xtxa+8NmoBfOB0THYyyxrijyTXCJdkQZ2TkMZCXuNQGMepdqenzp0aiJvHYnvBaQk8XUBrnel8Gv
OKWDr3lADIT3yBfb6PPBdEqr1tVKyxZNtD1gOUsdPQ2YvDpQVXx2Pwf/AVNXhamyqQ8ijXedYMtI
mthOJQvJEHbxfFDS23934+iRSmleSjYGDlLoh/JsRvn1hiA1vp2M3Z/BJr8eK0uQlkBlpdxGpMa9
vS9TFM/h0dcbAU49YAqmPK/7B42n1sqNs2YYTi1Z49sSU5NYF8+1qdpzdEjutsLNWYp0GXXGLw5i
NWlnd6KQBmDa4NoBcjzni8Y7qzkDH3OjKiBHwZYni4IYMjz0XS0HT2NaMHyQJoTm+kcy8vPz9lS3
cqXUWPEAVtdW0zVdMYScjDI4dYI80Sc6nixC9oBEOUnmyHEiIa0b/89yd+JzltxSKkwXoI4v6238
Y4260HGOlNyhPpUCEI0tEe+YCTVhSzcXYgKFHQXWv+9Fkh4NtgN/PoAVzKFU8ZO3HPdAQXIVVDO1
3GtZrck/U0NpoagJ8MGJfQFF/r1KFnBUSs6YIx4BTHsS1FlfITnRkvkMUiPeogvz7zHPQBlYhax+
zLwebGWnJ5OVsT+5OY7zdoCvUdBa6GrQ9To9ZJmqGM7K94A8c4OwQXnoccCkDLpZj/DkFT/B4pFy
cyhCnleSt9XrIBMdiTLYChmM5z0P1P1/0VgkJzx9CtF4XCDIWaSWHaS86pzR0wQTV9xYEqk2giX0
hRqjq07T6gJhh2c1cZvWb3sXS1Ehp/pipi27Vs0QZPSKK+E88SD5/jAhvWYXRRJrqU5AUPi69Cfx
0aUUBuOWEnXn9oEQNgQcZz9HhGDGULg2g66u4Bi34Em/TGMksysMvDQg+iz+gebzEyuut9OyUKG9
1Rw7olJx/Vv3+wkd8EOi5B9Ith++9JuER3sP6sgmsMEqPMhwfUKRs0wcf8pKvYZRNVMqezurYZhD
yegfWXimSQL/dVxKXeimUsV6NEr3M4QeV8CbBCHnPVODRzyj/C2JYrwfpD6c0WMXDHjCUN4wz6d7
ZY6/9C7CG7qVYLCWX1pQ99d3pSYK8bkgVlTNFYuMfMQnZoFF4E+tp4M8pNDIcyS3/2fG7HAHQzmo
i/7Zwtuw0jjhkXnH0Uj0EF90X7HBAe3RjPernUdVp5bRvAakTJUaWd7/QrfIaxdGpqtX/VcmczCP
IZKzB0VA5LHnl8k3qGkxQxLas2zG5NzGOV8BipTCodlS8QZ3ty0TARKVYEljvZ5yTh22Qn0toIxO
L/wysX2GHD5v9TckKkF5L53B7Afv+mGR8Sc/YXqrbivraB2nFC32aVbN8I89xQwKEtpBOdgU5eRZ
AQWG7/QKuPdKzp+WQMvQ+yQe0I48tRZUnXvjElnGlB0n4/wDUJIRNRyKCT7An1joACjlAidSBIsK
bJoMYHSn9NdcnUcBBTtHQr64XxMtHeW1SBilU61qwSKkxJ26hWFbXe2srDTiiwJHntw1wMmoY9YM
5Erj4/+WfxDufSinSahwIJa05Bz/3fJqBrQI1eVVaNsnVJLjBUYtBXSpFS7QhbiKQFyZ7pRHCuKY
SgbAnlPzQY8yu28sAdnhiXFEBrV7zrBZgIpDwpxK165QvF3GMMc22Cg9Lm/LuqKVkhWGHD3LRAbl
/FnXBZCR1yi1a/e+3iXj1ou80LzBy283pgz1K5uXh85VEOuZB2+KUXUPMkPZa0YvaSC9Zm/YHxic
tW0EvIGOzvju4ZfCFLa/7W/RTuQtzQeBpGqBLyCF+56nGY0BY3Y3ClWt/y0NwC6A0/nmodLTvYEF
WtCkv8DUWYDfvCMRaKiPg/OvP7dzVPn9UvMWj2gH+HD+J2/rVIobTCQ53fNEkRUckzhq0AT4VQoW
oGbta5A1dvdECOoHdRY0XqApxsZIKIulqIOLdQ4u1DBokyDHImf3a5jycsVPqssCUTQvBcmhR1lv
NXsnbonFGj5P38WHfU4zgyYEYilxWXSCM1yiExugQbr6qxxcszv+MIgWS4sbaPBmnUpEZOZjQR81
c5SYl56L5oIjGjYgVzglzV4T/jyzic4jiuEQO/a3NKJ9gyUeCgZy/SCMzdgHmXjSSF3pPJR9za85
8zfROVPBwzM6lA3qYyQTSv0euKHc7A8ct3+pC2PAOapEYZAhRspz37udweX4Vkc/dW9+XFolOGiS
BUd0yNP/iArYMjapUNFIk584IAff9r5X8muKF+35S7SSJgBd6S7ws4+FbWJNKC3ikzFkkbpbXcwy
pl+vUUXJoW9IrHaZxntKVVjUwfoLvtRstY5VF9vP3M5bPLzVZumT9fn201E6oBKMQrNXvK459XD4
yFLZk//GxRPwWiFDiu2Be+njTezfCHaNO450bkh4n//O8Sl/M/iInjXUMAffq98qSaWDyQOsolfI
9N34iy//m1EDDEzn3LovLwFLS8p6Q7Zf+IjbR8ABSGuagn40llGQQOavUgYc1uRJzVNJnuFRLHcC
WqhKcGgKxLh2wWQQ6oASHhEvBzHj4Vy4Le2su3ZIPRWKOHFYVcpNJTuZu4qq9UI4FAt+fxHAtils
aLsjERkRzPpMXLSkalZ459UcjgsGodZGLb1ToI5NThbthZYljH3I3XYB04/8Y48d2m96OsZD1w8n
AZtl0wY5hIlVonLEuey0uuM8zFSaisW66rRSjnjFFxlujSd70M9WT/+D+VVPbWTg2OshqfVormVi
Gt3M88cjtdajdR8uAkkN8Mk+kGM47jNCQy0dOmF/c0NQe6D6rPnWKWjLzn+6SIPzrXIh8N1gR4Kb
32hNn3qJjtRdACBYzxlAu/iabH3kF17b9AtpE4S87OlXNN3oD3ZEN7uRHrZDAX7nPjbgSRVn6uq2
KLmqmYhMmfnyKgWDqzyipeRchEx5DNKZnp99ZWPwjTJsihg+T8eXB13RGdrcRpEmeYYoH5uBToor
ZB84Q4AaHwzZ5SEIp1ju9TRQMrOU6NMIAgRikkJAOQ7lDz3WvMeasutqvYZjKv3oiPUu5rFB9LFD
wh13qRUpU1eggsNdfvi3ZLpwQEb142hHmYqUbZ5PmNz0FeKHd1W4kxhDwxb6JNusmdQTsb6je3Eu
3k6wXZAbnoH8Dbkm2jq/wWNCWsHBAV94g3g6S3/BvrTqnd1KInr4BoA7U2b0xDqNrUgbeks7p616
T4xMs8fiy8/uHPC9PLrcki57I/oygu6ysOs1h/x4cAWKE/ylouzJ9cUG8opSdPfGAg6cfoetgvBB
krFLvEoC0Px0cw+0Z6u5GG41vTHqggAx0S2lwQ7SB4tu/BmfhWwQveNx3R+L4fpAKDsmWCRXz8ye
g5YzIL6jz3O9R5lj8wV6NjKtUDV0j726K0R6SuelcwnbVuwjYH9eDqGB6bKKYD9F48SQ+Kqvihzw
bpoefCtBx8xJiK7245hqZff9a5C+aNPQc4F1F83IvAuwVDMO71O01RD6FkrNWVdY9nnxqJE0ARdo
Be0wIkzJGX4oOocz2z8kEIgtIb39csLjOe6QTxtxs8fTZK3crqL4rvr9UtcwcXt54y59zlnTXGEC
uZooocg4HlDrfPp4txzx5hLJMkts/fe4ZlI02sfGzrymcPWG8tWFkvn5zLPgD0+qF2thV7VL/m2d
vfnmD5VWIkya1QcTxumwi/KImISCEpHLSSIfvMDt7tWpKoN8b2lcOcIxD4H/yynMU1dM7dHyFRLR
kF/dlplPJ2qctpHnmvmWOh/pwk9hvXrLFmW4JhnZXpJLACBpZdXtXpNXkyP8TwWk+F2NFJjxLvOL
A5sUIjPrurE/En871EYBIiZ9Kl9Fwl6fKDWPNS9oI4Yvto8AUIfCvn/lQKqNYCgUt0ufORQ1XHrQ
H06P5+bPDNhXGY27YQaqE7I1irAKep2gkEScPIunHeT3SYaveHu1HV0qcjbonokIlp5PTxxCXDHF
47VdKeAle44u5bcvoGJ4YX2wy+HPOXCf2DP/oIDG2bUSYKFG2wpdJyNR6hh1sXtNflTAJK7vrRIK
L1cV/u0JAQ1dyzGjjcr0VP4R7ftGaPpjwsU8rrCW2r5o4rzz4lOvvNnm8tBzoPEj80AGh86ZFU60
jmzhGZwv7tzt4bBg6A/qYDO7/MihRheuvE5jtuhPRAzaYrIZqmF8TvVQKTNw/rMTNItxF0QTkAtj
Ce4m6w8SskDjTPqH89Nbn0aHzy+9kd1rgsiaS+rnvzQFlbBdVTpmDFAEdkE6WejZZgSeyBjA4nI0
WXt7zPjRKc9vpcyfaeY4kin49DoamFYqvToYxIXMT6FP6GF0GQ7v66hNypjaOmTmyleFGfn28yTj
E0cbWtcIMplurZOhGe9OWfaMBzAT0JbAh2UnALQalIzloJAdhHiXQ8Ar2BPFwXU0UMjpmCeBj+ky
9E/ODhzi/ZO2VLrI1zZn/RQAnQ37G8JARnjgr7EhQDZxUkI6sXK9u3pycsQX9qbcNkmNqeMtRu8o
fgQ3K8GceXDL4NW/wrHDVOnYHJVAppusY9TgkcTCS7MlaEXih6BJ5lqkSpuA9i1A1orqe7U/sNg0
5YOWtwCMQIoLMfcoT2oxABs/iIq5KS2JqnKiphRm5rzEKPVi1mkIzI+bcubWSrcXpURaHqMpkHFj
YW88itRVpFQrgXso3A1Wr6ipD/C1caWYzuRSsEzsWbfOkGPFb3K8CaXUZFhasb6rFecBBpJTp8hh
7eaNpU5FlTyRT/kPjXryVWfB6R0cpcVd5w0gYu6WnEiqTl7a4qUK2VG24adUOtizxN/29ojSKRwN
F/rEQ9FrnpXTNK3+0uj50Sm6svTzX47NpdYqTs2v8ytO9PDRnjIK7p1g+SF77a6q7ybto6FKrVUo
OKkWukYgbVt3RAuj/31ud0venTNWwvSGTI5nWdGaiHjE27AFtAbsap/Betlv4eMfMZPh56rtY0TG
nDY7DwIdUdk02DLxAZpfrfsiR1jLlyNv/gSPKd3s5tSADnO8ymtyc8pvFKsiJQFiP3ZUj6KUdUfI
G8D2TU2wtgHmO7o4SpToxVHUJ4wNJiRIygHuF9Dd2P6pNKdBWhEFvWnc3rnYfC4Kq32fuHhkhopl
uyz2xwm8B0CSJljKBMLECy4Dv+vrzEy2gGnoQcNw1++Qgr+zqhSJzFP5PbvdStNlrO0bkq4A9OXp
C8riY8msCXal+JTt2shFoq2465RKHc1TqRBS96odfpIlox7Lu9vH7lMjBOBBLjVm2SVz8N9H33cs
UavHIK+zpfhJeCRCXEKsRnpp97c71VhT0yx2KKwXpGQJVzO5yhEw2P7Km/HZg0+jndlf2ilv2dgo
aodSAc4PzrSoLxBr/upyUwD3fcKnb8d7pOi93o3+7qkGuwGWml+TGKMgpqJLN6uV2D8OU384pbif
ISmv4xF8smuIV2qG9+OqnTRhV7wlsd23NDSRZkZzR5qelQ7LUCWcTIecjbQYEagZX2qaMsLmkNLZ
azy/rLtN0nNjb0YURfEGt06uKaYaR4oIrvqzqVKGKO2rmi7TPhySKeJjqvG7nLMQ8z+p03ydAAlG
1l6JSda8hY+uPonVsmggEwlhllEOnkSlFetbFWTGvnNAjZugrd4fkYWMmDv61TgJqs37jEKGFsFx
EJOQspuoZ9bquiMQReQwIYa3QWB0Lve34RHacHKM1RCcogifx4gwHGmsEDlDi7CBNdf4GHE2qPqZ
tXmybTglVU3g60Jhrx1WYLqUmK6eRnuN9rOPw3tPaV89obxjA2DImfv8ctLShbutPhrUDsLhqHC4
f22INuqFmQSLvmn0T8fe1yx6ZOt9GUViwwpM4Vhe8qyfwHOJRKEZYkLwZ9TWkgADvjhiZFZII9s0
Yn4L0JUddrRoJM1RwHzt9IbnU4uTVE0WUnWMkggnXNx+WwpLR16dQiC9amWyxMwBO8XYta2FWJV2
yytVG/9qqs36Ea249x3f6FScnIsGT3ofRf26Q9vlbENfL9rM7SvI+zWMiSaDA3S15JxkTjgkaYtt
CdqneV7I8X2Zr9Zs4CcYWjWKtzixx3iKa+MHtCTWyPK7NUXW1ahotocU7Mm0UfgFp8O2Qrx9xDXL
v5WbcWa9StasCid11Ll1/jrL3y0aKh0UjLCbswX6OChv+PWjhlKnI30VG1RDrAmEobDtMG3iSCkx
aFw9EA7hEhk9JGsGdaImtpphtxOI5kYv8FiGDRPlxlrm42wHRKU65ySZ6h2/hTsH2sTsdRb7Dk4Q
zD+4eU9lCYLEYN+FE0lS5rdeU9UHbtn1L6GX9S1AhJfGPjpbz1zE/inVN6Uzh6rDVLCyfEOfCaEh
A90ve58Wq60Ua8xMS4KfSUT01JweZgIObIAB6+WpTaEysmi5l0vxLz7RTjLpUkjXR7bLI7Zyf9DP
fZd9mbqWQTcEqOmk0dSoBmUx0W5AYJSWiab8ROEYNygoYNHuLbXhpbdD3on18Zec4Gw8mUoI6Bxf
Rpo0Yk7OZSOSsYAJRQZM+Qrc7WG0SPDmMup6gjSae/aLmwKXY/h0zS+40Fcyl/BJ0aGMWnQBvisL
CfruG5RdBA2DBeR6royz434fw155YUU4jmvUgVLRlnv2UsYbZAfAtJQ89mUdf1coWcldUPFRxYHK
eykD0GwNc8sCyib4EosemdMSBUNbv1i/j1SDGXGztE9eqLTxMHkcwadKsIM82Eb6aWcoqExNExwC
to/nQCV3S8KhiN1p5rRLWjOSHHOsJJr+iOZ7KDjhvFGxkGXdGQNgcEmSmmA3BPMazNCwPlH/HEh7
EmJxUAgUvaV8JZuW1BMzsuI5San7mlQNSW8WKJ2b5LPHHqaYUsokib0wlsRVnsL+wZ3L2SkRYJ57
kZEz4DIph/qMIFe8EbHS8qhyhLRlPz13LUPrk6vRcWiJuQSAi4jXltFMbCVrUN6aajhClptSPRrD
lZoHjJfy1HSi63+hxBEPgp/uQK2dQyJYipFYLrDwB9mNl51I9k8Y5d7XeaSyAbjH4a221p2b8ATY
YzW6A0Nj0Emj7ilFUxvxjc1/2hHEr7Au1rXKVkGBdy34dDa3c1ODb1rJShLyrYVzsUG61FHLrG/i
cVZhb6p+gLAfFLR/3ymP4K5C23wRemTeWt7p53m4U6uk40ukHOon6hD9k5hyCqu/KUzNEfjZrNKX
4B+FQzCk7n87Uz9W6/ZChFdFTslUfIc8HjIlvUggr3Cp6HcT3ZBClSY9hIYWgOMg651A3TSFUkzw
C5ffKHkS2ZVkLhK9Mt2dmxVmGamdhLsLGgxBNO8rM0QJO4uF9oJ3UHiDOzwjXyMrOWY9jlRKg7P0
/C3awhyloD1PeBiW9fFpzVqbnwywXTbzntfOkqOkMelTuFAMKsGmIOD/wnzMEjKfTyX2y2JiGcAZ
6ZWcHy9E1uOMnCaxQlxFJ3j1kcPuqBcWnrm8XW2/jpTd8tX85MIE/OsXkKYV4txg27V/DSUk3MfY
0CGCG3KOOq24lpuEVOPeyYyCT0FHq0uST55xKffpCCj5KAtix8XHURk8xTu9T74rMrZtMVa7hauJ
JADt68+pln3y17q2y4pz7cZAOkhixgUABA9uc9DB1zE/G3tpRPovAkuq2XXHK+Tmo7uevuic9gx1
4RNdnk9s2lO/kK7CWDjDO/w8kpRVrYBHXhZEWTxarzOYQ7/8BcBl/0nZo6FCKlpEwBsW/kzhjeOV
euODsCy5GmgKP3m2cva7cy0a10xJ2rybylKupwOAwelWtwEs1SS+sfYuUEEpEB/SA4gVvzk99ADF
iXLK6W72eA5zCIgMpE3/kXUpuJlGFke5TK3Pb+AwA9YQ8oZUtOup7b5OYmQEP0AzSfgZmssM8rge
f72xsbBY5y5K1kxUFdcyXGuGOCpr89H5k/0Ll28ZmDszUyvr2tuepmw8BxQ+8cPjQUMhy93FEStD
oRcv3E/nEpUIrvPxjSqwd+3hpT4A7c0GtuNS3lEj10OHS4lT8Wo+EZpExs4LmGOjBQ08pV9zg8a/
tSnlVOB99lX0EWC0zAsikWd/HCJlrIsqC8jpdUWFJ6HM62dmyruSZ3I3OKvImczYXp2A3kelWlm/
m0n+Au/YzM2bpwhY+n9k4dGkWqxHEQA3GJUd3m8bDvaynLb+jDbXnpNztbruuho+HZVaCsX8TXns
DDWTti1iAwx2nwP3+MVA0MZk8ifEsESrS+YU4AY3TA8qqLrmvNDWvRm9qRN063pQki/0viHkZtns
bYRa4Q3J3QJZmbQ1XdJpo8mHHagvSMENUjBFDxaAlj0g9SgDI4gvhTCZI1EdgNKRaX0H4QJWens4
tHc1JkkQ+eddVSjJge5W93EWRjKOL26PtQvFJ7HXR5Aj2ljwoexyaTlecb8ck0Pcgfdd//A01u3c
YaauKnczu1NunDQA1hSszgWoRs6SzmWXhM86IEK98QND6muO2J/VrxdXlUe8OWgLrSlFXGqxPbxo
RrzR0V9LgVGDbIssZsIjhDKBDaEan6VzWwpN7GPVdFffGOIaZFXzGTpWnVS32Qa/D1wfVExtniXo
F///gq/3H2b9V4N8fxRNJUW/TS76jzjBB0OXhXAx8pYe/AW86dqO/DU+YPjrvFi/NZM3Pwd8BVVu
Gmix+mewq8xSSk4JLoZ4Y0J/iohCZYXq4/ZeguirRvfzsEhGFE5MVEOpq2FdFUV/dInyeAVxhZSM
Ap/g5fK787531qHwy5zlRjxkDH+NSXB3aLXnLORkq694GOsNJ4uoK2g5OTKhTkxP9k9iqFjC+nqa
EcObepHXMHgSIVbLkw5jBuEwn4bZkWh9W6lVGjrBb+3Ui47jmLKzeOFG5c7fPTj5dgLONufoJusx
9OQLU5BN7TgD0/C0lh3Kb+qX5TVF602OMRLihYIUJe+nAmMxepdaHN0OJxJTtCXVzjf7K3KLrTHJ
E3c+ajw7f1aZ2l5o+ZfW1PMZcApIyQDmkFJx2B++DWMdUwUWlrY0J5QfeTQwZPTXSjVbwifwIol3
P0qruMH78i3DzdTS83ev5hZxNIVVSuQyZfQJ+VZYVojunRKzEVMDu1Ja7zsAt183uM6yapfPVJgs
NeU6Y++t2+5J7UndXwktkAU6qD1thf9N00PN2ojzUSyc4Hl8g6dIgg9awhI+RH54oR9ZcsXIP0oh
J35cNqYYTbDIfD7Jvi7T7Y+7WB3WdxE3kuwEjyBcwieYjYRxjFYXIigRmFAQyufyo8DRlJq2r4N3
x3rUUSV6Z3qw6bMPJo7LYVv3h8qG80mLZOIueSaRGeT33CjVyEH2vrf3rIxhHHwHQ6MoQ8HPxkru
PTKnv/bp5NfudCQduIpJ4T6iyikVwd9dwrbOWklh8DMPQJ83ibMIEr0BWWmwU6An6jdwNv0ySbV0
DXmgYdbPaGu21pkIl5DzOrI48tiPZAW8EBrazOu3fw9nFHi84QjqU6/6759BVxy9hlRGZfDsQPiA
YEJFcgKY3m1Kr1T7aT+W3Hh1aHSi+uPHcEZZVeP/3nI7lzPMXKWlwH8mMIaEdUt1h1f55dAV3sb3
NQK91tj8fLoTJZ8NHSV35m1rCFCCIGRZ7SRjPl/g34NXwnQRO259M+kHCgX5TNkzeY4MbSA7B2UD
Dp2FOwxNALj1sajIpUwzOcpJ4giiO8rBsbLQtGRpMOFqdqI9+2mMfAiqgYMEoS1rKCjx5W2a1r8j
2wqR5wyFI1sLW7Qixdjhby5oyucgHpJ/BuRWAtjMuYnqpt39PCS9HVQXuVPkuawARQfzKO8j+20N
CzO/ctSt5jnHFIogfs8CKepQg9ccMbNekn9Pzx561/EG8Fb3t+QQ8Lg8vvPhzRJdIgUKYtH7pgpr
nwLDoAizaJ4ok3p0/WN9A/hmvNSuGWaZyovHMwK6DLbRsDiltxdiOSDfULq95OUfnD6QmThWey2d
6HuOCcQGyxnnjyHH3GBQpTRM9RQM7SV84EQ5K3ysFsGMM29ExOwik2H6iluKpn3PM/mY4Yej0Qd5
TtiY/0+8TYeJtUrkUNm00JUzjPVGAaJQIGbTTB5OmBhavMd+mTpySwG84n54llBSSIisvKNxLMem
LLqiJ0EyfcTtD/dy05ghv/iJ6/xYccnHkXs5KgjSWF5qDcG/+5XdIlpjZJ8gNYFN8+bmXYGeuygv
yPpFpd9b/EvRo1GH383tOn12SEBKBmxy8/4vrghl+18bTfgwjg1NpTlgr/wHF+PKBv7Xx2Ocavz2
tOiCd/yLWlktOxX2qHxlXFcXwjh2tSGhWCL2BNrFJcOQeKtWkvdEp4jIdnC0fU2SQfZNufz2d9ro
HoyaeF5IJTiRehsYvwqCI8MC9hl/YJsV5h/sjqegk8PLFqL8WG4mIBnp2R6J5D74J+xjW8Q4p9/M
5fKV0ehXC3aMH0x99G+AnDvpFO6WST3C9Op3BGxlE75tCS44E5c9oZASm1STzSdJMsNhTwOuj+1O
qrCZDaQzNsVY11hc9VUCrMyv9AyowNJAfGjj1WyLwBwq3qwoeLPaYCAxJoM5OXDfXDce9CMXd0XA
KwEoqzHOYdAiZXQlrP8s5zm1S0P2J2jK583iA4Pw1OuljEtgKRTtmI8VWEpAFPGhq+r1ik5hMW4h
uBvaB47QWfwO+Yb0DVNpSkf3xao5yfmnJmf4bKf+UAqHpvlaZAYQ74V0lKfO9D9PRoSDQlHIqg47
JdWcqDeDwjFXROJfrE/bSWPOyPuYbiJ95301NGgUgjqZZVeWZ6dGN1tLwOa6w/yxZJibTLGHKO/K
678VP131OPjilTOY4+KbqBpXS3PYsDeg76kMyLpKCtdhL2GddPvi1+SFOdha//+ZoEIcbNfN3p/E
5s/TQszREubeCw3jmjftnTtb0zPVHEkjOElFF2aixwXMUXsr4Io2x6KhlNLdcUhSIaIQpNxZPsgm
3x7a0DWVp1ygmJX48prIiW/8LKnqTSQDw6q4I3yK9YyFhNOPku4amMBO9LC1Pktz7t0aw6KJO9sP
LjoRoaB4JCzZuZ4nLL1Bz9hVmu1lLDSfBsO7R/PKIJoP1eC5yDSJjK14Oz/qyGSc4+D8M/dAgQpA
ARZfPYZnlq830E3reW+BkfoxVq37tQM/rIW85S3jtEaIUPEfXXHozG8YX+kmKaoFrfO/Sedlju5h
JejVFERIMW40cQ5Bf+hl/ytwcCekO6wCfWUpoQVmqa8O2YHsGTo4w5ByZyduLc4dEmU+djgYALwr
fnjHyTU7NtSpOwNBz4w7gP8uNOId5RoS9L23or8S/m63szxXzz7gJdRPRORtp7YqZH1ILRlU6OgU
Z8OxdjNVanHLrN1BMDmviP/+fRVT/OlFDkSON9wnACChpMVmpjQwydvKjnRpwwBDhLWam3Grptpn
CnBrodp5aBWF7189kraxHr/ckH0mc2KUy7PoWDE30JQLJUx4N/9dojwA93rS7or8RpBSQpD8oytX
Otud/My5jxFAigS5VrnDjTQau2JNtt7ZWBUoIaX91u6U8yXd/T4gzRJiZgtO9LMRHCwF0X+r+9cl
E/cN7aMHqnI7/ybMYShONGR06bH0AzXK1qwzD6l+ySM3masvSL7oovqgvASKY6tfwTFcfsCrTyIr
HApL577p57ANRltXEeI5SCnBGTsRsWigUuLiK5NkagbAT+lus4Q6a79PqMehQsxLaoG/2rPLwk+N
4heNo8kEtnmW+mCF+wspVeQr02vn5FvTU2xyW5YCabEb4ZAkBrhkTsw6hkE4+J7bKi3/XTnFJWob
N6z/sD/29wjIWUCUBeeG8CzO4GEubeKGnlg2368Ti5rgmQwPUOFxIodqY1fSRDX1flDR+OiJWasj
Np+dBn33Kb2sH75dAdTXBqJYSEtuf5KvDU3Ql82vvXDaVorOAdomsApbslqalZ68tnA4AX/BWtKC
SLNyi2/cEAQ7II01DDNHJJ/U1TGFGxuImZ2tZdelCm7NL9P/y4ka4jdF3DUcqYLDYwkhmdTfuU6W
CQVN+QqDx3SQ8QDtNJI3d50coYxGaklDEiHvgBJEHsMOkUWVrv20BkuStEOk8gHeI8wDwVA2yHMD
bF7xMc1FaIwL9wYmt3/pyEdHWtAdtMwlaltbjBK2ktYtbf1KbagZm7OYl4oj95mIgXbsXG6dDmdk
a2dneWMbJtjfn5F8pt0unecPVMqTyqdVybG01nY42rLU4VjVO3yg/CHFaxwi6WCMQFQl0faiy1/a
0Fum/0fbmPdMscTBjk/99HVtJzErxZ69ScugsCFUulCIRoeGBN2r3kDtO1KowWqP1IRmtMvXGFzw
/OqDwv8sWzVwISDdS/L1Xn8IQojeE7pYPNyfVROQks6hckiMkR+IEk/VuTyS6fVufyDC99mPx5gO
jOlbFWqTz/nEoKKGJQQnxbQQho5LaeZrzPATGrDioc9dUaqkcGyq5E5WwWXA0w2e6Hn1gg8Vjjw/
P+AS7xhJyktajhTxf4BfHOky2sjRnEoLfujW4o5hLcPyPph3ReGOtbwP1W/xkHY9aH+70zb0lET6
Gol3bvOSwIlOkx112/fT/U94lQyB+FURWiEvxlC0sOk8+ZH4XBs6rWtKl90wmlXgi7+5Y4XH0zN0
tUpUmtTVrhfVby4riMLGD5kiPk2jh0ezLOFfo//Kumnvw7AxiaBbttlHh395paE73RKtyG3Gr9x5
DPh6edSfOPLVv3x3oj4OA2Uk9dsmOY7FzpHkNWgxR2wLpXFC/TGXKpO3eMtEQ9d4B6Ovo2otO1p9
/qkNP8AYoNI2DQ1GDQU42Ymlx3AMxJT+La/5w7bZPrQ541WnApm5+yhP7IVzDEe9aC6Z5W4IncUp
sXQjLEdZ84BbBJZ/sq0XLjE1SPKygBfcbloQ9kUGaMPeZG0WZ3DGEoTDlkrqiMsdQFHKaGLi2/Ri
BDLkOD4E2AUH5YcvrNdABV/jvxAcTAJwqbTo7ZIVJqIldk8uYM86GqEKK4oeopN9PAtmlw7qSVMy
D0nBbiDKCEDW8/xbm8YoqK2qs5NgTxOaex4pIQX7oYpC3iTuYd3+eQ6cImRtshQ1BpG21JOX1hb2
v1GUdaj0tU3zi/LiRwMAxDP/r1+G+ThN84rd8XF72guYsbZ1+j0kVTBdocmX+mLJZkoal3A2qMED
TEfEt0j/PU7d7MoCJJFvWceHYuxkuRzkoOp9+XNkxmsAEZVXnut1fBHAyfKkDV77/zxcpqah0btY
9mV4eTxtni1TidqCezzpShXG4nNn77f4veGGDzeit3r34V+MH83l3D7o7FatlQjBVMzRmtSg0ptz
JdtE7HkOBJIiTMMuIIyXyCuSqoye6zYS6xffyzLTqBqpdnJzxhvpi8zFLv2JBYUAyJL3BSIp2saY
ye3fTjgxkMPJ4uHYv6CVbaMOx1VEbsg2/Pm/fTm8+mYXlJwbCv3M5b9EJXMtixX67YCwG7zvXAkV
7JenNPBHxtz8p7AFSod8KXrfuSh2avR3jv/liDqvGjX0ZMwJIzD7V2uWSi9nxHzrVBKL3W55jQKO
H/awrHnJ3iLLCOenYfxRn7OF0Yw6qzzYAvy8eQmlIoa4brUbVQksgyyvOq4cagls6Gv5sV0T7/Ic
dL0temiQNGJ3vdUGJzFvkWfgopxn1jcUB0kvdKM9Cr4ojIcg/nkwrzD54VjpokXfjryLsgMagERw
oFUMCPWYVm3uGj+GJ/BN/buAuGRt79sd2LRSB2nJKZmPDZBqLSKMIyIIMola9V2EPyR9zUgV9bOq
nq2xq5sefPJJ6YzN4pnribfTqnoqB/+D/vluLW9uM2VqpZ+vw50x84lnvUVDOjxmvH9QznewhvXN
9dCPxwys0Cy/co/7kCOZAr0nJUp6m7DWvD9+Zbn7mlIl9u5Q5ABwHpTbIME2zz+LEpmKb3XJ85Iu
zeYbJyMqyaI1pw6eirVRoboBgE5NblPFBM/57hj3EWtOaMb0xGnsAKRQ40K+SbCXB4Eg1Rmr4nHM
1ZRoffqgNg7X5LZS9mzD9r46ZrqE53dwEqoN8YRN/x5N0qNXqXi7zdEYzRhU+h9BFOeKIhBbO3mR
I1S5QLwHqkNnzcUXnGWfNYw+bFUYRUkUG25rQnfUQd4PWxt7fK1oUkonqzslk038ivPpcyzLfFzo
P9ZDQBQ5fMKV6VhHT63hfoaJF5sF7neZf+bQ128tIeGofNRSGRYv+XzaFykm0Ifxkw3+MzcmMuPX
SA1KFvM7+XQ+lXBRvnUY4/HquT/C9gK9hfkR+Oydosc+kUZ1alMHLDMv7eIAeXUY0tMStcs4IotB
OVVpzf5A4qCEMvzkvVeOKvi42aYgo6+gG0L8+79h4AIRI0s8m6Krl6BM81o46+IWaZE420b2l7/7
LtAKwx+FB348UFjgfDwxWMBAsriyJF/vhLnYFBv0rzYWg6LdgGSZaKiCw6p4WZ+Q8/cxl3cDC61R
XsEGCCbo+TqI0xKxMF3Q/nfburnYtl76Go2/WWi49i9o7kt8QJX3TE/qR9gO0/O6PvFvzXYo78bQ
2yQpcIBQE4Axhu8UmxpzDTgis50rtt6+cd5LyQh3Vite7dPM1oR0aKCihfvjGjJ1yIQyo7vdxQbi
WaK/qalStdoPS/Vs1fmhCarO0rPQ1FTJkT8xI9hhbABQgQ46GXtgqSpf32D/qhFQlXNkTJQiF3a+
p3XalaGJ6TbLiyxaUWFoPf+pyk2Kc44ohRcDbtMIYjVrLvZeQnn+9T3Wes3uZyxszwDeavAatAV8
eh8A0ilFd2lM/GJVjQk5DJA5Zlvo+WQKNsVbqUWIATM5xh8tNaG8QumHJpmKzkjGgRk4Lraj4o8I
pr113CwZfo1669BYmpefyj5fPc+6r2glSuLCX7SnJ7fg1sSCnftoLjwgBQ2nSa7ppis1b1x1Z7O3
BcYNWU0BzsTu3y3yAgp8wALnNJ48ohyX15oK/B2oOhaGAx3XWupQpjOAx9JQcPjDhLLVdvSiCgPJ
fPW+ZlrNKLO7dnaZLRJveKFAXuvPRZd985XWkTRt6ldhCLWW93MdTM1HwkMAyLZZEz9XoKIYVKK1
TZyMBMGWoNW00UHBTQx9j3IlerHhmR3hK8F0wUW69sV28TVc95K/bPrHtf87FiPvdSzQtct/WFHt
LzCt5//5Eo6Ri27n5sG5kLRRpF7w4uagRtw+BAcedHaMOk6fZGS/0cYV/hfil91X1elkLXpKPNN4
LbV5BnDon5do3QXtaJzHfBRpMeB/1qYcxuIJxFlJAnXYwFFQCW2ZRYxBoLTTjnDA2PIohFimXoiC
aGFy03zcGnRAy/oY47ur18oQZpW+mQTFbugOVVhr7l/jF8c7AZ7pJ8y6BKwyBI2QKi2pSvQlxSJo
hdHUz4NtjDPXZ54z+polyx7l9r8hratirJAMRBW3+EPi3BPVUatTHGzPzBJ661VEQGSpGUn6L9eq
jGXpKOVCQvRy8GvQdf559gtpB9IoplnJkJqWnXmjk4sbqMMFRepyaOAo8uu3WwhQtIa2BUlDgRde
kr97WuOpADu7cOZHYR20wsyyRTjZMvmqNtiwCTWT7TyqWk1dE4DKblKK1cVLfIfj4iQlIBrYi0V7
AAVz5K0+UN8t+c15b5hnwZgzAnIBwvaYJfjjORMqkPFzWA0HM2i9u8Y616rjQ80yh4jCes6d4xNm
KNtNM09Zm0yaneCNmul7Rp/rJKI21NYZs45A/y9jqBlQp9jCrF0r2oicb2wU288sjKl1O+ARAr3S
kvlfQK+gun0nPgJ32fZ9uOFNc8ntnJYR0c7xc9O5/p9IdetF+nQu13DFOWDTVwrEBBWeJRVjVj0b
xFKWWHGDDhkwWnIKF8+XaUL1JvR1DgKp4MIPv9wx8N3ILeL3lipGlk3e+iTCXNBgMXqcOLPIQq/y
g0ZLhiaV7Ml7DKarMMku5hEprl27Fk24zAD0+hc+NNn+pFwkQOgUMShuqq/tGrEOVNmL0KopAEGp
v7+CuQeaht5T3BHgLpMc9SUPyBNRWBdkz8kHbBTmTEg7QDw5MZpCad7NgZQSqavbLzg7EdO6WBX3
sOXt4dKPyHhfm2QQt9oxRZpeKOeUKWOFmvXERNdRwOPYmQYT1S8e68r2GtPfVI7R/RAAJ+Dbkwbt
hL+GBVEiqSC6mngZAArL1atnLS9SawWJk4sNXLV+4JxwSX2e4I8SMiefhEiMVx5mKsNfHcu2cq1m
Z8hDBaKR+fqiEnoVeSMHJR4ABwEDJr4LU96yoOrjIDxnbziZ0ph6CGFLJHGOZivogmhO9+dfJxD7
J984h9urVuqr9BdaO/fykRAiJdduuO9C12/euUprvn0JMpE4CDS3S2U6ktDeGItZ2O0lnzNq6N9D
NUtVMLurPO7Z8vQLhAHidBqaM/ctVNeYYkSI3HKbOtoZNr9VE3kQe3VtFL+q+cBSladcogjjNfLg
UbzJ02aYj99eXRHhGrzdgsVrvo2shDpLy/53t/atEPVL4qqqvRqGPxtk1lRTKunLWBCmM6q94eSO
fU6zOvLH6wPkh6KtHtEB7Xoik+GRl++aiC5JBQ23z0htlLhSIyYSiqQomI2KyY9SKeD5vhrHEYS5
faViKoswW8nNBqMTLopQGEUsYs1uempFXDsPCF8u1PWjDj4Is2B+D+M3drj+kgZ0ih5gBJXx9n3Y
Sn+jqft23sxyP+TA0/57/Kuogx9q80/YLrZigOzaZZvEjzDCxAxo9rn53HyPmuwzeVeoYOlBFosd
TIkwk++d+Ggr5yPpZAO0NOdcXvFpzSTj5IOvs+cO6POeYL5Jdfo0ffGqFGWiuN0UtOAdpHYFgBZW
jEcKt/gRiR+cB07WfdatuWyl1qzGojwZJ0c0ITGWKF9JUuVuy42UTIZqR1KPMryNe0nKUxdWmZUa
DF374R3NgtXj30uU51kF1HknI9LlvO0if1ZT0o6Kjs3uNm8Rt2bVl7m8XG3fQ2BR7ERCePhkAURF
36KhiS6AX+LNM7MPzk/5iBJxkl/nGqd8kYn7PktBqcLo5+6vXeadYWKNZSthMmjT+l6iJ6izW5bx
1rX8ulKxxg7vj2EA3wyTr4AKNNkulTmQEDe+Kwe78bSui2iqYKFu4B0N1ELA8OGS3Xsp5jbN7Ufd
nCVPFTmgbsh6s5vhkymCxfij5zMf8eXWwQaNr7bLPcaPdM5nl828s3/GnsbkXr9luJ1mM5u1LcXu
CKyPPCFSwd3zCZbN425Ha0ri/Y7VGYbum6hWXsYo76xy9Sv9KWk8g/Wf04Z/UscOwrLcmlwJMXgN
QbGvIy746GPYmrwLkRwWtNjOEstZEckQXuW/ukpe2dbx5A98bPWVF1Ahk/Vzv2tA8gi+/Tt2J8X8
QyW8rhVzCrw4cE6W6M/12l2kd8IKGRL0c9G+sVeBdsTcbZutFdNH/06PstaoXN9Y3kOf6U02zRJz
Og4PANacXUrsk074WCV5TbVPs6MqWAyIa5NWBb7WC9d32ALwheybMQor812DqeTGUZNHjgZf5744
S5moFICSs/SndG3oDzLvY2FQP6ZWu7fnO+N+wgwOCO6HW4AwMlg8JzVAm7lqC+SQsBMX1TOGxkbY
WHbjyuWQ6tQuDZaCjS+XgElzq0IF7H6YwAYvGUjSxFe5oliohs9jFt/+x8HAAFZwsp3jPYLM6n47
Cle4HrsiqXBhJ0KvagVGqtf/EeDiAPJAv0algPpnq9c3fg14UjVN9gJDFzmxOEL/qXbZ1PrTnsW4
HNrAx/KSI0EVSBd2tnZN/DYHSSpHZjJc9sHM5CTGwg1KAPLm/5Xqb+7REuMSpnCeWOAhiXX4xhJx
kcP3DQOESB0fxHgVcrehQrUBiGSe1JC9TCePDFoZJDdIMtj/OD0EQlgDCrygLJcsHZLSMxrtLRFI
KsrS2OHBV2TtzETBP+s/C25e/QUX7H49NJ5sB2fDP3olOMGwmWB+Xios8PadtYE+c7ZTu6JquZpV
RRHH6MDQUuwf49R+mYmL3De49WtgcZdHSu8/VoSejlwIfMChNqGJRG9dNvoN0+3cHDGzq/FZcg1B
cX1uvka6GL06QymIHxyi3BkMcvoYvT6OKKe66rs0x90NXMC+pTLSzlww5FPpJT/aQ3XvDE4pupsE
FfXo3/mWw779yrojU9+vYpIWvoPlGrmhyQJmN2CSwrJisJDQOz33nMRJJBRjpuFq0E8NK4PnC/BF
Va1sTsrbvKCqznZ3fOnoDmuoWqgaIXvPEUETUVcFkhOjluwtfcIW49SPza/YDDjTzem3HkvDu2U6
96kn00jmfLsA/zRGqyFNXFA6tN3iqfkVIgGOQedfmGsuU5FKp7PNaWnxcolgopmPZTdz960I8bRf
ebG+Nhh11E8dITlY5GmdBlz0dQieIqYYZFWfrJOfCjOpG/d6TxIa/1HUL4+vLTQgexheXUXgEssC
LzCzHe0VY2JRrPic3MukwJsttdEkuvKwyOuURFFRRN9Mh/t8NWuyuD3UbFE+H+CILTfajFeWBnLS
M+qeuE2/bTeD6TElmVDFhynAS7Slq4CZiWt31gL3L8DOwWrPY/pMSurNkn4027FKxk1ofR87RNvY
Cv50E3bHgvJeolQR8lJ4K58qxGIqU0mpMUJwNcj9uUO0vQCuYcu/8t0xVjK2lC1VlyWAg3GK9HMz
hKAvFPSUksvgtqHZMajFGTrXsrqLbf/igyI3DRo60aZbZBabsQPQe/c7/iUbhSSI04n14qjW50pw
yImRsbzJAOg+F51MO7rzP7UzUibgAwpcAi9Fbl4M6Y7yuopKqe52yQV7U7+1Exl8dYSKuusip5jX
XYbzO0klmmI9SY4TqJJa/ReZG1gAtm6Hl6DhBu0OwYg2i76VVOP8ZJC72CeDWs3d2+XNw4hhsC39
Ji0iVQ4FqAytF8fCgP2X+Xvr8F4Trtu6P6wvam4hbDz2Z/c7Ty8vOzYGS5hviC5BSqbGJeaG6Lpp
g+jIQuOircSQ/Z9T4wdPLtxo6BvjdIx0AtA95PcbuaZDhlD8Uzrsmj3ryv4cq/hFt6rw3VjbF9ne
uEglM8RhviIugXjMJleVwHand6s7CxSfWTVwbovRllVProem7ml14t2NdRFlUDN0eNQpxRNiYoYe
LzM6OjqSaZJCnEsc1oVaXo5jui/0WxTC/jxkPxtfkRJT9D0dKZXiORUQSb5bZSbKA94aURMuH9Sh
pJqiHtlumJTORVx/TcCBsRiFYjLQ9tL8nGzxhC7DahxzRbIQwbic2hl7Zs2qc6hTL4rYWD3hXcJg
c00ZYytv/62eNPNsuJ29NjmK4T+eulEceVB76um58eEiVM9bz+lMw8+J7HBIYWMee9QNc0S12xTs
D+yh/GOSDwQixVD74OkfgkRbpw0eHY8WvLi3BkiYz0MXMzSMfXzgz5rbGzJV7jQVYp97fseV/XrZ
Pd0K14fsGQvVYsHBncFr1nCXmZmafiwG5mYvtl28Ox0cVKSvQyJUEJgAnZeYpART8nUCjfxYqnxj
EzrbUAxmEzbFK6ZvRrB3rcB1NV/VD8EzvlMqmTrVhZUOlrh5ECSmvocKW1b4xlkuxRaQaM4tdE9u
iaL3uCqoepMipEko40qy7i1vxyRjzLXshT4J/L18IU8XCadAsxUovaC51kJmXTK7J428r+q3Ud6Q
NZrynYW7ARDeGuuX2HnOA6psu4KjplwLiSgerBUgB0/8j/Wn7K0HIunCEFEczVNNU8+BHTbFtwl3
USJXPm6zjyMElOEEGoedkRZq+avzZoji0BUZmYyHto+vvGuYTHGwXfM8adfNuk5EgOWbVPggn/lu
9npbD2l0eT4f5pEPoRA0+5HVLWSlwhWNkBAxHzNuPLxV65BRmiXUXdjYwiulrg18Qls+7MjHNS+F
jWfuOF5bJWJ6Bfkvvqy6bn9BVUuBjVas8rmvbA3Nc+EW7+vZTH2hD2MITXlinmZrbD1FFeiYsxln
U0CgGNMzep9m7Fg+DgIawLbfz4EIEO/D5/HCJArgZrOsYu/UNCazszdhDvy/08boxqzo7aycUk2K
ONkxjgfoFyba+eKdf7WZVgRXoE8nz8QBxa4wOOjly1venvNixk49p2RbKAd958LT2UEkWr7PZLK6
SJQaVQa35YE2vyUCoZjRQV8Z6dQoa0xxGzoU6t6HqWcSttrIrmfn64J5qB/fB2RYBtEJdM/ew6fA
gNmIkoI6cwRSXCt305IYtQ3MrthW1ss5bnZu1Z0ARQjKIFszMrZHJrYZAUy7OKPmGjD2Tn/mI21B
vci1lbsrEBX4Glt0H2vH2/e3a99xy5pBZqdgSzdQZ4HQy1r8vUB6uOaFMF3iL1j55ecKfEVO++cZ
pkSb3x8MQ8f04mrp7gE7wLXp21HDYfOVPLuyG305Ae5osYOL1S6LMqqx0nj4Va0nloUKD+bWeYhw
KQUgrc32nKu6STPHfxwb1xhXmE3ogDxFWvme3TfBkZktCzWHskj0QH4lHKZNLVJ+qy0HPOFT6kA2
9qzk5oOQjpBmqOUj8w1W8Ge8bPElX1YsIjtIDRO5ebjDAhn+QUmCA91z8eUE6ypsVD/xwaoY+Np8
P32W5wf6XpFMD8GWgg1SJg8xV8E1dhvUrhsu3+7V6an2xncChbmftZnk7SFjVxhDBS9qi5X9VlL5
SaVnskuiR5cPjks79xOhukoFdNW5jfatzVdBdv1AyvxteA4ohBXMs2GMpBfgr0v74WT4Ipedmc5N
BbY/NJ05Hk5vAO/ytokqv8e49sMM9PYoqR4EjleSCMqfCB8UaMuEfTTHaw5nL7tsTm/8rA4F1otQ
xsfqMUetCiS/JVu5SN30aTy55jhFthiubJLx01XjeKLqYLuWiz7Ztbz5fzH8KSZxhpwvq+teAe4a
JycuS0+JxnPHiEJ1LwaABUXjund3cA2YCRz909zuTNaZ1X/+0tOG99ar6/zl9GTwpTOc6aO0FQHn
bvjHsA4dGZaAOg3Y02gP/BmaEJdA5F7RCPe3Ekm02woKEG7F+XsdjA+HqjJfx/G7Naik9PFFoO8u
L426VPlDjFHyvikq24aw5dtw3JQCK9ndA1jrIlmJy6xHYihWZeszQ0WVgPO4Blj0Ek5Pi4RfDlq4
Ms00nnRTPGg0d0H8taUv3ZMc2PHBWo9wFhuNAVcNiku8NyaY4DCKab9aajNFkjNEIQIkcYCecxpc
80+cHjobMs/udHd2e48xgPv9TSz/ktcPjmV/T4eZfIjjHlDcYEonDfiU3S+EaB2BebIKzm6XCeNV
EsjdxaqSXjqIirGZ4yHQBBXyIoJ1KCJ57NSvcavPFpZaDE04hIYMNDkZpH9NbMj4B6ZCF844hpJA
TjR5gbSh/RYgPPnNGAG2OBxwOgORWAZPkNf6aVHUIQ9bNf76bcxkQvD8GnMBjhl2DhYLLTCokn+1
un09l+867rhpLv7dxw+ULcVufiyE0MQQqatzeU5s3FezUry8urXWoeLvzoWp1huKLXIKP8drzs/6
ynvKANN6ji8awzKuSiZ2IfDtnfMp993apvk2FCoaE4c5egT8tl1t2jXff3D+NW4OOfVbboA8RVR/
NGC1FZM8h7JBEyVw0bD0XyN4OiOmWHmx1y710p1Faf1sJNLyf3UhHaOl3m8o63qEXQTUwXmUVE0J
3N75DFyi6gTrhtgni2e9mRBJBkkzjKuxyqw0si8sRaksVHPbxuOVKjblH9L64DnrL0Dh4DlaCeIo
AXeNxCDMM6WUaEut9g7Qj7akcv7XOI2vHiNSqdJjUEHNPvqFzTebZH2OLKnvh0xvbj1BRHzQOsVb
KM/D2qrmOQDR+uqLlhMPDdUEZpGyMR6hXsV5yuYmAvKhJjg/DwOA/vMKcEdlgbPYhdST0tmWkVJ5
fcvcD/74Jn8SQVZj26dUA1l1pIAI9bn+bPW5w5UVEyQp/CnM7ntp5DPdUXtQZKrcmFESqxZiB3Ca
OByX4LI635CQhBxoVgQQstibH+1IBEKWmquNGaGN9bwEAWC6c4S2N97NqYAs7CYZTHVC3qP62nfY
GyIR3FT6ZVwB6vqT+QwNZsA9xM7PS4/Aq6Q3F8laWFMi5rHWPxE10XKuI5u4zAU6oUSWkIcs9kiy
rK+Y+1rzgMzGqCwwTSYD9dhS+jkbvT462a8NE278jPtsb8cDPtXbafcv3i91z1aNvIMn8uvaDVDO
8Vm5Gh1EQBmPAJRRrgWONv6ml3KbUYKfoZVfAY0/lHdzpODk7DxJ91TvdOwn8/HgZsq4zSINZx4H
tZtmSyXOsoc3EarTxMxMb9hdZxEYeRBTIcpi6AP9OlIdmQibpjs6xd4EXxUTw08vM7jQZP1NRuAa
vy9b8HWl0Hyp4Po//zJ078rhpe4u3z5lQ/mI8Ixc9pQfgMdxZ1oPDA7AVJNUsPjQMRduqOL8QWYn
KHqPmSzgY9aA+6GpJrGpvb4CnO9rfN/h+487oF5s5/g64IQwlOVnJtjP7jhP11hXV3W8GzKfSRs/
iUFXmRf8MP10EILflxQyVFecvh3MzeS3hmTzPhTW4NFI3l+EPPpy4buWIhBvFi2eF/mqk1jAv274
fCjHm3+CzPJXmAQwC5RvwNN5iY8Fa6hFJ5E7cSRz8TpPimGY9mC7RpYDPnHHHqptN+6YqFiNvT/I
JeLpzW8UpjJhDo6ia0f50S6JugETFB31TeQb2vxQ20K+AFTET8Uuo6SHRiU9/pCL7X3xey4oC/wr
iKjvKS8QQ20x9iHeZ5n6BRX4NBht0UKCZOQCwBhqMDz6w7xolww1BXrdYgEIbs2sVxOMmu3U1Uqm
sPRDlgn23hgZwz6k0zXSDQuOSkPRQzN3VNgZkct+sD5JjzSKUqdUvMHI6B4x88oUhtUToDzGoICv
6aMVAZjvof+WErlAcXVTR3o8BvGZeUtfEuKJE+CWXUGc3hXH1+XMOEmbQn/+TFi/LrGAXsu58u1y
wNBziVfKXwU/jfEhvWswSgLHwhXYKtgamZ4MsHx0Fd6oXkNasj1xhs60PbmvXDs2UJZxvj0labm6
nh23iE9PErbFPqxHP5ZgZ8bndGunIqt7RCCw8Xfqemi2eB2673a5ziuhgxkS74x8RuRS7qULAamq
Lr1dfmWnkoI3dymMH3cop/fPj1GGfXY/lmauDwmeE3iPF1P453vLGXVc7yr/qlkKzf4KigVEkgrc
UpNm6n50G7xdtKEN66bDGuFuXWkYZMp8PrIdgnx1N8iWHKXsGna7wEESKsLt9BzkaJ6ACDiTsNJE
qHUURledce0eFIpoa+U2rUn7kl3cwItFQu1Cb0rLMSte9EiylSmyW9Kk1DMzTWe3fEtZd5g78Rjt
DcRkdfHsUBo1U2TWiGwoUYUduFbc2xT4CnCaIYJSe0MWCPPj9dwVYtDOHyf6QOhHQaqBMHKe3ADw
FWg1jv/MI/2+oS7gmbp/ZIxTv/3Qpk0Kzom/aLYFRpagB6C7KvFM6E569zDZwEwPJ1aHf0mxsfp2
RJRg/XdBn13XkuZ45FPexLYmc8Uqdm6uqdvJQyrfQINI0hFnVAdcTYu7jm4acdECoSQSOgvGCA9l
p9jVF7bToZJBHMPjSkRNjLUnVpACJpXQrAtCE3EUER8Z5CeYStE9fzarRrPLAvC9+95vBplrKvVY
4Ao3ofOBHkzTO3M0z0muyr6WMcwa/7fPp7aQRE6U3hvznVfStpRfSNwUSRKBoPjK6wIZzX1XuEPx
l6gvWtGjlNqEUIEL7SXEZsRxTNRagR4PZMSNLPgkvwOYuPOQ3dkqhgfBKFTkBHbKooh4hrlPtJqA
jnT0HkDx+KXGozr2ROLfsZLWvkIHzYUTJaLyFxX5sygvahJ5M3r+e+F6GecD/6w/EDZ0WPTiPVeA
Df1YPK2iU91hAb/njrCxlnPtQl9GGAlOIVI35B9/8Pbj7B6ntqRKVNofVlQ7IXB0DbONMe6f0Vrw
6DM51y1WT+RbCCx2taTsL3tsqBeA1amPHiQ30zeeR+72Px4XO14o6M2gdxsuji4YPWo4wK1twHQf
beYDGAjoMFJFYP0YApulLPRONUm6f0yo0iENvizJbPiPV9cCNTO1GIhQ9Zm1h01CLdLmLaifNNXz
8IeMfRUYA/SIae/klSnzPJB0TJ87LoneIx1n7PCHhDHyFP/NbUSXBxxd5ozjUbpEqlznnbB4Bjxj
D5lab66WWKbcQL8344rN0+9QFn43sTyjb9i1O1NdAeHb1C6wt9o0x3cuPlUKJ++yTpaHSxUuJSMb
pZ+UGME8EfIBYl8KG3Zu/CroyXQh8sdT8AacZwFi44ekyNQDjUDW0+2Xc0gq66zlURIeO6udSQDK
/eb34mpYqnQu6M7D7NLAYdIrqvUQmDVQw1D0HKH7+29Nrfp8Z7Erwu0zZPzukVNYSZN2IqUG8OIr
9Xbo937bC2lRV5T+2//gYUc8e/vW5ewV3ahViOxzxnH9xf2+cwZ2lNz63yafdHjukhpI24XR9pWa
mIKsDMDdpF3GGQ5bGCMQu2z7YM96CU7Z2AOCMX9A93ngVPYEstFwOk5MlXzAoV0sGOZVDA7p5bd5
cYh0GzD2S57LarOME71PMw70ipfCMHOvXRqBxAS8GG1av9GGZSVSi3gupBI3cJnZ4lgMwhwC7Xbc
gOBciC4lOT+a4HlF73vqczxZ+9F5rvvhtisEmKE/mY3OkOgDhB7s1XQjj8BBj2yqDx0YhY7GjM4R
3Qb0HYoEL22N8oU1p02Q95A7UtRjMwLsdUWLGin6Im/pXXmZytpvd9X86Wa+RN9j1o4ZX2ZBg3LF
6yRey5D6cR9GpDeFXdfhD2BorxKJF/0HbYQvHRUnaX/Xgnftq0ZaIP+qNoFnGoUjGHHpZ+YbOdTU
oXF01vEmmjvS7ESlC3zc4TezHpgVBKG9vdN3pbeV8v08iiGKo1JagUnht/XPvXfhaI+pyKdRj/V6
6njsJ57keVzhrsJuxAfM9vcOhZ0TdOHerAtmV4QxjBYZi+jPWPmY6/Hp+LD1K0a+xloloodhPx0y
2ei2RdrJDdv+aRLrKRlKWp3cKsREvJev0SYZiN/Qu8b+gCkZOu/PXnixfCRqd6jD4tLUWSN0koh/
NT5B6kMxNKJ5dhrcflTcgBC+cDf0s9+gkzExihgUZJ2tfXpiCba7hZjTzAUI1SOcIuxnCBG9Cwpj
0fOvJtc566SJeuFY8hegyhFnu25bm122Gv1RAh6KrNYQFjtf9NwmqPQuo1ORCb7yO7OraZ9z7w5A
iq7KC+dwxwFtexAa/oirajurrnW59oAWptUr3s3KRp0qB6sMEWCh4uO47KxBPp9dkppeTe2eMzFA
3WMmMoZv0NQpAU592YNDTI/tYkUJnXArQhVWKzWvP8X9/2RiFwL9fHfhjuvJUOY0afP47RLjwJOK
BILpOG3FzMlBoaepnUU5rbnPUY6A2OjrZyn25Ebc+mC+QS1ZDQB28JuBOvM8iYK6wJ1CWzaH2iXo
iF2dDVY1q9CB4jC8KAQuH0SnfOr9cDIpXqxKRQDfdBMY3fusy9YJLpuOv9bL0PjcrIXLWOPOHRh6
dgaaw94TYLaZcxK14CVb8P0U7B8pUCIMAYQzNIHBeOzvsm8j2zdcyOfL4KOUJYT+VYGQGcVCaXIn
SNap6tG3vm+VSXo4WUAtIXcVCf1/flFNT3mB+VepZriADcOHGjyG6ySqWpplwPue2VUjKohtW4FD
80Uq3pBoBwOc1mmCm0c9g0GYAUn982mmPG2e3E6qjAiAzKkORrQOm2zqp5ahs6ksALHSCzL/zAIu
WD1oeCFmYsfVLoqPcQnjMIGrIUnvON2PmZKDQFou6Be91fBStt8TKN/QDLrwCdvuKAIewFuKwwm+
LvmsIaM+Yu6cQgX6VKWFoanSb9mk4jMUvOCOAHgw+EoC/1af5lxL9ajdSuZk2pt9vT+wkI59CWiC
hA/9rBCOm4CDa6t8sxipKvRd5R/gLhgKfq/vbrkour/7t2qHgf8wITotFdt4nFR8GHVDRd+52BhL
Cl/S7vSFwR1WoRjzP3AHUDwEkqsC5xFKqUbLk3D6MqklIYkjiPf/bpo6DRr45Ok+yQ+Ge7S7IGRd
myki0n3qnLs/fmztm5ZMWEZGxd2fqpkpR+Cx4U96FQh5FHft19Kh/xcU5pmKXq2FkketpVa+AkLF
8htuqWebEuOtPzZkENLXAxA3izYTQ9xu1tlVewnWSKwr5Ggk5YTaGJ/nmjtkQeS4lsN6w/IaGA/A
C1N3J4Ra1Abg/VVbB/pzfqF50kglkK60kfH/TRDb59nQRNGlt+rUTAXTI0fIL0tdtdzglS6hf/ba
6tHxQ2eiIVlE/zke0mc/5QvYQrGuhPdQhLfic010OY+zSYmidpkuiNnpW8+WYGAr3FsiqMJ6Npy5
MVqJG61nAyj1Z+sZbqL0OjDz4ozXz6lRmwzT6onioe5CvO5PQEXhmHNh+puI2Yjm7zjM9dVOFXXW
6FfebYpooRgjkxc9l8c/WJZmg2w45jKMydiucv9Fnv1LkZsQPu3WyJksFx/4hSXhqo3iOjj6j4Gv
/XipAYoN20FEMuSnrSWAiVIIFp4IbO1DsXrN0h+DvpjRsJW8JYdRFl5RcDfZ5ynKfMihrHiN3UjW
ogLlBI9UMm9OAgPtcUJUpryT16OyqODdRhU4pGKEbfz8u8+7biq6w+UEqbFA1mqBzsTkv1jR4hKf
yyVODWM9VaGdF3oqtgMuNj8fj1FWv8n4FiEHi8T3CrILDi4eGVQ7aLedgvnif8tzMOvtmN8A7ZcI
IhSCsSt6As9aEKrNPTwtcWsq0fJ4QF67NFdrPoViFx1clN3pgKC1OQoMmbxor/oBWkVIp20nrPVQ
WB1m9/7/AhMQwd3wTebwomvHKxTleS1hXNcf6YG3grBQ7NJCqh8iKPQdaLvt26oiNcchCYyzBIHl
FyI1oCQWE4JpRRdvR3XjFx8ef3lUTuz0gUh78dAlndDMclgxbRwECt+d+5pNuLPgko6Kj1QJATeR
Qj53BaDGI3/68Jchws8ZTIpkRgwQQEeMecbFvVtlMs89spK9NGBZaCUYXb8aW6JORaob3/pMv820
zFzPeeHgBuK0PLIqRKIXnWWzLdOPpSOKtt/jKUwI/RD39r4i92aXnQRHjkP7JS5zRKN2IXKs9ygE
4ImpjKanjTTbIjHlCoyMicz1Ya80xeYaQVvs5d5IVmguKS6Xh5dmBkts8FJsFcLVp25ijHUHkPmo
QgfQeYutLqjzAfGMgUinu2V/h/GHl9K0YhN8THqw9ryyX0zfFfqEeFeZlInbcd0xN0QPjtuTcpTd
Ehhj6dx/DfNp4XMqQVxjJEHNAjdkSYZhY89cqmOajlbuaq9NkjuKjss4bDmwTeaNSNZxiu9BePet
3VfD38iGNyWYNnX6mZRafqj4vaKzKehHIvLeMlGCAKe0e40Pbdu1QUrQ/Rws7TDsDoXlBJ2vCARa
f58V6DQfbBGWyGH1rlHJSxh1Yp1ryodYHFITZaXl+L5UspndnUbcAhU/tVcfrmqBxBKz7MfZ+5HV
LBKH3CyTP3XvYNz/IizqpzMHwJsWIAD0UHbS1yHK3eovYkY5Fk01rx3YbJj/9NCoKFuB2y1HiW8D
rRKDvjEasjhcSB1HIZDBzvwpy/w30soqYJQ3y7m7CIVUbM0sdqDiN9PSYiuIeqpNPOBjg+ZyzQXj
tZ5XbVkU/HtwTvPGYS2vhCWsRlUmrNSv50o5TMu+QdjTjEIPYFNxsiJ8eUrPoKpKgDIOLXboBwCY
s+HhukHVv6Qo8m+LwWVtAwQoo+f7LAvLST7Hxoa29Vldt4Euxhe6Ili9zK54VeKhZWQsi2H2bcPF
J2DsTI/DsKGpTNxLvuQRgFnMEZNSQZySkx9KiFQjprTMFwvOXf5nekErKHoJ00jXSSsAu1tVYWaN
wF8JP4OUB4D+qV0bNd4a+QgwvOi+6q8nHY1q2wzH+eup//w1gSHQepPRwciObxvKLoHlXhqsvxl4
zE7Z9kgkB7RdN91KhtOsG4Oc8YVm7QHBuKMBiPWSLrNBu3Z4t/v9LUBi0Ag22EdUyiiK9kmHeQbP
QFMmDvfPKa/ZucFCIjAIHhWqUQ6XKoRL2UNQP5Ylu6aXrFCvTOqLjXCdQzs5KhAaaNCSgCg8rZYy
nKm2EMbLReTb+zvPQOH91ci/NwdmuB3Ja2PQw3SOh6e8PsGx5JESMs/WNxspgSHF3I0jY/srsF9u
8TeqKMsailvqXdVJNbaBxsC6ODnjMU2LWQh+MDCReC0nDbxUOIY1IUXM5CQjh4BSkr19DI2BbIMd
fhBMtwXKRDwMlFirPflATCAHXKHbOfTbXBB5FBlAtBpC/9twt/mb/AIq+BvnXrjO7jbiEnONTCiF
Aa3Whwxz3XsgioJJg5ekLY6rZYztm+RVMSP2ED35hMp0lCr2VcFjK5wETjXeL+tpEhrvGe4zIzIn
1zsDVciWcUANkdWWUUi5Zks0TwertjEVt2UUY6yaRC/WAoiU8XQtvg3rc0NqxFTmnHQAItwZ0ER7
mxGVrUYb2SjwkcgeX6uf2gE6f0N81ZInlUUwMYXDEAgIC0XIgH5AiJBUFGA2ex2lCeZgRFPDvKQe
D/IJ764sB+WkVEHkqpjZdakoiSXFMKurKlBcRqhQ5cHgl8haRRIOEhNHpk8vNMqpbXkMrJqKEEms
3G7urQBnIPzK9JYx5nZwwO/tmVTDvhURlNYagZoNNKueQaeOvclp3Oi0Ge2XemIim1wEA3y121X8
7zLblgzdTN1dKl0O6NKWPNrXPZtCJPmRsWySEbndgFLeRVAYsa5sNiW7ZspwNhWmFP/2McmkvHk/
gaJBafK6hPBJ6QeiXXXZG006gs738UOONa/D1UKYbKb60D/zoTFfkW55F2ClEnFzgDo8gbht5Kfz
hm3feghchI//VA1Xcx2voMMrxTntKqo4IshAy9OG6HJKRuGxtbX8Hc63xI/NtkY5sRzi3GZ1VS6o
93rBJmihoH6kgE4vOKDfQKUlSRpxl5uz1ebw/qoeBGuVs3f4/WFKe7sskLVulYAF+8vNpXWVyC2s
LB2z0epzZsypywZzTXFKZwhJJYm484RZ068Dn+aAuWT4rVIDL1P6D2bELuNChUthS6SbIpVKTYyW
09gNGcBG/S+RazmQU34QadiswpMyLhQOMSlbuAnd9ZK/Wu2g2OKO8buRoWm2fFIOte/eG0zB9Jkf
5PDF+pvcRD1RLSZu8VR4gNsMYmcfpHb7aVX/Eexx/oR1WjlAv5Eq0+m9sTrzBCKfD+zL2itYMRtW
qovuFpr4aHZu8EOKrN2vm6/+h8hu/xIYSlSD9a5zHQGfKgorhCXN9W7wi5UZxD7f1OaU6eInX+Sm
9zSM4sGkgBEnlhoMDeQtpX3BE1uUh/IcFyNypLQBWxoHWKhwKBD/XdOVwNRj0hT9dbMnzzvPS2vD
/yeU9nTUMY3ud2E0BV+2X4xwlQ+ITfieoYQAZXmYmejaC6z4XTskIjzyTaU82MCuiQa5fis4VtxV
DOHS4b8eSY2X1tO7Q4BqcwFOZV9bckOO6DYlPgcFbrBG/hQbT5Ak6g8dTzmjTutJ4fjFl+gab/fN
ygR8f32e2dqnqTXG9EEC/GQRRoNcS+MNFLjemZTqvOAy58jJdQlNxSesFfIKuv4bBhOeVxq6Ah0q
Qu/06isf0g/E7sy6BrHO1NU8EQm38kT+n/rBKfy54RKEf1sqCyqX/yPLJ7u7HH2oqehHe5ZHuVbQ
uDCE/Kv2rS8DGuDLHKty7GKKzrgC3rLemHkJUVmJyN8WOB5dJ7k6e2PtHyQLY8hioRPJ1FeHmjzP
5LOWkHA7AU9hJ+iTQfRRBUljwEpB/Ojv5CqnSb0zZzCkibmjXk2aYHEN9idrZ5uHiJNPjvo+R2i+
MUUztgwM/2mo3SSvo8ZgUXLzlqq+lb7NyQkjLVpMWEB/Dkcxlyxy61NNfHimHPtqkAc6Dp89dCC+
hqxzk/nyWj+NFw/nQt6XzvWC2MGe8MMsJTbL2NlA2qwP2fiPPR8e7nHA8KUhiVT5xP4WgAjOBu1N
5nl6how3KhediQ6G3FLELKHlyUxHyS6hgf3xrD9TW7CmkTWDvIQ4FQGLTTO58UJNeRq9HveYJSHX
/8y41QzNnixPa33M+7uAo1rmj0a1S3fd0kDxmCHWEzc4q/tgedEjA2W4FhGv2oj0V8A/NOzxy65E
N+wfxonpToZcY0AvLYktamSm+CnQU/MTT+vO5Hoi8EFElgs/aaTC/6jh8f1L97dgEwSCKHsXjGye
0iiE0Ud4z2QeWFC7KqQUKl8hyy3eS2534ZBseZfbNMrW2lAodHcY+WK0fOpCAU0uiFpXwn2VYAfs
XmItofNo5D3nqLwuHdhOZ0GLdB7KE3qaF+hdCPTJsRKyMjU9uKbp91iXD7/RG2Swyu8UEkeJVIhG
wHIRlD5D/8NiBmMvCqYT+XFEPxoLHObRTGZ+UaelMYo4dIrcRMNM6oIEOd1d/nhVLck1FscbZR7G
M085f4vmJKI+Lc+6J/YzunU8fBcB179CsPejQ8YALFxbMkiUCMr9G4aMd0JmcehMX3AtXhAduVXS
I8TNlCZyxGdDrSI/r8j/bcd+k0UgUvP+VAv23fZNUPXmPKvLccA1cpWs846z6/zUHoiGpCaM6iLa
LP3MD5BbScXF4poO8LSW1RtTIk1GamZRbW4coZ7QP7u0NT9y5MC0TdBBldkYXKuYuDySuPGQSsag
MXwRHBrzqqyC4+f8gHxxDiez1vxVVF8FaCGYiTTNib5yGp2MCJvsw/VY/UkKQR76mlNlJav6XBfy
RlnTvdxt+6B0daKyeW0X55mNwITxQ6Lg1QkF7QB6EwD5obnPsRLSUYG7qnHldzVGD6l0K5Avwgni
EMIsUuaW4HKhXt4KaGj1bPq9oyNgAuy1yQXhek+FGCAuy90bmOEkT7Uv4pFK77q9tpYbjcPMYdsb
ZdFl3cuQwKk8p1jy3DGRVnmKTZJ8NfgAs/t+nMjl9YjmRSm9K4kvCTGzu5gwmPJPdsTmzQCDos7I
+cLWlMlfqHHFbL1Yvww2F0S6LEruWPeQT1yJmnJXobI9GV+1w5+FCqEA0DY7XpD5mKAUtByoFs1N
7yUInKFeTQMD1LovJ3gxnlDGFDhtonm0W9SdbnY96C7Tc6M9d3eWboj0+214TqX/w2kEkUt0HTQD
tdNtSrEh05wjjwW5wJZC/+8UIGE6J8D4wrMU8VWnx78rrU0hF4e4HofI+9TfSkoRbW2GbwV+ywCd
P/lxxlUMmMvVCUyxMN7HtdJXIjYS803GwNuFoKawc1QFfjkxElJDogFsg2WyB99XhQeFAkJd7YOK
nbrQ96RL0idcLEc0IZdqz5L4LtMKaomBHoJNLSiiQTSb8rlG+BYyYnmrSlGVnzAE9I1OpL4I3dVN
XGxUvF/YAjwaQ71p7Zvone0Lqx+/P2kFapG8+HZih+SE7wuFqvTUHVodxB9L+rb4k469XrBgP5tN
+zjCw4A8Q6fczhMwsenTIZxMJiCJUq4FmOZtLmLiB4nODbLUCqKPg9aB7ad9JoIYAhXTroo+xwIZ
L2TlbLDE5WetbVax35ZUg6sHYZJQs6zagJfybpUpOfDbAkADPJQpldm8C6/1+ymh66st18EafEat
wQ/rni68qJ4Pl+ewMxxVuCaQbMCYZvG1JuaHWsCpHfFQknR+yi6hCbLAan6jssVS6rGx5aodxLkf
r21X3nOfpyctY//0g7u9j5zpDRdwGSZMTvWLGcnVHDwDy/wvKiSRWwXb94bJcScGPuZIXYzoL/l7
aSQ0SItv/8zs2tOtoWPCnqrpsQ6DO+m6rIspj7SmIv9zQxJUD+K1368B2NdKZb9Ty3vTWdFp1IeD
tj8HGTZlRwLvb+hcErCjVQUMe9AItovwkaJh6QswBlscKE4Ba58yh6N6hvi74zk0MRpfsd0bNZtY
M+qMkOFDCPNxWGeV8FHXmyEIlf9dgOJ40WQvFm2dUnag0ah+rDgBBldLs1DevUuyYSGYkWLhIQ3k
fIwXx+J50jmmwwdg6v+jS8C8A8KRyR86vm9ttuBpyGrm+/aI2bqTIErK4s7FJANdQSWywCPHZdhv
JAT6SAA9srTi9nmfo6bt7WPgsn+WPcLYt8OCLKyFokHklnjia97fcl7zhVQtx2xVUp6uJcuuimf2
F7ujVqA8yLltibSplWaXGQWkuETRo+eGenl36EHqNMHT5q5AY8a+dBu+o+tvD2O/gxxjoH/1XndF
0Ia8p0XjeSMYDHQpjpj9VY5aSPeN0VprexsuulfCNu5NiEfhE5A11TRZQ4drwoKSW+p3IkGkIqF0
fT398s6kDQ7VBDTya0mBLfD8qv2/c1gUUOzfGijwST2XsoZcJdZ59PioFYKyya9yDLM68qCjvL77
xWA98+nbl8EKmKZ1jnj2dk4PtyZXSImY/ymv1DVrgyUD/OWPdmcTTEuBKKmRM1knJb+7uos8NLt8
QXVMNxlLWQt7vO0eORlMkKMOFgUGfWP5tbAeLnu94ajMpd3iz/KNKMWvTIHwP67iKMvBXs4/7SJt
AgfdpW00Hahs8IN2/fx2a7ZaTz0ipe9k75Lyd2RtnDAEA0rH9YmW6UO/A1UOQ+G+7D7vr+u3u612
7c3hPC8MnWxlVcB9FVGdOV5lfl2Hf5p/CgMtvUSIn7jJzIm6lwv0ywjmNUXWBzI20YxVh8LzZcEb
xzJ99BWa4RWaI/8Zow6ABzV/U3avtZW0MjRvogs0ht1iEiEL/ONAJ5Y1Yox47bXtea9PcNbHLAAL
2pEVwIwldYHzxV3bNVaX2UFwlfK/eyVvj4Qqd9JUHfEYyV8iPYBoe0HGq8jDHxOkt7qsLA6nqemt
rZMW44HUGBHDygZYUkbOpy31YwCN56liHE8tI8xbVACakev+NNUHHS7SKQRjnFZrr8ej67S2GzJn
rfykzVEOLLP9H+kcYvNM6kkEIU5xz5duL4INhuqEvklZ2GC0LQhu7U7rSxeFkRfGJTnVzEEDqfsF
dzcTDUKFVHyXziOuTSbx+lRCkg7un+jFg0Krt9PmGhqSZ+rCxglCkVrPbRK06QECAgIX57qHAyhA
AAeNQdUWnH5eGtsaJV4DZNGxWqu5faZuSorEOPdt8uiHvpDJtiMgy1BP7pX01BNvkPnCe8M3Mv4h
/I5eLW9mlJdDzUaouqJYymL+BsPe4h6sDm/3iID3So+RNJvqZ44gpFh97ms5vohD19JTyLocft9s
3z0Hcg1tBZzBzb0kjdh9ZKix1R/kM5F07V5pgBdoOl8VFXcVen23IkgoVp1xkkXZHDyeRuy+uQy+
tZbHYGYeVoijjdqnAodT6xv/Q9iI42eY0Gnv7mpc2eQogZYzDirwrtYz5fhRU5fV7b+JooE7mZKx
VgYFwD7zVMNH9lmmakdiPg43B33YB38b6otLoMKtWV9hRnrexnL5cKe8KkrZTXnv90M7X2F0mROx
v3xpZ6U89EL21pB17kSzUW6ym//PcXqBzC3Yz2PIe+iCbI0vfvXjBAZEXJC00qE+Zcath+oHQ2dn
A/VITixpipXGRT3hdNXj/utBwJ8uJ7LLFF810y+Ep3nPTslDBxf0sH5wgvziLkYlrX1ffO51/o+9
TWfvP+Imq8wTZL1Wa7kNczdivg6FkdXajhPETEJF2y7KBoSd5eqUel7E/jrmyBf5L75t7xi2RATK
d0+ZBs+hlPCBkmtxgvL/NWJKQm0xi8AVCR1EefAhPeVk0ELo1n0cYz5OhhNhjr3sxmPADDq6DriZ
QciBKW2fO0AhUuVAZ+iqfH35tyDrs0cMGFhYvMDebB0lq2cfRRGmpZDnrdVv6tMRYc56PraG+7Wl
j1eQ5ilf9mguX76b52mcP9/aaQbYPWXu2FfyD4H70g+EIYXo5zhXbs1+zafg57JH6vrgH0bQwFcH
ea0VIODg+tQmYTpCFAijifeJrIAdmmlEmUnBmUbUN9X2t2Ts2DgIhcIeTI3cS8CAGkSWbpAvk5gi
XF+Ld2+odOmiC+u3vAcWTk/6NefW2FPLJlR9rtAKmZy+ru9gjgmmMh9JCez9Icw1vytOn7oO7MzF
Vx0Mo2uxTxAVIlF4sXt++weRdEBtEwqkAke8jXJ/udsvtTe/ricET0V+pF/dfpT361UmF/Qn/ZqY
650VT83GeTJThzxpYpjHirVvfxBJpQDW2EsAdrhFdu6AmBq6yqvl8EvGlKguXlxV66XAfMZaAvsU
gMWPjWia2Li6EcBDlBFDUXRdeLym3duHkYHY0WA4gtwdxVofZIlTfZ2nft0q0Icqb78QUKoa8fyO
2SYxhiQjKukIB7bOXjKepE8blJBA+HqRT1kRd8hEt3hGW2syBOWcZPJRg0ovJmIRp5xOEw9yGCi8
j0k4uhgnKAjiPtxHmXf/ePLmdvMBMdJjBjdRJM60/oenzfEbOPfhiNwVtVYLgUuJRXvRVPYQ4w2h
LIN6HKOzQXOlYAFSrozxRcECuMRI/pUnIoHRL/BFNIEGW73Ipx0ap4eNhRBbXAEwoo5Fxf+Nz9WW
hZee5wZtJTjpiKitPbFV/uWyOVBLoclbtFJEK0G/ZvvKVwmmFsVHHD8eCgwEJHpsomtcx8XBfBwB
6zBhoSj04MBVBg+fwjXvTrlHCJmY4CRBPZ4kgEiN5+H3ocU57iOVL/AlEE7ApSZkFhDfH4x0MAE3
Gr7F7dbWBybkpzmWxdkRrB6cViFjmIy6yB9UbFRbBQVzygtUiJmG4rKoVJjyPH+AefYQ8A7x0oe4
clHrAnZaeFQdxgsB5rB0+sF/E9u1wNejeF1lhJjGeSzA7k/SBw8I0saGtdDb5RacXzVt7hmZGg36
RrRYK07neVYqD0eqEmGhUJQEcIiqJF1TyS+VIZrpxjqfhHSW1JZxROLjzOgntznM/puIYVOaX/Hi
YyaTSqhggrBRPHeOqmJiiEpZiA5r1QUytFt8oXgFgmrKKxX77RAqwMuMlx7Bqg4kpv9b9Ax2IVY4
bN9ffdEoIolKSioVFmiPccKjUe+RBnfY+4lIzQJmLaG4uw2tD3isTpPSekTtQ79K01z9zlVRhabn
jmkuueEgIKPmZLwJnNv44wfrk1dwjPNK0M8lVKbi8aBwLVL8IN/PCxASl9TsFBVQ8yccWLW40abS
yWIO2MrWwcRBJNfzszWJYoHggRD70Wp8qdEQvb3Kq+uzB0mJu//U15dmSXZ20AWjyV2s6kSNWKw8
UBTbOqu4SqHFY8mMbOVFKEV7J9M2S/U0spUfeiG5QUddA6nBY5k2NR5k29fJNLELZ8bz3/3MlrCS
XJklz2sl9fs1u+oyyVUzWwovL42vr+L3HpqTC1OKTrgy1JykxQQQqsyeLrezcauP+frSoVn3gnkl
HovPE8WUSXlErimr0xhy6/AJHcmDlpyPc8Us1Hwkb4qdhcHUBMMPcOozsFrfXB86B7ZMA+eQfbLg
d1GRBrGknd5SimjulU8I5YybJ8C/vOhPum5p4MQMs3pHCh3/c7WMj9k4iynVsSBXtUW5kEueDC1U
++er5UR75uJfNR4xH6eJAhT3dnaNWZTy3J9IA/Oi/h19fTyGjv+pn52fz2Wy1RgQLw1G38FkpNR5
OcJgw0L96foIA3lkOYmCcxxJT50m+H7KeZeP9hQ1GBRXIivW91rBX4fryHv1wWp2F7rBKhJkg793
Su0s++j7zd0aNLfzgTxP0g4EEZzZEKS0XPsF/vx8nBPyQtSUK5XPEA2I5SwkC6DzfI5LT4vGNJ4x
59B9dtvDpky02yIbm/5AoxezpVV0FUhhrRiG/uyYArbzZ9SfyCbB923cgzglZrqdmdWrohdtsLWa
UPvsPwXoq+f17s3DHv4fxzIVXpKZQnE0GiwHRnYroFdnfXitBz8Yl+lfOwq2Dg1KAgAEB3H9TaHQ
Xa0RarLBhkVviI4CCtkJBMrOkWJBkYT60yt1LdWcxgXDk80P9DiKbn3STSZJ0fpfWCZPtVuIlkaL
PjAGc0eh9wG2JGK7PXjfBgZWZjIXu35nuhXtStyRTYdvgBVoltlaW2V6glVssLY5D8cBvhwvPd3Q
6q7xl8rIUAF3fQ8fqVZMZky3i+j6fs7hWh/Xi0P2oMqFLXG+YnKXhgK7f1RzRdVZIbIMSDuJj4i+
/ZJyBGktOeevJzgJe3afSm4Cpr/DSBV1VitBs4yEGO2NGycj/XlQ3IdCkNyR49BiO3FiV+Zf1Ezd
iwRzhny3CXrRXraljXYuOFMGdp1udVn0S9IORwEIALBCaBH4F1KZIP3a4l8EotU89pCZP9+xaZZK
AFYCM8IiURPNzNzTdGldFS0tcxvcbL+7dvDW5A1VhEA7zCd4chl3mgyHTdTNgWjZwmkBO6ols+DE
XgsFf1Rcvg8alAnhSZbUY5VElbfhXjmVgA1eMcdAKGmpuzlVrFB0f1g5woTtcoXeZyMCaSyJkdfV
CIBaYt99QDb+xsz/VG6J92DnurKjMza3Y+lxO6mQqRl/Kmjd/C4Ar4SWUlC8SGH33nN1xmnkI/xA
LSFdOnH+ohNpE45e+/4/Sggk/eZeyi73M+sOopW2VmUSPxM5O2h6VFPhGmM0Nm6bynDbSpRCmt5b
fbxHCmSV96j7dnN3cgHA1DZCF811BIOUZxx1sfPYzbcFCFtcG6AJUrE2M4Wobv4sRRgzlSnYnQiG
ew565kHVf2s2gXtmbhFg/8/hf9MFkgF8sTKOlfm9lmo0E6xx2Fq4kuHUwLi63+5zfjs/6nt1JuiQ
a7AHgC8xAXsPmaHXIiCL/AGiGsg/OOfjrn5K9gEZhwTGHYebA29/O2ltphT+fgsIdo8/lV+rJmB0
CBxmMTUVZHgLmRSkhWhzIu/hpgwCFnmRZk4/HCme11FWBveq1/+gMpPlqYXgK2ovnRsAgU4ug8zf
4o9pPpIOt2LXZ7Ej2f35URD57hzLsR4a874cVr+lDoemV+n6tZxUcXQytzkWQmC3g6M6Yioc9UNC
ualpsq+EhdpeTRPpAC07cVqg3T/z0cokOvwOVq3r2xOt7qReL0cfT/ub+aaUmdWWmEZf6DrWC9Fg
K41w6pg7rAeYxPCemYKa5wKJYe6YCXV7XKNiPmEg2i3R/ScOCvljacRVLxGzMHWGv9uWdQNxFp3w
2Q5TkBcIfvpCJ32HlzoTcn1zngai0R8rPRxWTp+3v7FkKKjJ7yJdjRktEHVBHKgt1JKoXVilPFi7
gtPg58X1Vf0ZFoJpoVbyI/8sb08RSz7aPQplnmRzhW6Cm8Jg4WBxDjWvBZ93X368gfde9ahp1k0c
i0CtBPnlCuptL5dZnJdbMuJWbLaGSsK6EKPAiAIwSDqishg4kuC1u8x6sFBGIcBdP5ROT12mwijw
mDCOWv4gYXn2BkNN8UJ9NwSt/3DrGgpMCFagz4Neu+5frErNr9gHCH9RqkA2gRt5wseMiGDvK3Fe
a9Nq1Ie40XouDFgMo23b8VvLMtPHVdWlCOFY4sPk1mPdwY5oGVMng47XRpOW1u6NZV+6HKMp8K0h
FH4hjMwIDlYegw1cFgqZHF33UeI9n931AEjpFkxp9HRA583uebIaJYj9I3stG+bWweNyRs4EF0C/
npW+JHOppUxXrK4U19tRG5icl9+MjLyfkrvnUKUE6fdE6DXiTz72PMKJJUEwlqlWXbElY2m7AEdO
TatxX7fnsZUV2728ghAFaxEP0nVJhgma5Z6rzV6kWZRhaQRxRr99XfgH6r6TN+r1QpxVLV98kLti
v/NCDQhllAGoXMGN+qStl8qTznTgkPGGAVMCdEQRvAuOOOQUAqhP1+Xwdxm4jzZvbhp0FALHSNKO
rdYU63JBjFfSQaTC2hhc2w9ONpkU0BgqEuWmRl7NMKdHuXNitM+A7kQdgik8eMYoD1gSh/tLWZIh
az5GbnkxDCVU4nUKLGjTZpUiL2K0rtfoQINspEueDLS1ILWpqUa+coiqzoMbwpcJL/ZrG75TvgAV
lQ0BpZDKDmyVjWH4C7SsnIQhDniG85G9Sb+qO75SCRBvjXeHe2ZIiPlwQyIuCJFDPfDK49MoFVKL
37pp8lI2tsczQE3BRcujvqOvF6CThremfn6Yd9VV7ybhaBMBpSwUnPN77UIqdzw1I3Qdd8kU1RH8
CvdzAFnca4eLW5qSoR6u4Pe0AvqDEXEe7XpHaU4oPTe1QH2GVpz/LOys6EjSppgq31bPCOZHEqz7
FXB5hs/xbjEAfXyjbTT7wyic4nU0kfjd7LDf7rIjVba4YS7zl0WRNuSPmNd89Kysf9DF4JVuFNGm
/RyNqeSDOaHMiOasxqa7Ipji6WD4HaYnESelnol5HPpYiT4H8GrpfrTWHdHY30wF9a4SwkhSgER+
o7ToyTySiQzhes1jpi3XX+FIGV4EC6Dr3XwclypmjlGgvOKjqYlHRj0UsvXHQs6zLtJyx44VHwB4
rSdH63agrfeml+/fGaEgx65QmuT7ireNRc1UuOMC8Y8HY5CDsw7z1QzrzbSNFolPJvzp0AzuC9dD
dVBl2FT3b5G4HOgoTAl1cudvVwCvaSi62VX9Mf+go12fL3i5BptoMLuvGCDXxBha3oyGyZ6mUXAj
yy1oRbL14J7rZJFW/sqJQuBl7gMPpUjHBVIQIHawe7UaS2gxz+W/cZs+a+AOGIf10+POlTK68iBq
BHQZW4tYfdvTXIDavJQlQm8g720K6YKOfmodmYp8lDYUC3UwzxOYtYtBQQ59JJzmiNtEIJTc4L8S
IeTIxbm9VUh2nKUSo+Xc+wi4ppQkRACmNKmBLyQSVp/58VWGyWxAoueXXWp273fOO4MUDPDoqPGh
VfZjcOfhXv/W7qNy5oDMYQqT6ksG4V7OcgBG+n+2k/BJ0WOIB2b0Ck8UcnnZDkXITsIgXUjyBFwX
bp2vfzws4Sy/8LiVoAYwfGgPihV5n45VadZrKt++Pn1tACcGo68vw42tvsjVZsoOWNQ8tMvdiZTu
EWdz17fl6ozPQHCMETQymyZayjJgI/bVZIojCh9xGbr4SyjejeByEFj8oAfbxVLyqsySEohB4qnD
Nf0YUy3o3oh1dvGOOql9y0ZDly6j+n8VDNQTePOZe0fWCK4vIIBQz5nQYhd4NmyXFuQW8s90sSyt
2b02sf8L/cajdi1Xoy3PaLoDoXsgjoUHD8VS4r2HAeHASat1Zq1nZGDs1oEousHbD3zQa88bva4y
KV8qLQRqAbz6slodTog36vy/pyMCEEM0AZQUipg3pufTFS7WV9YSGXxRDNDpt2g/CfJf/S3Tyntu
wi1fSyK6oXTnAxBcf7UU0/Mw3L3407qs0fuT1eqM3k6ooG4vBjwfszUokcB3KQF5ItN+YcQM98dz
8sT+9aFRj25XdpsbgAUtx/qByaL53L+SG08ETYy4pVkTONxJKqfeJ72Nn6/JTekju9imMo2R44nB
DZfFCEUXQRYZXs/3la3PQVhm2e8ZhrbR+5xx1602dpGzBIi9FBE+KlzV5QYZHbTaepsnzRUuR0m1
YIaGu+SuMBBnTLBWF96q6y2UNFxCUHI8koC3mFq0vXZDS/DgOcyIkQ7hvMmo0kJOKG2GgZcKczhX
3DK2jZnz7SK+v5JjAXNzkQhTbDR6OXuIeMnyQb2BJb5I+PpqywnrzoVubJKDEFQ3NRhwgwiCAom0
/NaMqrPpHyL49L774I+Y/+c+P/J1fmhcd9E4HQ4HgXG+8jK9vfB+a9jbp2ilEOviAme1jsnXVUsI
l+Udqxo4wzco23mxdXHXTYcaQnA5lkSTeqBTcvPR8FhCKg3VYbWqVqSuU8V1kU2n76XqLGI6soLV
NctSuJZw23frYgCwPvxGH4R9tVqnJsOa6e1dv++5JQasNB5f+QE1NyGr1q7G1MP9S/VQP0QvVC6c
5J7/DUDQUNUQQPMstd6ld2mluFkWw+omc4XY+3V1L8THyRxlCdRBN9dNbBPNY69Agi4bDTI+PfOv
lijf5q01zl0OnktF+3zWqUhTh/F6fbJsDXgEUxshA/nKwsU1S+SnNkV583vTk10qaAaAtvycRgcw
wG9RnTju+s3rpFhIlLJ3/BcvMidRZpW1Y9Jva9goCX1Z1IDL5EwEIVM2TdklHnUOv+aD8VTZHL7e
1q8OegJiqjCk09RgxJSG1snSg9x/B8cdlcJXE0YpagUSz+EalZKZXcfVZ1x9WwHs9oFjEVLvI/o7
uzT9caVLAfcemv8iIY3aB7pV6SugezanorsZJiFMdJphkndUnTFVjR2IBNqFgcjyB2uOwOvzHqRm
8cSDYqW0OewXU/X5PM7D2fG7y6/+r9vwHFL2eTt4FOd8ojpWWlv3W5spfS3GZh3CkE8Z6jkSEbo0
oo4e1JL4fc6doulqbldk6Mh/rQukIevKImmnyJmNoG9A65ZHt03UmrHJdNRl+yE3sivayoZUZfX/
FKK3Gv475WJntXIRSFO3O13NxM/nMeI+I3KfshXttz+NX1eFhEectyUSeJlo5ZydLJUI9nByMx9e
GqLGcQoappZ++VUMo+b9SmfMoCdxqLPBfrs0VmL3+JHNUkgNO9WxB1jmAW+9JMr+ReelPXY3ojc1
h+7Mcb6Xu7Pbd7tNi5k51R4KLpbUp8dcRGkuDoA/mVYjg8v0tJSBp5cgikwuF9WR8wi/ypxciqAm
a6otT8RFo4XfNCouiyuQ8ZcLtYvAc3K/uFg0gVcT2tNG+NfOOw2802vqbz4THhEVEFgMrFJggXTk
16mQcqOZH8JYSnGuAVbFXeP7GxmWvQk6J4hALa35Tfrk4BL0zNMxwiHWW5+SrKjelF3WqEyVirOj
7ovFRJl8xahr4egMr14VRYY0Rt6qYuFLeA+G4O0qK51UEpcfMHqbSza4zjduGwSefkjvU62GmH+e
OPQD5CcMTksTOyOJ11Qni9PXCgM/Cchf9+pKLyMWgW2GRKkthTpG0XFFAlCeM5wBPCgkfVZeAxXz
L8B4aryXZSeHzdRuU13uvyatQGpMimDsSLZUwRJMgaFMEIy8mMBTMoKhBiQDCVaOXdnuyqktdK5P
+c6jtSjQTojKF6dwKw1rNI3pdb1ZogB1cl3TLZDHVsvQkKGw5k7xF7RlZzeUrG3ViEXjXmn1iBoA
ryR59Q4gpjIygW6glgq89jAF3b3fwEDqXzqVPfc6lqTWhIBvXO2PnXMCgKh07lPFL+4MwZRByEOC
DVHmNKXikU6Ztxfp9/ZDua1E4cnZ8FIqyM8cOWvi2Bf4sjkbEMvoTPo+fLtepplv0oSSJsbvu8sp
eYUvyWkcPwnhB3hqj98P6qFYduNG/2hCjy8VU2cYg3972WmjEyridnYaJ5ghKfSoq4VhERuQcc/6
LOsr8YzZoFY6+7msP9HlPhTg2PC/rQFLKmYeR8Paqy/nMYn31lQtpuuVp+DoDD31Y5KXmxStbFre
pij2azwVUa4pnt15jr4i0e7pUahe2098Uhv77foCew6XzjhgSgLmmPX0fokdhfJbjqabfk0Qgc4e
Wk4cgeWwC8elu5dF75TiBkh7vTD7JTHQzh5veWUKJRW0roereFsXFDABT+uzeDgywTLSjp3LxVKq
YU53m4zsm5+Z+M3oB3M96hXqKaTkmpE8oQmBfp/1xt+QrzNUhPc31Lc4kGOy3QTUrErz8S6VBcFu
RTO06Fs/yuh00l6ABJm23ByQKx8ANEUPYQw3MES07b4F8EaGRCG2r1gtCwcDv2nyRcSaUkx5uWBj
USl1mar5Np6/6C0u/Pc9pA5WKRYU/KUHdwtJ6NV4cATXCYuOus3jCjo940iAcqlSbe5O21/fC4lj
SC+9o6CmeGc75WaNx48Z7xc7PoddDuOAt2McY5tOGjZ9PI2mzFtUWHUOWcAwz4Ta5nVgrmdMz+0C
e3MjsAUXScvkU/EsaPQmthUZjhyxd5qoAiKhKJiwCKgxC85xU56LnuNaiXBj1ub/zrlHkNmXcfhR
Px3SoNKxc99mbCv4cKfhpHDLcGRfhfN39olkfDLntXUrbPMOH9EsROdpzLtnQJ7pn0sn+46MEcXs
n1jqn+ppucSpHF5Ag6UJrWd90XG+l7GSfUuYLFVCKiIK/J6xrVW7oRrkLzkTJGeGjqv1Y/hU3R8O
Wzxw2d9eXAO3iDEG3nenZAK9oMjeO96Mbqs+lHzqna14AOkUbxYOzEFahGP6qC3nokG8v0mXKEUQ
//kKbE9prLSdSD9RyBAjfLcYRUD8J4o34fLFvalgV0VANrQ5mWDOcMaObjp1vLOvrJMrblKbP2Hp
K+baFqxDXODQYtPMEUZMZaE7AzqGDjbw3ugKpvBRGcRUqTRZB4Y4SZTsUIpFBqnvpDABpyzzq2Mk
sWEkPJZ4fleFvCEmyQx5UpQdqK/4FTyMT5VkaBiYP3oCPXiJlCCwOctObtC1Vvo/a/lkeY3qpfzT
RpXDvY1GDEWx3QP1kPB6s/DvO2gc0RQ8tqa3bL67Bh7/wYT6yiPa0QlH4/s/IQjq1MVl9xlluKUB
G06FSswwceUtgduz9aTh7kOaqWr4he/p4y8X7JcA/XTtdZeijPbRdZz8v/9bGv2oedMYRM+tbAMF
aiGR0lL8HD9hw07WSwW1ukZQkwhO7SPaHK6iGG2RFsMPBwFMFDdONTbCyN8FNYUsV3Xwid3tsmSv
5i+zUsAInd6YpyqMV0HpO+QV+UZwfNILnni0jzMvqA9IrsGXqX6N8XELQKQbs9apV6J9Qj0c0xAu
Vr8efj96DDB0Uwa7gf34yGqC64DOXPC9IIAoZFrnl9QnWh9oIx0iGHEWY+rHzyHUvfw0+ZiFn03C
ZG8CVrRx1A76JPj7Ctvg+aZp17LRLMpDzTpRQiD8rbZtj4HhXazLJ1uSTQlh6YTl83A4SWX2fWIm
hQ7Q7TDSK3WdeIkFsuyQ/NH56anlTMsI5TRPFuak3SNhdr4mGilBpN/RGQlp5Hv/PE4cuK91XwQZ
79KXR2xjT7oSu+4bqxfhJU5YBy6g7rsr6VwTkTyE3ILO3+6yehQwKVaAthUKR0cjsJFa2r4cqqSc
sUA91abkq4tDgvKgS+24uavU+RE5dp5fkszkFQUR5OJorgPwansBPL+QI5vNf7J8Ca/Ih3fK/kmA
6JDlWjaH5db5nsBPjsR+zV5EUqGrpSN9SV11S5tJgfNlkrnwSbfa4fPDVQDFx/voA5zSpA+2Mukm
Xxd5mHxW8Xa3gDhScXsVVJ0d71UxUDHop1V+agE89GsrIj617z9k/sJWwaakUcPZWL4MfrqRjlMw
IITExw4Za3mrpH1pqF9vNaF8ft/+JS+1g8XQcSPnvVHxrQ2UxF7ASfplLmb9Sn5c8/+Ptv1qA/Yz
Q95t1jK6PyQ597tFfF1g27dGPME9nHnLlmsnAuF3ic92RKywMbIUUs/6kSHeXdF3TiR1/4lYRT7n
y9nfVbT+3iL0UY3W84YCQ0rOO29e4SYGjBt4Bv/FOYKArXLPUpGA2WRxlpPIbJ7inw6rYhHAq41X
qu9qMS1Uu0SaHeflLyJkfYTsfroOuKQRyaRypx9GYATXUW6EU/I43BGX9FmfX8HqfPlfee34BTko
s4brSMHQV0fZ7v7hIC6va5+1jMvdFutK5qzawHyaVQVyD+gQXng5zUnkj358XoShqD6Gj1tXDKV6
uO3u+FEFbrM116BoZ4KEPCTqeH7a64UxIAPkuQv8z3t+PaFlO+4k+L+iaa4yCj//3mPSb8M6EGTZ
s+6fBM6xEoe5hSUOK2SJq5qxwjyQP+wF8p8s3/z7IDDaXeiI7b2GVeUwNfjgmGTY1Nnuxk9mIquO
c7ZEYo4tHAQUlyA7EAPWWmb3UASbdoz8JdE/7cnHRZeuw+rV9olgHVL8mjzn+cCdSJikUtv+30mj
fO/pR49PxEwyoI83SCragKwAJyLTbAZTwgSE+l9qqL+FoGMwP0GazZZqUTENXFF6JWc05D1ly8U8
B4uiwPrBlAHA6mJ/igt101ZCE/24kjNdSeLLlwJ2iCNUmdNL9Wmu2Z3uXBOg5KcYn9YzI+IVIjIr
5GpxsBddd7tPD8cXALFK0KK4dOqdovH+1VXZFnNfvlAOXKvRox9Oby5R/Pm3AEL6eBK1/GaTHLkj
fHGXItQP+3KuNmg+nWHZ+/PZnlUXyE3drvKeq3he9gplHZgoBHk7B4nT7NluhbMLCFvoLvvPMGFZ
CCBlLWOyX5tHrd9uTW+Nu+NqikN0t4gK68wKPNXMa3EClu1nBwVGgM9NTz7uoOqGTYKyAlQYtAhH
yMPSRxHwJshu+Ov7Umos+uZcInulnFGhjiuAibzt7Qx8mOZgr8yTDaY42XcspoxA1TiJ1C3warrQ
VwCYh/pi6nCuiRIWeB7Zx3PpjBoP6VboyQ6kX5Lx598nOsgnMGxrdZtwBhnO/7vinNQnpW/seYmO
fIpAnoU28UC7nQsumcfBxJP3kv1ZQLs+kzrq9iS4BqCgPpG3aDL40sbzyn/Fg2+LK1HE5vPo8UUI
oBCKD6XlXWO3OaVoyYDnYGzOavtn0fcTzDgwmilzApuSWDByIaz5ZuUKWh+HQLyCQfjcVs3AwJDF
pbB722fPTQ+ZBZfy9HD5SuiwBLS6qmonHM+5CIw5KdLQjUJIEBCmwtioE5r4PmCRaLTXZWjf5rA/
sCvd06jBH4CQtZwIoIe0pnRa2Iqne6cKjVfPb2BkQptzvdrQQOW+TSKH57QLdK8LkiNZlMjatk2g
xZxal6G4HJyO3teuDNbOVJe34jhAudZhiTQRdB49w5BaelJgCmpSUZm3GU+Ziypc9wJ4XnA88LLT
KSStKhdo9DpXggrtlPvKxPv9rsj4VuGjWGKwB9a+Ti55jaH66NBnngc16+eD6mOns+i+OYfMKi0G
tn7BSFcYKIGK0Ua8QPX/caG/Q2kFvrud011X7oFeYurNRyhzEV35o8gAe/PzldEFu1KX8cQ3FXwb
HaG5BXkjv4blgdB8Fiv0J14xK36V4waR6pAF2pLfGdfylvaHxc5r0q/2ScCfegkqYgh4lu2TzGwE
YBxj7kYTXKQ6hRanCjBB9ow379w+j0NZVrKcccirM5MW9gNf1G//Qvb+Gh+5WVnikwv1AiMkJ5jE
l2+nOIYEqGjK9lZc2XIGGJWIG2Jxy2NqZWKNRpvZpMSDTMvkz4M7KeY6nVpMaE+YcfIueVL6P/DI
UI1MUmDxthTBOLg0byr0P84y+kPPvF+8swOsTzqYqEqjVGlRCTTdN5iMFvHyLt/0UOJI+yw6f67f
bT+WiAW7neh2EUVQ/YyQE4cLBjpQVpm5z4D/8LgQCTMzJDWW12OkJV1HWY8E75vynG4+LfaTRtPs
Nun7fXhjBjKbQ/4POA1HWWYbfPOQ635lKKDw/T/SkjY9DUeJcSo3RVFXB68y05wyxrMQiBbgzNvQ
BKhl6SC14tPjy6/5awiyg4r1wSmsWop7Gk13LA4+Occ4Lh8QHRYWsUsHEkL04XxJx1lz9ug1MkbH
CYAcOLtbEO0EPArcxLZRdCjesmyGCQR4KjelouKeHU1+/cardkaDaeWVYdqs5DRXuMK5L0Qs+5cY
CwoLO7K3l/ZpC+PLans60N+L7IgN77x+cjAN0RIJJU2MpKkYqZdGtlJwFYc1PlH/cG/4VutjC4cH
KbBxStLsztVeqmO2E/OwOYnU3U8bLa7evPiVYPVYxfw59yNWSZCgDPPbC9FApW6goH9YtP+e8eXk
Za2mPLADuga0ydbfZJg4ip1KfE7uRX2eX6LjpMlEXAZSsToE4r8/GO1tiFldcWBgoTBMroY5QqqS
NZ0KJ1kqq40FVKqUoh0LVN9yemVizj8LdESeBDaPjfMegPNLvLYopTOaadqB20XZOIj7ioI4K1tt
XTe6dUEjtyQxD6Vxq2H/RO5f4NNF3j7e3+563qBMqZomBDn5F97JG8ePfponRBt+M2jYhmsZc3Jj
9xv/IfSa8P47xAQAPhKvwNaPqC3wsj9gW3J2OE6PyN0Z78fJRLI34Mwp/oCMyOGKDNy22/7eqpst
b8c9c+cdGYHNwNHMBAh2zhtDCKYx4Uqs6iNoAIY7zDjoZHTUZVS3OIVeSV0CyWThwG/03cS0EKPZ
47UzIrhG6AW65smVcx9NejW9cjH+Vom9JZ+MB57kGx7Z20opaxOXrkh0XYHKnWGBqg7/fa0r9iNG
yusREKv5g2CcBudgKsE83iNp3lsWB9gNQ92ElANyi1damps5fglaAVmgF0KS5iMlssadGoj8jcb4
B8iih+srzHNJyDPQMrplGNDyZE1SnMmeGY1SIz0bgIChtEFxUfD0MMXYXeLDI8Tz8keYmoTFPr95
1YhEVc7QP63Z/4zyF42SB5omavFf2kITLmixz1tTpOavJ7gOy5m2KEmMIavFsqt6pBmYoM+ffHAY
j3fi9oPsTn15ih6GUgHcSfjZ/QYXnnbYMGduhopi9dNgEGsaUaR2d1JKspOpZB7HDnft7UP/3Q4Z
exAMgdAS+MVX5xMS50apogHbwxC2bJHqw4QT83r6KetsHOiybfbuoDqvtxXka7dJcMo+2CsvV5HV
1rpJIryhDWRH3o524RYXFvMbrK25KGSXDl3utp0wwPFOvMaVBnts8szaDvBpg5ac3KERfwPqzzqn
29j3DzLeTyz9Q4U3vIXbZ+HBTqK1dZDoG3SxgQz0uMJYuCKfLNvIp8DEap0wfSA6C0P3KYr8GeT2
OWQMeIz+S94rCC3uST9h4OqgR+gZlD6Njt2KAfPfn7uMp4wAXAcVXWK/4a1Vdtr9qaOHCRnlztyq
oUEh9H14UZyBXGRq/6IVzxVTXkeAHVqN2mNdjNHHHFEzXOL0a6Hwl/PGGgq4xQ62wjBEaEAVSwk1
hqpwcJsGsP03zT15TaVNQ6MwFi9DG2TCUmbE/5m61IL72xUrj6aQwDCjslkLCZ+LBWWDbPtUb3Ni
Nr7abRbOCOG3w2cOCHLZ/RFP4EMpbgYD5/q5X9sIss7UhVcsLrtIvmM5zSi/hZC6f/LHOUc/Le4J
TTfW5jVR6clfziHvLed3H6xVpqnHana7IIkMDE/FqXPZjetEzKvkF55VT4CT6mnJyfH1fl0h7v34
qiN6+tnM5D2ZhMLA7mrmHMqzjaagTNxCk1oYVibDdZA86tu4HQO9u9S+/SOjjnb6xG5n5A6ljyUP
fEZzYiCU1rwFC1PruHXeW9a1WlMG9/2QZCuMUQzPDaSAK5pCHv68kex4epGi6a3m7k1QmDKpXfsx
+a1PVF8v33moFp0jCVZwWubi7xwW4riLaUmRNJf/QcFsBKzUyNFWksMkTt/6Nk7gnVFL7BB7C8M5
rCVwexIh26cDJ6aqWCNZ98azT1L8x09dbejEzWixhO+BMwHLHLKKhRwNOQtqvfUf8yc0CcneUO2i
LgGaW6h6VqYIRgzWatSz2NHa3wSENZ3YFCE/ADb8oMyLqPX37RSZP/RRwLASn/5RGiRLUBdNkipq
SG7SqgL1H0kKq/qZZap1OMkp4c7S6GOLcSWglae9ygoygqEcXt0ZItWafgR/fjUJb1SaMMPOX3bO
hj6kMC8q5wyA9X6h7dBZ1g+ym3eeo73w2kneg05CVTqQ3UMwm2RpJijRj1V3d+HU1iyFU21EXlxE
gUjIW3JXWOUEvpZSbeSxnX5uzD5efBG+oZShBSOFGex3nuLBpV7B2X4nfD3tlyH0/7YiqteqvTnP
VWtgrthZ9o7KBmMVu1x/cN0m7Ou6h98CFNznt4pIvHyP/qGMjz23nrjPAgnZlSGIJM6/vOdhAHQY
2qRQFyinMJ+rGmAn1bxFlgchqQGkc1XPCRK0oubyu0nkmP5/ghIPud3F8A1g5ISAxpwfynH4KTJA
yoKM8l01gaVy3LWZWsTzxKpOEGsmhx1Oyp2cp0XNRKEYM6gZtQhZwqKnea1V4//QzG0O1W01ayo8
7j9VYNSbZDaJA680vyb8191j5J5V68euW+TSiLbHJvneXOCCU9XKWlZ9kHaUeHSY+1MZGZDhFM6g
HIjBBCoe1JoKeRkjDFGPru4XyTgi0TcDc3gLMrCm0+cuknbTEmc4ZfdBrC6dmSUDvI8AExL4sTCh
3QVEFL65pXW2Vs2skU25ZdZ7M5yo/jFY2ZjvT39GrciKkcz6glMSNWh3/XIzit2lCVYCO/GMoMQ9
m5GwAK0TZt5k/4FzS4lZRUYYo/ff5YcBZsFgmljXjjvx47cDlVZQRM5e/iwC+hvFzp7rqmUilYbR
Hu4z6C3s7LvKA923zl/0y92o+Dtk/VPcmJvVA21Pl8KaXT37aNKzNFzjSEGoMySmvSbRmq4MKvrp
B7hMbm3mVX7fv/gYoNNa1U9EA7bclDBuTjczJf/Xeu6aCPeiDLuXK+ioegNh6fIJM4dlhfnVwgs+
zsIAqRLH8Y2DRcUmF9zyF8beKTfW+EqrIYRhar6Vqc7T8ns8/DonK8Ttb9nWBxGvgNxH6J2YBMJk
WeqIGfn1392HY7hrXtqm90JSdB1W/agWl9VFt/n4Cbezf5C+d9oEcwzpCYj4sd4XNuD7TMxwPtNl
+NabWBf35YVfluwEkrlV8ZxIACOtQXoU96wVYd3xVSagny4jSy1NfTpKDUReMgG97y+w382UfOVt
VxfbVHa8otaf7G8PUpB8FlyHIkEGE+C9ArgR1F91orVPb/YkpRBtTmPyJWhn3cYDaFuRGZNehlOK
pHWy7nLzhgz2MQQ+kxyJZGJFIyjIP8MozA69HXG+Xu7tzrSRXhpKRSGz9LthKzw9ovYz1jwMJmGk
DEDOHmpdcglvnP91bZrtgVAW3WxuB2liSLrTUFEVxnAfGJlBQ1yNONDKJTYYD4QcmPtb5N0i/55e
Kvi1kuMaRdwLhX11UBZW03oN7GBY6WmSdri+6koCoNDTrdOOLYkpH9JeNiyAFhpoG19UfwHIVwNb
Fy1+HlvXkliZ3/lCRLGycH2F2ocxPCx8jUhzomX+Id2N3mIXcflkLzrcxYCdzMxl9LIV+nJLVdw5
dPyuRcyFwe0uzt8sihhxY9EaYwC8yIWyX8Gn/DVmmi/rPqiXT2Uv9+0/kXLx5dW92fpSIZH7kaDa
hLE3vGO8k/3OOrE6w+iIV/b8yDt3iXGN51czR+g3TC2DSf+NnyHwCtbzQhup6rAZK56Z0XlPqRGp
MLcX4GEXb9e/7YgQw0AQY8pKyC57tRa/meMeW/222JTSn7R6WwVe3O1CMBplcq+Q8+qx9fNy/7Da
jCNs1FjJDYBKQh9E7MN+YY3xzpt3pFlVcizl4mHKyYCNw6OUr954rwMb7R9QaEHUdnWdxHB2r11u
nNiCGlcISHxBYLCYDW3iVwl6xYfg/H5wHOwqpzAUYijpyWhjx/xY5cz8BEzRbR30PNkJ6NoPeR2z
qFQ7fOvz5k/zsnjlt+XDZn6hmJmTeidliovGlVkAL5P7BvE8B3e/lT+yOr749i+aBOB9uHpPV5Jb
wln3K1gqvbrIgPMTTi9taMByKSv/X4CLr6ARwsvxSnXfc9bdKLasyUogGbwjKs2BWf/S2VqhwAk1
Akr34LASTlFQ3pNCP8OUCo94xuY8iulLKZ00FAC0OibjlfRO+Xaqzp2Q59ck83uVFB+Bjf1iF/FD
GDyeE62dpP/YZO4RbFKnV1gj1/XAMdVzdXIRa6kPkVDQG9BgEggtSfs9Fh1ay4+LV9d8iDfgFoF+
8aO5F2s2DjGfSe+Fu6LTPMSjvaylgsFvP+H6b9nxLbV12UchgHVhZ2c6IgEDF0NniJ/0G/xnQ8um
NjrPDsajOAbc6Xj44uPvTdZtMPU1o45p79SQygh87ccYQCEJ3ZIqzhahtFetRGdMOKoiGMqe3r3M
VIsrgW6rirfzXSelhjytA5MRBcdeH6cweaGXPpBAzx2w2QRuXKL0C1rrUw/HuvDRgtR2cPaUTGo2
pf2b5JJlJmajdaNRAoEjC4xmmj/O0vqTagL+Y/Y4gRfaSH+QHEnJDw+ieBQwWy5nN4eR50nmMA4j
qOFrYWFjl4CwMNuISiYshdJtd+Vm6seoM76miIVelHv6JwOA+Kwtcs8jhfCx0O/6XPdl2CAj+xYO
zThmR6Xxa98Fj7yheAINl1Q8eWNq23n/cdHDN6/IsNR2jVfDqrXrrPU7kvHBiqDICWmzSPhZN5wL
tS8YKZZZw9gs1+shaf1Bfia3DankYeArkfm+q2zaf/BI0EDq+yaTaqcC9bpLoqcb9ZlBpjZN8aeL
p2AQGrUHbWoY65GOO4hHLvC4HZ97mprXeZo8LxVcTEP3G3Y4DirBmJEGlMNu6dsg8S1HbdcEYJJn
cF79xQov7Vz2gU019mOuvw++BD8GcXX5RQh933EAE+qkSxh2fYrEbGzlDAJS/Bc6amAAVnkVH2lI
kzv3wtJyhpNfHkjwvmSOjWS91o9zFSUOEuXb0VfyZc3vmonJ+sD+FfTA91MdDs5yoYYXWWonzuoH
uBPWUKIECswzKsNbX9IFyiCu2ylqwWwPgbB3XJy8s85/JHHhPC6mbxVNyeeAU0coT6Z4+83GzgIe
zg26XjaU78Jy4kQ2AQA3p/H6iFR5FhUCjsBmpPQfNmxUcSmK1Xes1TtgUnRC1mdCQ3x9p+sv15xG
RC9j7cfBjIlBQ0rKsOY+VPoqdUYaGwoe7sbEsUCieUrboydXzJLaGcwraQECLfXb6/l79KEmzmEn
GR/tm0K0ir7hmE4aXvWqHWqxDdWE+ob5cA44cxU+Y6LI32iMiHow8/5o9WIivKngiJv7V0dSfpi3
+pfhlFRxLAblFFU5nwwnTEMo5wVNsqrkfIdvzGAEF+aOY+ghBIjktKASrR3qcKO9euDvda8yfnaR
k3YjizwcMpr1bNRi62G7K/BY/GxRrLmh3xrSySMnXyex909vmfjkY6t8RG/UHEe0wsdO2hCwLKZ4
Uuq7zPWOeat2P0EY5Uzyqd3oZcCr/xa195o40wNKy/LplTwoBNsKYOHmSDRY2e+jIKo+Rlci18Kc
+k2XolCUhOU0V/HzbdU4CqeiNjzin+Vc+PSCVrQl2NbYV4DSMRi0Vb7Rr1zClRftEg3DcAiMbfWI
ZwhhjkjvFXZO/0WxwcB8ICi6HoPu3Xn7EHncsB7pS01GPoWCPOvLPL0NT37BtNrj0rpzhjJEcq9l
616eD+QwyGZRQQd4KgYe+jG4GC29aiipkMbWEGLjLIGPtZVPf1rGV+5ALHaWyk/5BdUHqtfrmDxI
epcgHKtT70fLKlOEKYODsOg4MLbS4U3MT8VezAe9Y2uJjRQ0SbwzdfDgxJaRGuJLNjUJv4svl0jz
H+MMpcSTGws8TEc1bbNjaZCMTj8l+lyZ4b+RZ9XtcYDKn1Bv814kAy8WYZDA3BLbcnyi+AtyX/Zp
5zj53LYFUDrLnTpL7vSClqzXRsbKjHQUqhdhrcPcfsEtpJWE6Qt+Vv/nAs8hOntKgzRvwPutG4JI
fvScaFYn8vaq1Wc0+TfBa1dyb59j2Ize185g0JtHRyDYFOp/wlRSwXnDUD0eUhzo/MzYQGovmkMj
zks1qD+Y5Sv1TQLODEqlugcieaQVKvMcMOO/rstSpAtjy33+FB3LdtEa/Evt73/ET590qaizLYYk
ucZJYS2AZVlEdPwJJ4fCVCRTuGYKTIuJhGDObxT9NmGzS+54sG7JdiCMUnkKEgb7+rEnxzchjS86
GsKkKYOuGhB0mmLpGN+XGnTCUCpud7Zfn0CDAFbvWJNFaH8fIZDjokn4YyzF3OVscQYSMfQPkipp
DQQ6+Noalq587ADKFxzH4NN9fqYJfJDxkxft2nhSXfs3fmkdADmOS2jqpWZ1X+36d5G2DqxA1slA
tVXp7XBQrvHwhKa7ktr85QyaR0NR0Vpg466zvQKqyMTR7LTlRrLCv3U/9iuelH+/lfrpPxeunOCo
2OO3fIZW1H7NoTQvdN/0HJx611UH5psZVlvrK0TocT+bu5w1gUp6JFEdVXYDLg8TgOUBRkPIC1sE
wirpg+qoG64l5pPjls9ebMMgejwgQ11N7S7kYC5FkiNXRC9O0vvYL2CTe4MOzqy85l0TcftDOLDs
YpsPca67wn86pheBOrpK/u3YNtz8avSLopn8XomhpKocxwy1inRZ6VspOSJEUhy3djwMQJ4BsrL+
7YtjTJClSCW8vmKQOCDhmfXJUW307i4SW8Ph/4n6qjVZH8IOgt05k7ry0DNIKjMFCT2tl5ASScpp
GhmC9Zaj42vuWZWAsA8QpJ/nOvo8/uQ+e6jWNxcEC8GB1uP49Mhv681sTJ3exb1BMheAJwti2x1M
yptX7X3xN8IndiasJ4brNL9VS3ROJN453rgsR4tNcPrMfsUaD13DlEQw+VxK/xZcPC6jAe1S1dUd
3hybwqWJMoYqbfqSHG751eUe7Lv7ouSJ0UCutG1NOetP1Y/cZMV1iWioFhHJVR+i4UV0n49g1Inq
X+v+0AgMXoB6Y/c5Zmxdg8XwUU7EkIxf2OiuEG7jivqmX8nyqHN+5aMLwmL//9rcaPtJcu2pC8B5
TSO4/VyzTQDiUl+lBQProXkUvXcLXk2tjAvlJBnoco81rAZ2C/1hozsiQ2BtRiMP/a3U5i1tyNEa
k5PSMfwTf+G6pcCdGLqCtNpj5NBW2tDrqPRop0DVxh/IjwtVnLFeKVKDxAJNIYfAvRZ4it8zsVmw
UnphtweDBSlo1TltwqHvyTR3PrmAabOVVyCFt3Mu/IGDizz/O11w1O58/qh2vLJTokXDGQyuBRq8
lvdXTZDKC8k2mKEU1YSvA2QJRxTogbSa8F60qOY2gWZD21QI/CV/5X2RGhi98C0CqUZHkm6ba+hS
Q/aE6umBvzTvf5A1ARKLYkN013g68RmgyPV8ZNKJCV80HF+B5+7VxMsIuRXL0TmwpSYrjxZPxUfr
TR+/kyo9wnSG4LHMMm9efUYb0IoJW9v6qLk6CR+XAvSpEnYma050yOs5RFNlbn1JZmnDDkwwTKbX
ssxpk29y9DmrDS6jPcgD95Wl4bsFzPlJ5uRr7Bcqr/m35Yh1Nsq+Yzt9zDe+bwEZiwlhnSEWq1SK
OS5th3bxMfrBlUEOSPfB0ZrQWftmtDPW+uZNN46ATrIyhizZi8IgriJQvGPBuRVn8P6aAgn87ZZp
/iCDT8b7iaFPyoTIZ85xXPnRo2x612mJzmkgt4EzdAUSxd/xxBEHhHxkZEeIpQSmdA1Gjdu5rie6
TWwZfcGU3RAWWgULRIs8bcyysBm6ApM4zl9ul3YLoM+y6ZbkoCq+dwNE0hqt9dVOm52XsUgm0dEI
i8JMllcR6Q96DU0stnrSoG0fF6g0upu8LA0up7C7LW5Qn37nJx7WZSOqOT8FO+vv26xph+GP4kHg
N/dV3L+0OvypIxF4/Z2TVbEA597fwgUccedlOsMvThghB/ZQbU0ZwurISmLlnO5Fp5+9r3K4bTw6
vTzBsUD0sZ/e1XMy03qI3+S2Cbptq615SBm9kDs4GU5R9RY5yrbv1Clz2poDmPNezpWUO0CyvMAv
Dl51j8Faf7Yt8t0L4IAkNfOXgPDJAqqX68tQg8sjQvOsskdr4VlBmrib+OjGdwcjahnycHopyRDp
0iHT66+JMDp65ZQlUUw3NNV/dmwypyxe0AJoplo75w4so7WEowpxD0vEXH0rZGlDMUWqXCkB8pmD
TaAyLzDVaHH56CFuEzqQCsjm3ZphXpIzBZ/82mZeFyx7zHD1fNaRF36CgeSfo+bYemlf8XBpMA7i
s8N/cXKVW7nDhQYd4XJd7kAXqoGBCirY/GiZWiKel40cYqUuiLOUqYtChMBuWOMGS8RVBwKBo8i8
t8JTGlgnQXr6PvOqaU1KAfaoB5RX71dFo6D7CQvI7yEZs4WluRqPGKuMKr9iYqlIbRX8lK4/Ot3N
pYnosuMZxZu6FMOnboifS2z6mxWnJH6IqafZym5tEBaUtiffRs/9kd87ui7zYE6p9hr+zNAUwjQ/
NSmO/fa4oKYpY82VhKO+WaBJtuevX/64deGFTGs8UjOoM3FFQ82osv/sEWKVwYL20nCemPaHwClO
9CS5hlhIESL+oX8PyLTIFPau+Mp7qN81U61+5PlvenAL9YqfFdf1GeUbvOGImDjMHOVvqEDqNFAM
O/5yuGlqDgtengtzCQLOVsSSOf82OYokeWfkvuKF31w+CSFsayz7+I9FRVVOwfp6ssWXrjURi7M0
CwTL8S6C5oc3yXruLgbexX0T2Xkm8SloIxVjrDTsaW5iGGNWU200ZcTftaffNqzDSjAE/kFXPhPZ
MJEXXI9tDqcgwEPTzY2WkFt3/j9G1mO5pETclIeIyKhkjBD82BoIti3FfKV40rHBy6kq/Lrt6EnR
VMvwUezDJtY2h+L08r8v6OeehOvyXEz1BMhU6I1EgdW/QoL6lmQjIRK56L8BgtNXbi6Dd6k9Ts89
rKSsoxVobquD/vKwGlIBU6XCpWbRetYVWR64p204QXO6W1ocmHMjcpjHMIsQt64TT3OitkHRMtGe
WAQtC2uFrNh9Z1VOyp4qoi8B+IbwsuWUzIK3j6cPme9CLVf6DGUADbAh4nt5fzZ6kTGEaZcrGpFd
yM3Q9/8/PNieHNUQa34IgdtaAecpiJcmnkYhXjPfp1ts/3/YHGdFEwE06b16IVYLknIDj5R0JhG1
VgcWgsKK1QYjtXI2LKLYkWgFfThQF/nh/tf1kCIfEwuMZHZgNkiZuZ4LmCVGFtfDzE5+KVS+sXSC
qyLTz2dOHuIjoC/zUsAM8KHSLUFZw14gEhe5WVoeQ1+7bzllmoR6XGHDbRHopywVOIX7267/IF7T
dbEQgObXGA+p13KaL54sKlLKIyregpZQHrbqJVa7GQZRqfa31LepjPa4aEuDqe0TYW+MkwqhfSTe
zqh/bREmy47R6vYUp++F1gFEES+3k9yuj+vpb4Mus3KrSZI2F6/yzmpznL+9qZJhzmGy0tdq4p26
j/LHLnKw453yZONsdtHWUBiiEJkt8IaeBvy9HfT84SYhVld+YQtdALYclAgK+Zk7fkc+R8c0ljf3
8XBpP5UNN/N8j0zbG1MbslBU7auC3RX81LQ+dkzUzGVGv1o/HsxWVQl+zxncPdaaMiSQMfPrws52
Lk0tDnfefKn0BSkm9DrOV6zpIxm6NR8dCJLPWyIQ/40HEXY/OmsL/N7GgLqECLC54xWiToNKfuKG
CDtK2BYBsaDYuus4Bao9mYP/n9z4ekl7KShyPLhhukFRqDYekSYLsnu9XfSdhtEhtHOIEd8MNDOf
GLpbxBGE9JvDhjkDDURHteEIwqq1YZlx53cChJQ0nWU3pacyk0ctmNNXAEzfVWIC4hKKuXXPcMfa
wo5zZlYKpSk9vcgoO0v7ItkWD2LJa14C7JmoPyiKAbZhhb+hhhzgvqJ+B1ERa3FKbpMdPlFOougw
K9UX1z9akWsXgrMDZlzM3lyznVAxEMs2T9ZnIfqiofhZGoQc+QYPH0/emHDWjksXAlit8y5abMvC
TVISugNbMYIsmIzSveqgvbBnhVDt2nEn0jmspuo9SRKpbLf3GvoZQQKM8uW5cMn5zDNsIbptFIrm
TGPisM/NaCN6XU4v4LBA1ifDJ6E9DeADTdl9V7aBQrMGD8jo6NukydaZ8j0j3zU9M+EeMayloh7t
KWDIL6zV/YTtYOFd6aax2HbWWSCpbC+xroTrzHwSfxrmQ+oCG2tROSdwKIfxbovlMifJZPXKrWDO
lzVC6XkPr1UiUOSoiYu49uSpjKyPl0s2Nu3c0hwKKMrrBujce8LFQQaoyN2tMm0zXdhOwZaXs2p6
4Zth59sd+6wdHnJ1TQjShvrmNDDlQklfdwC0kMrQWLiRVLWalrlMj0dlvaZIXOlvC7NZ0Xr3oH+b
Pg+h43pa9gLu6vGxJPn9D5QM+9tkX1goCyTc9782WspO4WH+wpyywZJmkgvOTmgPSLe/neumdLQ4
eNN4/ycsfaPhjRFBTjCjanlg3jIkL7SKNnM1S7Gs24ZpU2B8B41SMBDHNuxGwqT7v8oQK0ulouhC
3guFXfK9iYl14g5L64aLuLrXxcELN5V8tg1cxZYOUPvbJ/4Jt6w02GLZv+9hl/AsMa1S7ZmexmvX
w5cQGX5uhodZ883zkM3O1ZmMt/RWzBjERO1XufguoJzy7oRexl1ZPG6lIK5eX4M0cwiOCKuw+3mC
PZwSgeVFVJpSMRb0fpTOYXn/2YDCnjpWxNdcXZCr2Cj7K6hPDfTfyWr4Dlpk3VcyeQAL5Utf9Rx+
/qefi0vWH5gEdvm5Uh5lvaRLho6qPxWvvE1KiTdFsMZH7ixLZBjehkZLFD9ZP/sy5ahX2q055xa8
eOehk7ykgGw05rfQdej3EMKoH0nlFNTDIaG5y9QHWwj/eNbqBTJ9HFI7dKINBD2h0lOJ+l2t+6XH
WjULJlWTPBd9HHeRA2waE0EJAB0i9Uf3ghEV50gLD4Pl1eJ0mzK+AGoZnq+i9YRrrN9JGoElbhZt
WVynBtQmOL8rFbZH8GXTCfsG0LVr8cM6iHisU2CliOErAYzMdkW/0HoXx8XB/Lg7Cxl7+bC1eO3w
jciwxLNSapDJGeLM+3ZGfH8X28SIsaAE9OjecpYNKq0NP9pUFhGW+Kw8KNRpwCB2NeqqnukWU60u
uhnLTKwSCbcBDVm3xdZtIfPDl8toq3IhfiNZfSIKw1oHuhur2g99gypK/VNSGVI8W9Z3yOU79GUU
CwMBj8u6UjWh9fcUbi131trlOrhoQPF2vERCkLM8daBZXgHLbRsOtyVj20nU0thEby/0+RCk3eLZ
pDWqBs+NsG9Nr2G5ZdBW0AB6qGDYyPZAgYkcOmaL9sJqOxqo7h945NNL07Tpen+qa+6wVjciCGxy
oDHV1ZJhBnHoFEkpaeWxDTjqJBpzZons0t2o7Je6BXdO9NK5Q0T9ihJKfB1KjTC+r3jInztz6ERw
ZoKKRFpYFg+boUmaOHOCvLvA9TC1mrlZi7oi/2oWcbIzT6Cbgg8+k82yW2fEQ57ezoS2WrTriVdi
bUcOaLhWRhRbT5/3LPdQlljMsS/24LWxjzFEFHoV/DYGfZcv9smO+foVro7M4e4O1iM5dK2mkMSQ
hUVeGRYO7YwpzlaZbtj81VzBS2JO15HoxMx+a4czP3CGjIGbWS7yQVvQCKIXi5b0xCF5QjAI5Zzu
GhpDaQ1JZz+ybHhC/XWXTSgfMiBBlxl/L8GDZET/9Ef+HqpYtyApt6N1NtljHHe69bbJQHEKcEKG
Xoj+gCU2zgDNXoJH4e4EEO1mgK8Rn9e18akmhM9dHBcMI+n9HYQFKVGc3x7LOU6mWrRH9xdkbLKi
l7JH0ty6XKV4oxU6TMlDvyD6DeE8FuI9aJsqz/l9xqLaoHJ9U2jdXwTRdBVKZVBw8GtoixwvmiQI
ptZMWH/t+fp2+Z6I6d2C1bOZxyg8rpKFmgo6sLxy5gFTesWKMtj69W/zNYtvwPvcgTsj13Zprpw1
I5xoO2pyGcdPKBfyPKeYEeJGW9sAxF4MV3xdWCaIPacdlq6rFtlh8G1AhBPbJnmrIDX70vDK59Qg
ulwr+3f5i5m60xly6CeXLDdDnSxwWcyEY2NsdhNo8nRznh+SJEhTn8H92BrYHeTLis0XniL/hJee
ln0hL9Jw48qzx7w26nGo6YOxgO3LEuZjI0SjQYQF9gCf5HSy2tZcIEvnQkPxcYvHfun2knr8rmVO
C5fNncjrXp7dWwszdhqL1aKzIryrBPXpItuT4ZNthdnPxoqighA8p4sP0Jba0qVFFqoHuoOp7gN1
I+ZXpLKxwo9wkGcGNUlOpg6lbApt72z8zQsIsD3CRjjtKP9KAExyVsziEYdSk540KEWxMXDO23+R
iD1QgbJxvXvafx/A7Gfiqg5JB4GwtXv5/euUtS/EYFOllYXE9C+XZ3M5b46YvWbGX8tUI0/VNXaI
oTbplA2xdNXy60OUakNnd5CZccu64xXF/6/h1Mj96IjsYSgnou7Fjrd068qmCotshX5vn/XZWmqN
pN+VLQmbQLEuDYwiyob5yyjbjANz/Mo2QalnyPgGjm4haPbAcRUMH0T8DDUt8wb5ObAjHnivr/ur
s24zr6RMnjNBFfMd/fznSgBuhskzzELvnsztxii6mMezIgCb2OLpWU2bwc7N/pISLjRRcpOu87Rb
HhSN0a3kLOC0zvll0rUCLzoGKCi5xkXeEFqOp5IMjgq+JJgTs+L7uOmmufewMCmJ3sOe4eHOUcdu
e8Um96ZGGxkVDnSUkkFUP18IHTyytNkCKCX0Qy8oM+cETDRxEdkSUTo2gebBYr4NN5q3plYed/Mo
WpxSv8VJv0YzqKOi4asIx6dTqiQm43sxcXn02wGZP2ciLHsmseWGrX3cZfWRb9qavqGp/G6RTVPD
AMwDrqdV9v3QyEgXDenOebUXSwyS75ih5n4LsJcn4ji1PDF4+zT7/UIDQ9IV/h32eG+x9B8NuTIR
k7cobJ3jRRL2OsIQM0nvGrjR2b2GQJAi8sL1ttNd3CaOIOPXImSomytsSyj7ZwoZixDaWc4s0mwd
9kcd5xJ2UpeJv6G/o1LlkuQMgTLfc4Mie0mX+Y0QPvOYoUM+FxHYchzqEsp135tUq+YqJq5//R60
MmtRzzGguC2LjrS5/pb8ARrvHK6X9gHuVTP3/lNqiBEgX15bVpR/67mk91oUp0mEXwXogWOqOMoN
GHwUoT1hGWYyL5944ammVnYKisfn9ccD23FpSGq8o3cAhZCwyJxi1A+r15kIZbWH6v/mB6QpyZw9
cmve0bREuZ3UOavJsbPmc63lqgEukTLhMO1EpnOjrz0++HH5jIrPgSLATn6YoTHWFRPnN2+yuT3W
ob3ixq1nMKbUppjK3N3JrgnrKjbmcioUhjbBccePYxmRPGFS2BX4DAHODLQv15+CyYz4w+phQo0W
xUsMduiwRcD7fd7JqPMebED/gMl1LSimi6rbbAnoByEkV9800IRxc19u0HwDnnjdVaHLxOiPRrI/
vG9onQCtz39gT8IZZfua4coZO47g2pM2J5cGZ1uz4CZTX3hC/0b7hVqyYL/Idoc2cSeT+UTwLJYn
HjqFytokOLi5oIj+x5zxgnNNIDJlNYktW+6Rdsk3vy/QmC/SYka01hhW2J5aJY+QLc2gvz5Q4khf
q6Qw1OWiymhF7+PLXZAdzUVzq9CGBH79IQvBiCvWZRQ80isd1M/lxWwwXQtER240qUT6ks3Z1Mcx
ikTqRzYm48Kl69f7YpCLzPwSSb6Y2Trb79bm+6eKkT/pIW7swORXJpmcLV6IKGt5FlUl0wS89May
QKLvv81pCnNJurwJQy9ZMI3GChCgfkErHhkrA9yyru7Qep3pmrNLX0cS7H5dAZquPyy76VgbJK13
7LrGNLxCcbPpuR7Adf5Rfc987xtgB2kmIPeRToDUwIHCMocct+1ZTWi+F/DnplBqW7TquuyhioQk
wph8pM65EarDdr4yGzldHW719SmyOIoGYwdBbNIZwUkg89EicSaW99LxBpBcL94JzkyDvktRfXST
Zvyx5x7Z2LHk3+vhBNPW+wmjFNDVnyzOp24al7LdAVvkFVN61ZjfDN5fhDgFbWVdcZZqz8NtmI4L
5bG6fI1SX4LdQDzYjZSV7NGL4nzr6J9o7nTp9YIe3a81WenddLorHohy2WOLKIXx66homXABHLkx
SJ75QA47dkf4mjDVDTMwv5BFzBI/1Jn/u1loBbqQmkWlFeRrV+lzU8e7leqUkTc7hXFkhSD0M0oH
4u8vcejhl4uNd8rJP8nzgXKrhu5zZmrCrpqcytInmIZvt/sQ+CnSsPQNGfuUKzqOmJ2XHEoNHXZe
URPe83uuyS10qhVAqwtUkKt1XUrdbspvKxqIsye7eZYbJbAhywGEpD+JgvhnU4YQWNjFsfhHrkM1
0s75gNnW9rfuBxC7ku4QL9jvE7jht7VfZmlAXT6Lt13Qa9p0Vd76hwfkGR8hTZbCJD+y3xkfNizd
3Phs1pXvMrI+N7UsNjgZ7eVEXxQQsWDDcIjjQ9cZ2q8QC+H8Dxkm3NLdL1dmRxbcpMSXBm2fK8DH
I6sIuK2bSfZOoAOVYqbokg/+qd/H7enNj8hPCR3BftgLB7BKDsvJ8kdAJQa9vwXSypGOvYSjYv8Z
JeJuRtvKAnxQtjKYJXq5mWE7qwRP6XVLDTkwiaDVw4Rj7J1D4Ox1VoVvr7GFPd1rrkgYabn0Ealp
5/IhuJb9lVhac47paQdYPO0+3vA8GaeFSFPp/8Bp/EnlCUhzxqVatHG2Gzi/8+ElNURJcrboT/AH
z44otGkJRxz9+7+Xxi99kF0FGELObEhWJC757Eg4Xrl6tXt6aH7kHCD5CtCcAktxlyTYCwAPdRB/
N1nspJfME6Zw4NXC6N+LXqYIsMpovOWxOGTXayHANTi0/qsUl07EOG4/+MsK23KIzd68+pDTyVRC
BP+GQQxA4t3MvzyznlXdDcdIrWNrNh83CLgtSuc9IBd2v+O8BTgJf9HFwXbhh6KAlZEgWlTeA6il
8p7FYdLIqyZlBx/zy2IavmxSLVSF+VbGYxtJTmjEmXe4gCx+69PWf3ky2b/7UyxGmomiWW7KMZd4
yKu4dAHg45/SIJA0jrWimI+TYTQX1dOqKm5BPI0pnjowWYjRs9lOeXu9oY76nA89srnCS9iaJtMe
+vC61BaQAV9aM928Av+lSa3U4G/CcrPUSocajHFPnQbkKsZozVaBejgHh56CtjuH4jd9L8/b9ZCU
mU+IqzG6yy99UggImriBGbO76eXQeb37wRokyBtxjVoiYjLnFCzR3xbcUq4p6hM+Se5QgIOEs0eN
6PV/FsTXPTnUjNGOs0UhFGIF0KIW911J/8ciKxZbYDdXayB70qEqCGROIjs3UeuPjQ2qShpNY12g
uowfrLcWUNcGUJbTzToiGRQsOdg7yObVstecJ8i3CC0uGbTxdMZmdVz0rmvTpzG6QEVGVjsj+zFW
EfNGGM4amCALxFGZ23uEcQk/k0yxrEx9kcEaDESyc/z8lV6L8c/s/8iyPTNg767AOoPqZ1C45UwK
qfSpPNsLtATVgskeIcOMETRLX6ISb4QOvgt5blEAYsOsYXbHh5Dxs9XsFrjpMcVQhIZXX0t/2f6D
V6D+wKtJhB6l4gmUUuWBW2kHmgGzzVPTu2hee23vXyhtf3GLSPkWZtQ5ZEzjWCghXMRY7wn/1+fy
VuzhdSiq319pFq14SuynV9BqVmaG2vI+nhdjNcw21YgPV0jUceKCXJNM6bCJsSIIG3bgaJqKcS3j
USdQF9/4EciE/RG/L91nuwne34K0zBy9WxJ9SavNnu1jk+29kVt8kMcEsbmS2HryWRXa41KRHywL
bTJb1gY1rQHL69aaUuIiXFDDgibvNgirHTrYnbvsgvYa19X3YlebGsWOtJIIZ8OwnQyBScNSa1pt
grVZEUWRHg7JflW+WhyDMd5waaVF4Uid4Sc0P5cHE8gVDUx2wrxNBIovJY4NyIuBJO+YGP8ZtWh4
jpT873ybjZmCtXG6kOZ48ErWvSoppkqQCuzp2eeMrW6ZKM1jg84yzR4Cx7s1IPB7LrFHnr97lU9K
TOpInp9qFp2fKlAIcrLBx4w+FSo+cgs6YYLgAhqwW/DEbgrHHVaJSr/rc28yzwOKaX193iHgPV4D
2a5MmapldB0wgFeBqbsc/MAMSWCXNasJGigWbYzZ+guR7OEqFvWGYz22gThc8j1LdKneN0Q9vrJv
neytiqE1FAA5EZfI/QSSIN15gE76cU0mDmSo6l7ViN4pJMKuVgD6RdzpcLKnwGqW5w+F961Ih0xQ
wRak/cV+HDJg32HvzqT6pNXQUqMuqKHDvlnqLSnzwYTsjpogJ259ObSgrRyTFXVUfSChpjQ+fX4v
w+UBtVZcylW3OV/iXuT31PsTxtSz6QvWcVOvHwRUABKnLfkzkjubu0lD/rhhXlADxw3kgDJSEqeK
IU76ChDzJIvormfhaD/GsoHABk6RiL1mEXqcchYV30+mDJwW3tJ5nd9bfwKlSDNoGmBE0BzpACvi
MOiEkJnbmBYlRgDkNGYgY8rk8uoxQBvd6R79sKFU95gz1Vkc9u0b+HkE0AmL80JC7A4hPFb2Nbrp
CzJVeHuA0643q0aKkROJnb44mk6PJ3fL42gK6vUIlGFYcC3R59SjpD9dejwGjI0VhimZ63uJNlWb
uExXRIf4tn/CeF033gkOcP9i8q4tv7FKHnyAIGRN5QbpDVtPVK0VCfhBaTkJ/w99mL0yIRBejGFr
6UtJUi6pcet40LFnuDDwmbbnTZCWe8FYrRU+sEANgBBYA52/9ymMqCvQrkYQDQkgHxRoHuBeArB1
gQQrmBlS3YRtzM4fB+S+dLpd3n/w762faI7JRAIV5mhHPwKcpGzOBRK4tB6vr19xa0aQl5Hk18I2
47ZZIWEVvIkLAB+ngEFpqthXM5SFafJjqxmoVVTtYsT7Hf66LfIdnMtRUbfB75nXcxjNqaIsBQNw
P4nZUGszJavkyAYSovas93ysX+3Ujc6+8beIzayXLeiS4bn8jjFo8IyXxcfDM/zppm7O3G5OeAa1
u3bx/ax/UYWuNaaA8ZEPjY47xkAu0CCp/CLn4iZTlG4GeRYLQ6BVcckZcQu+tIzShlFK0qAFL7GN
AvjxEVKaksv0yl/83/FK1WqoE0vNK3Dbg0S5kivIrCM5N29J1MskmWXOATHl/POz5Wh4rowEePL+
j87ijNuipT2vqwK2bPaJow+wJxpM1lZNNStOIzN/4/3PZYbUG2obckowIUTGf5bVlyTRDiSy3lbX
3sQjbl/sEA44CJO8YKEmYISbaYKi006pebU0feIOtbetsGXYhU3yeaJBIK8kkab5RMHC982MFEO1
cV320BmVIcu6fvTZiFhY25baZ7J34jF+7JI/m5oR4MZlyxbVMzH5vmIsIDrq901QSSEtNK06c0Se
Er9a2gmiWOG6+Ku9hzMXyepNuDzh3CJmJLMqdQldx3/SjFW6A62zwYK7+u4ABeIpZsVzvG+oSm/L
Dr8QcrVMXCcHt6BbIx5shLVYmprbxeV5nDgCCyC8qAtbm22gq+itHto8yZVlZo33FvlYX53HN6IA
1P/wOLqm8zatax/gdhA/E3Ox+99bGUsGwqwpyFGIRFUerRYLarF+mrpscJSpFHBMiT0cfGBUZ4Cs
n1pz27VLm/IUeapwQNrAQaMsDZ9SVWyugI7wsuM6BAVROEYbauie2IgBHmfnvWmJO+ZEPP0LI4Fq
Wl3Gxzw2cOgfY/ySGPH1aUrvKizmzq+APp0zj1h2ByrzV4YzLEkYWCnQyc4TzYCp1PvA+dFtFPqA
ZFRtb6VKvdCs6L9+TeBlDznWVJh7LSm7pRY91xaBvfHMSS+YMc2v+32/Xq2FMOh8fQVZma4Js7xE
gbYNTFHt+HDh1Tq7QT7+17tjsJ+Q/FZpFmqNdGaguTyelqIA2lNfcLrl1u0ngqHJPmE6K0hbn//Y
bZV5L+g0cP9Ca+Fs4lSnvDLmwz9Z0PhUGqu6M4SsvquMRPOB61eDlIBGT8bfCmFAG8jYZBs9j9MD
3cz43Mu1M71baESztrsqQFHvKPI0KWo41TcGEjyAnnSIxNnkUMypG7FPlQkVUj/XdTVE5i7eDrsc
zii3JQ6/wfwKL0mIk5ekBdCv8rhWlSqhgMD368LrOJhLYTDGbwq9d0yky3039e3g/W8PSrszOx/b
d99qgJ/DkF+llArVXQhCJATTtrZy6DDFwchNOMVrHHIst5jOQugJVm9+Datev7aFj/CRwubXOXW5
Oaj1IhhP/exF/YFx5VaH/4vZGnsXGBtGM3vn35sLP232zB0HIpYq2MkoPKGmV6NVGwj9Xb799yCE
zmeI42TwmBh/Ax3c5P0fOWVzfSv+uS3KYhgpEbD3fN17J1wsYr0vYs+aM19xZJuKxO2+WvZirAbH
9wWYG4+joYxZSNMyasfw1d73fBetgJM4tXQfAbgyIpKlyUkIKcE/DBWrajfXyqyXkPwmRHA0RLdO
QNV6M0RcH1jc3f8VNTKybr86HzuoZUx/U+VkTxDZf+L84kiANO5E5h/9PiUtwggvQWqO687O0Tp0
3GUIxRKZ8ZpwEVEjVd1lFdyYRrJMZ1fIzClWr3o1VECtebmuoe2Jp8IHxbtfN2dTCwTdr7g3x2A/
+B705Pa5YPC+EqOUXJp4zj4Blx1wL0DDzzQs/VLWA/9p8OaqI84+ENvRr1zUnkj5SK9ilkhl4NVQ
hWj15OKf+yq2GxtipdAgqT2/qQ7qIy3jsivH5mo3LUAZ4i1U2VW54rgnnnhrZu31iWjBrMpUnLK0
bfv3tbM3ixDCZLEK2d0rSjkjl3rNaf1Z7SviSACF8VNPGcAr77BfDqkPwhFYJwIn5/dQiyy2F3IV
0/cLv9+Tudf/YaxFq+4vemiakcTSn6QczcmNyl//5pllgtkxdP+8gAoILZ596aNhdih7+TJxqwWG
cTEqgd/QNqhfGSkfhfTqN8gKCfuGtAgTfw8UzSuRXznlpIYp2jc73xx7FB/+e/KZ2A69N2+s0hTo
QdiaNJFP1l3yD+4Cl83hnrI4m/ZAHZFPT/kLGYiJ7E7/SatW2OhXTWpWj8nQfsriRxS514aPxXHG
rkzZK1ljI6NAeHcbEVUDjxprckR7QSI1/G5/KTB9PrS8CUh9vOT7Y55Xd8WOtXrea6oaoZbwh7Vu
+jicyc/PBpKvBqrgqBDLBz3cSFC2865eytDck6/LmQFoMHrFYx4b2ub2DdHUXhr5fryPQr/mmZb5
1jqIgZO0X2mytkAiV/mA810a7jwW7/hw4DyZrkc6fi3bFbxbF9y9PPr1hbGMS/PXrstEhnt7MVx/
e6a1pfiREF9C+w3WJE0mY68IcpoRja08HOjHYnCPHKm1ej5AxiN0eNeScUsa4asqul2K53VCKrLB
PumYnILo1+G0REdT2NLXOn2gBbi0+jUYulDWQ22RuA2HQx/7/K08bPlVAOP7AUg1PsWFyzSDRBya
/2+qRXn2nQnCwo6DR8bfNzsiHvoEBhWtD7ljncYn2vIrucv/1/JlKTbmrNMhlrPsRIjesKkLs+uJ
cVGoHj7roff1QDEXfoS/eB+UnRwIT7EUqLLcZhimRQpdztBZyKEyV3sHCSy2JIQAn93m3ds6KaxP
YvLkokakazOxGV+w442a/jzheDAXDoOIkHg8w6Zf6nX5ggIpY4YZO7jdkNyNmOXejCYg9wk7MjKE
hBRiMg3I8M4ImtNL+eGfaW3nUA7taAjSfWN5/ixEJmShtXR1wvycf0MvEqHR/lx6CjiXT8PZDvzs
phaO9wIKBizlO+KyCXpXEFdBJan6/DcES50f/ja2oWiQzNoizq/TN6GcreVRLaVp996SkwJTAhFE
GnWSIk2+VnatLOkm6yZPdv1qfTeJO/iH8QOKjowlG3JTZzCRV2caLb4234QzAq7cGp2nQWMjKqBa
CBX2tFX31umnkKL04Qi09plb9g9niqmgnNI4da/vhragp097TBHO70p2nerCYj+QHjcZLwhpO17C
mUJcwgT6ftu9GzxIGrySPBGHNmc7ASnHXnEpJihfVbQ1KusUWSmT6knTNZFPEzAnsiJLgrzWUd0h
xfGA6IyeLQdJU1wjKneb6JZq8kJKXkv0hKT3Oi5ihn53bplqUF7dCs394/hf76IK+C2VDDexT5MV
U92p4ymIqG1l5mhFvR/8EjmqsbzBPHw+SgL/s8hJrRoFUoJSEM2XITBie4FWCLE8Jpoj7QE5JFGc
p5wEjH8Zn7Y56Qzshm4ZWW52swR6HYC70TBxSzod/jeGfih+nUlb5l5Hm9nk4sQq+OpI6x+yAhHi
RfJ7qq6yZHudphx8uosKK9WA4Jt+aa+oH9JrGrX3+szOh23O3vJWa+tRWOQeBFd4JnJugm7K10qR
VoUuHY3NoAXcBKZ/WAcn+MHUVdqdkUIVWCAYKFh/K73m03LdEa3TcMpZn5PrjmkucWBs8YCNHXfe
inhtupynu257DzzS9UWGlJXjZdDtTL4eAaCCdR6rgQYpWbgyLEMdfwO0Yi7JdhWKaNZAWVuhHz2D
/zs0nRd3GI03xl690jY8l+zbLHhKENqc2WT/zj3loPq9BpUBES6QN8AkfV+2MbDLJGyXvgCEtBP1
tUPnHhUTkdUt2TtMo076aCbBywLl3/b3hqQDZobDL/gm+zL8YlLHJxML/cSWPUawdxflh2obqsq2
sfTZm70TbGeAE18/Z6+BcO7cXpt6/Km1SK4TfUqr7VP8182pfDDTsoIT7db72vpC1J73BMND3mdh
FGi0QmAKVIb+BCKQ5/EOawaXi0TKvYVLbS6O03oplxv9S6snN20aBQQ69B8Pi6vZu2axWWOV+1Q7
EzyMe3LjI4SsLln0uBoUIhugPkPdyCMeMpT/jO7ci6AqvV5hwim/hrX7l0g5kV3q6dtbR/mOriRn
r5d3jZwWMc/e3tLcj9ZHXhpuLAhruNLZyxevHz+RcAfM2gUdzXk08QZHWkhvrFM1iNMSXPToL7ZB
VdljTD4lzNhs/SP+5o2EcRuK9OX3M4j0DcDby/AklPrZz/lH/t0tCeUzzXM/CMA6G+HROaoxPIrh
XMwHkUswqrLphZBCp0xVa+C++8o+Nw1DgZYabFhr1cPwbbHm+Uj0JhbawHEl/T6f4vObGY25ajmO
p0CgvtpZUQ/NL2niB5u8ylLYLicYXHALcCS+bIOJUy+JIvxb/zwBBSMGqlHYT6kieaBOM6lW6xIK
Q5L5gJGQNF2HCVM/JquB1YkHX9MHOLSabUfIT6uQqbeSX5vCWi0MZom5qsPszTCo6D4HWu5DY2Ho
iJX2gTPRHlEu+C+y8sjNoP/fSA8MDf1JMQvc1x9ErODzqT/FGZBlB5a0EUGJvVWjyZPK6inCROtS
LU1DR2bPAubea07Fx3D1N6czDVmZYVtgHErJ0y2MJvseynu3R40gKQ4xC/RdXu28Do9MDmQZzO74
8FAqOymV9zetXO5KImgzqW4oLJnWHvA3nOT/LQnzQryS41tBwQ2ta1WmWJmE3PNX0Ci5+xZ9KzsT
hYoNZIQ93Gn/AhqKss29eq6lqGZe19oT8+P5xi7n55kkYGQIggIntQGcITbtlz8ZEEbHYwjzz7fr
rIM0X8bR7LboyOSgNU9Cs74KOQrE2YD/MAi7Xt5Utr+cx6J7rktKMWjxAdVcrm4b3IpgjhSERd1W
H26WVXqfsXnRciDONdZw6rEBlpq2sKiebMc974ea/L5ogbWyA1BDEE5ErQM2EURw2Qncgw0YkwIZ
futiUNAKV8XhwmWNX1znTuhCCWueeEBzYaIqeNXBkMjiYRrpot/TcF1rtGmwyRxRIdqpO3LDFAGp
Q2aj+/Oxaz8duGAHfYGtJrNGdbrOsS/12LQ7aC/dG01BRaucV7bNagvNhaoKqWbmkK9vVQm7COwU
5aya6z9aly+SHJUm9Txwyjwuj+/8nICgW00gUhrWolU/1Ozaw9UfmPzf7yJAyut9AZfZNWZ1DPTN
35JawO6jcr5e5uKKhK/xGvdMsWd6F5aQUHW+gd1zYv6O2Y6aCtLulZvhKwOq9dkLxChs360wxJOV
6KXttzD95kjZRD0EGzDIu5l5c19sLI+wG7AYk7pcwE00GxWaLNFh9VfIG2zavRy1ezjSq18o38Ps
3H6hc/LOjdoRhaGrZ7Eu28YddQS2k8DdKKZ8Kc4cZdRzKOe0dUPGuVN6i8Bx9/2lvM4PC4qqnSfQ
g5bIBbYKEIU5lhLwiSp+LPN1QpMOQNrALWFMA5bQGvUhM+QzPliPOE8tWW/jenCOM0m3ZD7mMAy0
0NOXHXPnkGpFA5R7OkQYJVimoUj+O1IouWzqttQo1FQth/xmFl3/keuXjhVmmK9jZY4RvhEzkI5l
raaIoBJtr/5TJY9YKdKgHe30EepyMsTXPNduU5koXMizW7MZpu4DTvzUKa6JrrgFNDmpBRq+7+E+
cL1IxLWAkl7+mvJQJXfNhMTAPUxtEvj2whTticE/I/dsD8cS1BSqCkXNodndYzmPudgrbbdSU23o
BragEVbDoXmtquWNfxBfYQqHLLe1QC5D4wr0lopK+vf7xFcNUXeOPQySAapkAzx7tQhpZvc36hA8
EhpfsN/zPu6+9OKTfA3T4dCCBjXl780g51h1E0OiUFBYFgHYsF+HV/PmHzi0lZZ5fVF0QiA+gW1q
Q2LjYSWu6GcUgJEKO0BfZ+9C3xmH97eb2AS26UvHmM1bI7RK2mIixPrGnqzncoe154oNAxcwK79v
eEJP12mGGUNGh1k9iedgqhgKogPopWRq2CN9Iw8Hg3Ysx9cJTdM30HpXwoiir6P9smAS4kiicfpX
wAwLRykS+Sa5Gq1x5EJ41O4R5DJ3R29xN0gKiNHCM+0hrsTmZC/jZiBnYzoCtvQh5ihV8aSfcL/n
fndTp1qXKMIZmPxeTQ5dXZuR509GeBkzMYmq9VZVx+wHclTLjtz+npMpnidp8kceIRtbLMAg4Vrc
x4ArGDshSj+EpDIyPhTNx9u0YAgIQTrkHFW3m4wrjVko7R78XD6n/v9CJ/mAvgmLYs6jY3FB14v8
rE9kpg1Vptn03nnvsfP5tyUStccvRs6BEI4jfzdOH4/K/uu5P15XwvH0SQbwFJRLiCMgi0a6RSZ6
q6StjSaCHpGhl7pAS9OaK1ZOQh5wTM5NZbj+WvOjqaPPOI1pSPtJuYKDOpAUjKCE4uPPfEwa9/B4
KpBztD9B8dWqGIQpIgX9s41JG2AgVL/yr4FZsBYaEIs/sL982oOP3jbFJgXVNvrY3GHvcLDl7Im6
j0vO8rqL/s/reEF9RF+HMKdhO9cMvU6bNlSNceg1jEFHt3Kw4m3EV0lTVQbucfkhsq5GLHPGZbQY
MxtLGVJbY2nmDfjzLJeSDK3a+pStnKyLeHfgMyuCYZMUqH8aXf7R/5s6VR0mZqDhLUJcQMgdJ+va
FmNP7kC1LDtzhvj4D4Zawfzlkei91reS4XhASZ21lx3ihCWmXaVkPofgUw7PSsx/W1nmRGHysMwo
gpaBCuBmLSB9nFYCi/ddg3Ml1ws1nexf5+k6zaIYa0vVjXjw1LZQ/EFym1yKvXHObHRwXi68GIvh
/wiEqPfqYB+8v8H1uwaBgZU5cyFFeQxW/27dCEIXgojCcaHDqEjsSp8SpBmnRvtpSy7EPFAUKJDd
aPrgDf/9xAEw1RJLGX7EYwMlj83kSuhNLHyhPm/BAgMyjivrAX7tQrZkUBKXmzIBrfGt8/EDHEpB
k+NPPgK2nXqf4y5qc1P09MyzBB/+dp05ZNMiwqfzB0BTVAuvlgMbzNGJlKF32gKem4HnVr6HvNTS
kLURWgmQIRo5ZfEBpO6ZNeSHKi3Pg0Zo0kma68CMokxRHoJtm+M4F4QEAeMQJwNVnE1SblY93AKC
G3zewenvhKlv5RQl1a8UJmsE+Vmftlbolbz+1/IlYmwXjniJhRHjgWquXMyZyAN1lMAWsqg0UZuY
NneClxbx8WzJBgKkTav/CpsG3JTPp4exgoq45BWK0jhs/lS+znE1iVrAMPbbxmk5ynMce9jKr1dH
huc2PtHxZVq9OeTG+inApahfffiEas3HmAkVmQKl8NgzsvSS+7BGVOiD3+6176Er6/ikwA/XSjIU
0BtQtJcxyXsff6Xt//uW+1G3wx8zEbmpAyIHY9VaKkEIJk69GkyuJ5fa79OpjkQ3L50GfrCvEVHH
pwRGHcTuWyxFmN1sAIdnCW5jnxmVQcHdvaMKkyf+PJb9TweLp1q5/uCI32iJYOxh5alFR2trh/+s
Hv6bKaiIKx0U5zN7NtI4htIq/vjwHhSmrmFM0UknVaBy/2i9ggiy1XvUeJqAPeMvU/Cx81YJlc0J
Fs/fFC2yV6ZTbja/mtYcysbuBUS9hZYvkNtHIyKQVkE1k3Eu190khlzx4+o9XTCh4KvW3LbpYcma
GgeWHLaZo5gdklu/k8gnwn90ZLvdCGtB/L/kH84SEpE24N56FN+/z/bf6DB9vQIbENUfXJLk9HT8
xW0WHxAOKpvpqvO2AaEoUuU3TlNhDFBCF2fMA/rSbsXNxP2P4ujP45uwCmK89Adlm+3QHqizrwOY
gC7aE+/4Zx+0DQtXf3IrnJpQCEN1YhBiXfulcuqw8jMroUQZ6Sb1+zQM3ZHmAo+zEtPL/buNJVvx
QoV4eZJIUzsuaz5HbgapPrKfK28hb9iQbqew4FDs9tSi+RpJGD1DhsLmDupcwk9S5QQe4qqpHSv5
zXp+7fA/kmkjBchX2SQIkn+jls9bobtHXfloPatGNpcFqmfMDaj/eOIHJ9vMiuzWM90vg2en0Y+T
4KrPmKqUedByuDsNODohioZUaHjr2OWrgEFNwFY3yi8LA+l6KVK4wGPjtkRHJLAaYLN3TAm2dTFb
xUzOBZRM9b4pvkidiJXw09wIATX2Ga9oYDPlkYz63asDye5xcPNd8M0dW9ytPp+6UcJww7ARSVZ9
dAS+DjtkF2kSehkM/Zm13sZ/BjMA9F7Ol6ACbK3Vx7rUvhGE27cXitYX8Je8XNZWuMSLNkrc9mnn
nS6qDubr4B5OGLuqBQd1HdPCrMu/hS+ucWqfr+wOrtLAvdZ29BK34wWUhbYcD3Rmr1j1kf6RnBQT
B/gCFoZndRu2Fhtba8Z6KXbIm04UYaIJB3soCyDz1AaW43U3V52HYlTeCAXAN184tQV8GHdG35W5
NKduODS/nl4b3jiYWaMmyE/dzSPkeATg44jktDYC7tJ6c7HC84ciWlijNMtIzpsrQv5pGXFAbTAG
Bd5aCBj2+DNrnOaW0FHH7hXXSvWiYaJJ1fqU/ownn1Kl/6ibpblQ2ZgRzP3giP0W3BJCZ6cL0hZv
0vx36JLvkumFA95R7J6gHbDtvYrZejKHeTatZ9hOHQDmge34QKX56xEVYQ3TqrppDksWV3ibU62x
7lPMOluGBeMi0Cst0IxvrjBnam3qxJLbbKrXPxQpYSrq9rh8Q5PeXI6utHbfLXdx7YQ9TVtqffjS
jySObYdvYAehqNIAg8bZsosEWdOBmFN5AqAN70AVgP9QBJtCv9e2axEwh6CZudsS0B0N7naZt0kv
wK+a9XBr9qf4KhDXAQ0YzwvIAhVbIrh66e5u7hNZiH3gFODlWoBd8UQwj5kxWPzPeLusDomvgrok
iDX49nDbjmKXJZ3Rk4qgk/WmxD/1tZNs3iehVGc6nJiRD7z9hPxTTUm8s/unzg8KUmbgsqhzMn/l
rhUqLtyqLwA7qE/LeEIagGXcOtKFDlVJUxHUbzY/2GoT7XlIpGCdvWSXNgJAhuQrLYgdQ/JhiAl1
e1D+StvKI7Qjk9CzLxUlAsBy1CmItk9j1+bhfwLfn1rsoqw0Ty5C+viq1+Wez4Xk0OzXlZDpiS/+
TWIpvrjPyYSe8rZUHdD1BSs9AWhji3CCSgQ9Pj7KFHioPW5EYcORkuID60BBj+3IM1GTvlKgz/i+
XYx6nTh09Uq2TxeqYD2TSpH0/8e896v9MiuuXomOufqKS3JAt7h5Jsp6Y/KTO9sU5XDgjAclQim+
CTupqtIwx/RQ20aUYSijXY+F7vN2S9O4y5oRrCytSGTxvIaLxF6f1Xcymkz1Gi12PLUpWOlnB9+R
+H58QGw6W5Yi4JQtICPUMDtpL4qPCP0iCHBMmRGsOK1nvItQGZI0d70pMSUl2sMLduLWGuhjepjy
zwqK6GW204l3G3k063vZW8CAw8diVKS0/65xIjfcz+31r102RLXKvr0zWnZdfvA4whBdY9/YaKwu
fK0M/xV0NSZ1PrW+CH29euPgSh6pKYjVm3Cotf06VWLTAS+UoMgmmm1cl08bu/D7d4I8+dKUG6AX
xCfjR8cjhd6m46phARDYrxPG+Wcwgqc01ZhsrBqgHxaeowWD+0j1+mu+H62axqPgcRFofBH8ERY9
xmUu2cHdfaxmmdEPNz/XRcZ7QXolbiZdt45WWqvbl4Y88xBPtwk7bPD5pIDccDPRIaN/qc/7VJ3W
sy1MtMSa0pn+AxiqWeZgjgATaYwLHTky3l2oTusZsNf3oJHGZUcFaW6D+f1HIIsauNBrka+4FcVq
c2mMv9VpinHqh4axIup/Ij9GPic0+inS2NY6KTgkwPuhmC2tW6HyKiMM0Pk8cRO2l4j80ioVQpb7
TFjIkhGQySSlI8sFdhKfJYz1mQnHN3qn3nIhOk4a5g4Dt4expk7nUOxs9jyCtMWHhR3pMaNB+VoC
uu/C+rsQAeKnichUzpsVz/4CxvKzgLz8qk4PhfXzy5s3o2tM91dcw6bB9ATy+J2OqTlxvrhWZbZB
QcrOm62KTXfIRQgbTERVhqia1lFYs/QQZkdL2e7Z49x6wT/YUCZUCWXJ0Yoa4Fp5yb45rBfirkc+
PSclGFO7mrbhQsDunNTBSGYozEw7bdhY9T7hSwm1IaKjYhYgiGAkQFGFzLoOifIbJfDJf+UXXuno
AQtQ8ObTo9trH9qJDbnQb74oPunHxVXf8Qxp8eYU7VQcWiuOFPp44Vcnogx3wKWqZDe8TLuR9Kxm
eGyURews1ROkkWxiOO1Y1rtq2NwZHKCgKMdlB/OrAOX5yo+eFTnoIOuVE7xnZ+q3UMkm/eS0tfHy
rI7207nyawLRTY4F56KnhKIUiynm/lxZvA9iOvJT1xPfansr/d+QsNODarsahHQuU7elKxU3yNxf
2QZdpxhHIW5tlzo/VoOuH26OpDU4tLF01Z/wrH9/++n+JxCUXp3EWBcDWs/V84iXWlwY3Thg0Xvx
je+30xzxD57iAG6wh/EfyZpAJDnzY4cKgUklnZFb3aOkMm5roPgzA9DejpbzHw6zMGtC0WXpxpmI
fgsm+TpKtgFa0ihGm37PYLco2SgsdPlpTjR0BmE4uNWFw0K0QAMsLNHnM5wQ/rVBxshiMBZGIiJz
tN3Rnt8L+o+REd1V86sB3ojQl8EkH+yxQEZD7+L6kaxfqt4V1aQJ8gcDl/0c2Tx8zGDPMJu0hjUZ
s0OoUyR3zkjHD7Eiy4GlQjlyLduYTkYIgx4WW6TLO5X6iXmxt6Yf75+ajrenPQ9pBsbBD17lc2wT
WTV5HpxoX71Up/km6uX9z+ne4gJzlQ9zZ4fWvkaZgj4TOAsVTCkRrtvfodkow1HagcIgLcvhA2Bw
bSHn3Dstdh0ppYA25CPQRNzk770DgTJ0dl6gVkAcekoha7Sg9pSRS2B6pfZQkSWOlTtK+IFN2y+2
56O1NGQyZ1z5CzWNDCRA1WfTO6JJx40QtvbAhoThMKJJvcOH42lmYiVlWDAzUIBhgj6ZhGzjDq5e
ooFjwODAL9UBFmg0eZxv4ITUMq70f5VYqKfJYX4qabhagW+xiRXwNtqiZCTfjCsvcJfeWP9mID5e
2qeZX9DUtWZjfXNswC+H2h51br1J9r26DpELdp6Bl++zrLwPHDAnvHZdNBzM023UhZ2ieJzQkUlr
/bKiDnVFnFxC3LT/sjCcUYpJ9060ULDa7eFnGsmHCNtCd+G0IG4t6ZjQC1FIaqhdmIoSfOmaroVC
1Hx3nTSdrXpIjs+TsJxh0Xn88xS7TuAtc8EqNp4uCZYvoBSiyd8lSX8xMhGKWak9jh51EvgXXHFQ
Jq4gsaOHb3p3YaHHTnPoCcz4v4v+IdcHC9rGLMpKL0HkGA8ihOehAhE216lvghF4LrU82WAqHbZt
xC2PFv0Ta5oBiP8aIKCLx07xJ+bZzDUzAa/NwNdlJCklYjMO1qIVBYrhOUeRu2eF01OEXcsL4/hL
ZYjm8yPGUbu6rhjwDJi2MV/DEq+snZPWYy0o0Ka9sD76G01hFS2HL9Zh4mEdTqr9Dja4UA1XsuMd
YV/cNDbUYXSfdLmCD/RQ4jyN74LRNV/n/vSHwTJMzUIqe0HTrm+V8wmAC7jk7arOS7zu431H1ull
eIDh9r9PDjQCDQ2qKVOWA7y3bwtgoqi1P7bU+Q1E4080gdqujJvBe/weIKDbfMApeq2mTsNevsRb
HkySC0dwMJf0eA0AyF3fBbdPc52JQ0unrnd/+n3gyZmFlpFDkgICMz9qgFrGRGiaONur0GES1mws
K2o5y06b8mJjnHdbbJQ4osLq+MkByc2f6v60qOoL5MXKqX83g7C23MAE2AjspF+QmbJCTHl3Zf42
zEjUEu2vAFM5QDOuUi/pMI6mXGxegW9Op82iZWd/6gpFxtzrBflVaiQPbk+m4W/Sjvo5dJBW4g21
+eZ2mtF+HnoRu91x52DGqQ5OjtPjIcyCeMqgVRHvuIWnh3IOSzHZ6f14SQHEZGhaiYuMO5ahkSzh
tyTBF7FBE6Vzy1sUf2rPzZV4I7STQALYzIsTTAVLWIv2jX8989MPIGJfU4T3LQ2CaKpZdxcyTJaT
COtKMNNf50ABb5FoGwnMIllqCHM3pFAqPLECADSeQ6S0Df5QGS5VufGOQas1S3BPb9LU4OqXg8bH
tOAR1YenZCik91RgfnCt8CLRfKK5/mE8ZMwt5Dp3M6WikmFFdxBvGWDGY7fUAXtYnRBeT+gSL15W
A43eF48FSAoVZZIk5CcDZlTBBqmB0JLbtO3+SgUDNw7/QXvFKJbLneIsLw+LLJKjkQMl0kIzQKD6
/+m+EybNzRaGKUoJkjxMj9TdBgdOI3GEjXVrNWWJCdmNzzK2qj/x8wJyUyVjLhbk/Hkm2dooP4O1
uYkK0WVPvmSwYuZmcCHXq/I1jA4xpEYGFBQ/g+us1eOkMj3ElTyMu5wck9srsXxuFywlmizuP2/F
mVBZkEPSqqXokGIFPQxNW05bp2+tawUlyq/48cFhdhZzQ5x5mfWAVJOKcpTi2X98AUs++MBICQx2
nCAXAT4tVeelCmWHeC4v6HHQeRaPTTXnhPrCq3DHj7vbNgTcM8j2Mo5wOMahFHjD72/ZzIKZbboh
zygGJOT/JfzQF2GcZRJFjR3tda8LnO+UllJxnNwaoVpJiI8QDP1JA+yjZiwUAZ3t710I0GEPTofO
LPLEjz+yMR6za7F0j2QHPE/rDsZwsrkx1fzkZ/5RFs+b/m/bb7m+KpiJorx1SaqVa2BGWX0os7f2
d8hg7vamso86S3XZGhnfcbXYbxKHHPBGSWeqhxCqHB2WLEY73UeyFamjtvqoYw2vQGZtg4pjOWrP
T+MpfjO9zn3+3SizS8PvvJXp34xrmkU7aJ8p1QcS4beHssnXNBf3iPgBoste0v8hyDK169rMz5g3
/XGtBd6XAxzEKbvHafmm9p4L8sVWcjtHC0/phE7GUFYKvwJguBka9jA3trostjUaLk9+RWuwbytL
Vi7nd2Q9p1MzCwZ/tTMj1hN09n9AWh0OKx9KSrBIOpbN3Zyidp0Zu4+ELuodT2hx8gIMbmiYYifW
W/Pc0CX9RflmCodrgQVX+5rLbRyevMRPGOnrfSMUF5DsCbHrA6WFgrEolAcpldEy9d+KESQ80Rg9
H3thbiY6Xf0ZmZYHuuEi6fnlm2HSb4cUZ0n7pl0LWrvH69lhp1+jH6DOAdg3naSYSRskjPHViwiU
1rrcTRyal1SHthHChF3PXu123ozyNq6KY/o8CHQK04tJo4ohD1PQ2PvLohf2cnel2cy/gdpTdEB9
ywR12mqt0dMsmvXzALauEqUPtlx7zRZl6HHZWv3MUF1mZnyqWRctfZRa3r3LyNS16CwWhl1dbo6x
hjaWHIGb81LU03c9G/gPK5faflf1gSnISvyZVfCNPAEqCcbF63VP4jqJFYEDqdv2W4J8oyrDskll
ywL3snXgFS0LoYBg1llDx0H2tW5+rpe6+MN3+p/tGWvR+WNTwoiWBC1sFhIgCL+6SrbMLqZYybgh
myQlMGnyAh2Byw9qHtK0ltXKiqD6GZCkbYIA8SxXeCPwjFwWOT6aStzgzcQ/lFQVcwBF9SpkYqoE
r0OIE1jUFIiWs8fOToXlk3SZUzhwd2x3FPY5OQ1A2pFyhv1Sh0BkPBp0W8ouQdoOOMp1PxQ9MD1v
2toe7/f3CDS8k305KwibjQWg2LcB8Imz7igjlP+7dkWy0Uo9U6NJ2EOtV07pc3lCHmXiv3GzZzkx
JK8+UjvVGKb5il/hWdbeb7zny1vHz7VfD3cPaQwhweokGCsYfH5EoTtXbXjXNvWxYe9OVjUrfLwB
U4PGj6KTnRepgWv0BZufYDU0BP/DW7EejpjVLCECt8COCfIusWw66LSFERsBQtM2uRm4OuVd1nJu
RNQjpqF3RyKZW3KOOUXm1uuz6ppkyHwUI29bmWSacLzHz7AcNGJG3AD/JBmG7DK3T4O6PnZV7h/e
iU8P7dGxiDtmcvo4gPEEPPFCCIwwjh2RIp4+GThAieArtD9/LRjjGZqx+yQcPj26FgVFD6Xcz8OM
fRl/WQ8qVNG3Afhs0AIt2hOn4r8A3Wq0JG3osfPn+EBeHqrBOdNBVF/zpso81yk16/wc9VCvn9qF
DiYkvrVt0D2NxGivRz8ORzemTi5J+pR48o4rm9VThCQ6nJizfpt9fUwaifmdfw2aWiFoIfbEkpdU
OYotvvZC2B5Scv/WH8vmoYd6I8WpTF9QgwRcVMTH8/W/NUbEwtimkqXvuOso2mEmkHT63pVBgZek
TldG50Dh937ZGjUrh99/10aAt3tX4Di1TnvQ2kO9l7PCGffhznw5L3uBuiugkOF4IOqH+xSGcPzC
mmQYHA4DiGkjLqPka4f0QSNH0IMp9rDi9czL5VKJmqNDcoqkYlKhFSHb4suEZzJH3/oXRPmX5BCy
6bidFv2n69i6ImYefcIPJ0kXk2zeUQ4Hdd05CmB6H3BWRz7Fq5rdSH54ixhA8M3dYzJmhWJjVyIi
VICxvEY4SYZkHSEjjUHR2JxCmtkQz/O/gSF60/f0sbbGeHFy06N6QJ4kv6IZx1hUX7l4GyWp+89Y
5tGooSxXd2FqOsXoOkwqPpgoj5RqrTszgee2LIlmqkyLn9xy3Wf4iO39kpiJZ24HuOLw13/C4Lpp
ZdRu3gNx0NQf6qAbzYlP1DP4VAovzQDE5tTGpEXydGxDtr+E4FcO8vYg6ySBwfSy7dsVd1yG8Dzj
K/bFmIK57t6lsouaLcd2sQhcXsbkabu4MzsVGOOhpKZoYgCuV8+c2wQF5DY2i1M4nbSYYybo/JZF
aayyrNsLazPxWkbJMS3Wyaum/xdiF3SHDwMdVmePZYZr7Z3DfjHNl/9aAgSNWKnWpkOWBIynby/V
DgzYpXkQM2tRp4c7uUlmzYCeUyum3U9RuUKd1x230RCNM5Tc+IMUr+YWvGU8Xnc1QN79O0DZeb8s
Es369sxZhRzCHknGaTiOnUcyrOHR+4cx4Z/uFcNkyC8NY5jHwwtFOBxNwZYcSNhX1e0UE4sqlQRB
HNZDcxi7/7NlCZWzw9CVyYNaAQJudlAISp+eKrjMhf7wXdqZo2gm8bU6gEdUpCqkiBm6PE3u9vwx
HAZThMmhZh126yTV+hEnqEbwio2SzNlLOol9rqmgMKb5ewhyZh9hVCiysQDJceHbehGVmO8GTbaC
qTMbrJWu+gMCJBMrmWQ4ccMdBZXUPJGRbPUMgxeFVHj1DBuhaT+kGSh/e2eU7SLk0o4/MHQUX6rA
UGwIIojc9mjWGEjRh6zjPfOowlXfEjP3AjTrhBlPzUXvOssE9WXDF8U0v/bOAI2egesy5CbfLGGj
/eQKyVlMwxq1wa7r8EnFLddE7YL+wk3nWdkQzJWu/8at1Z2Tzf87rCnFCVnBszHIOuz3nl9D0R1v
XbQQGuWo505L/w45ENwRkOD3DyWGBc/kGnaxGvyzt/APn2VhG1BnfO/g9sDFmjm8dNL9kPSgDUW2
Sg9I+ob2Tp/Xth4beDUYYWDYwIiDl6gVF2xucjcjJSOVkqnU34XKH/Vf/ReBqfDVNITNaJG+H2rb
jCcei57abebyKY0IInno0AxPdLP39frTlbQCpeD7Y2LsPNvGuxhvFckByNm7NmovR/F1OSwqlgf8
aDZ0h0CAKCkZcLtyNp5f5Kp0jDXvZCM/rRNOdXnt5l4OIE3k2jaEadqjLoqlxNbr+wFnpoBmKqqw
jD6kJyYF3REqF/4Q5MRKsmQXft7KwL4Jte7gPSFQxcfX5Vw8BNMG4A8cSAHvBgZvel47UgC/0peT
BGV9YMiy3/jiIqTbGw9zgqMNkV+UusWiJKx/6ba9kEMTq4m0Ei3LqnsaXEcswm3SD1cOTUnKqZoT
6aO54n0qEEyunuP39I5KUwXmYV0GpFOS2XwLcMXD1exK1RZ7m/DbWSiiGLqJ8BLSDiQ59zraeBmP
wCjUOlTfxHy0bwU9RGlqYPieN5dNw43kPLEAhhp5j/0NII6wxX8cxfWGxpThe5ghVtmIk8ZrYcNl
hQvP0xLpoeHRrUQmLFmE6W3ruGPBEyQ4+q6GAe8xNdt5X3FBzKhX+FP+8sZP0yB8g02W3FBUNdv4
sIboCSJQ0ofWF8CpIYf+gHeNgiukknfHnxrx57SGT8AcH4iGwzRS15meeHr3WYA1QNxHCG8ZIACt
wKplIaizvtvOsplSBKjD6i6XjSvqlqoeOBP5ThR6IkDDR5/RH9toeYGt/Gww5cgGmNhAH+KL0ZQE
ZD2zjPxPD7cw/FZ4xpXye6tiR5M8hjea8YvM16MAdUdzSQH8A87wU58wiFBPo2fPf8YcLmJT4FnU
K41rX0LIzWJ+iREWjYxRxlN+C7qqyyoxOsll+0P9NEkyQfoh4/jTjiox6YwXqajqNuKmiUYTK1s2
4/bO1UEPjNa4qrJawbpsJqyv2i6o+jSLHkje0G4QHAqrl1s9NSO/32+oR8ta0kUwbxwG5wHMnfTf
1yqeFhJiHgP1QOuCrdbnCFY2ju3ro8W+5t+r0UdtI7XI9MzeTf7Qzjre9wiO8XavUGf9qQRPHGyS
SboSJV4hl+/9EHXg107NiXImfXFW+JVAlaZ4B4CQisxGqxrh5KgBRhFOnrclCgtZNDowHPypFb4F
uw7+l/hf0hYNy9EV3FljZ9vzCTq0lHIHnZbCL98uJKEQwhlhbZ2AwOIEk0X3azaY22fxUvT8caJu
6DxiTOhmTJITIzBoSfLtVuQFfjeO6VeXA9jELb8OFSwqLXhGL38Nn1w4PulVYAVkNt6LlMbQYuG7
u43qe3STBGRiBHVwxJeOOWdEKBaAHxS1Hf0twe2zCvreBcdllhkFcKE4v7EeI+0ldO/tv1MJMOMZ
yVstLpIoBoCCOFHSBifwEmwKUoBazVwK08asF+2DIoDNm4gsBUEWOtTeLLU60JPMwz6eF8f9F+Jm
htI01/xksBqMazOKRQa3XmNP9poiH2lVAtebI676sVKjGrqjSURubmc4sk7XVyrSPgbKYBDoR0Dc
6o2u/iL+S71lFd9qoTG1JoKt0TzXSDWRI6igzX7DuQxdrrQhW7M25phkBRdWDBPU9yEqbNB2xvQL
N6hzT27P+oHOGLSoryenTgoKXXeezSDGAzPLS/i4qF976I7z5oQ2EvpNY/cKErGOIhR6WY6eVahx
LNFJtABzso2/F3AddbxZHocoys7DF+SbIRENVgyL6pN7IhaXp6UCOs+Eff5GMfH5G6Ab4i5qCtzj
SuxGIIpkOhS85INGvvLe1r1RMLUkjIIXeHTFnt6r3T6CUyAw+HhBOKjuf+BBzHFDIGprEmm1uW57
TBzakstSobTRR8tNBY8FRzw7YY3BUVQgbJowSbT7o29nULa5K2g8FYCAOEOKK1ZTiM0oG+3UZvxZ
7cXtpcmgZ7mBxl5cu8oseaAdJcMqbzt67Bv0+NONxi8Zjo41lKWtBHm25PkDo7gL6xwYC/0Xx7vG
0f4BBzR6JXgvabnBtQTPjy3h41NEG0osIwzp2jfRO07iawIgazA5TchmlOIUMTQh3BYMH7/MJDXP
0cw/LgyPuCuVPqGVzVXUEnx1xHBNwNCm81w76Y0kyE5HhDR8mMf7zVW7/LvEyrXWw7YmzJPW658Y
UpME6ssv+7adHp0zO5oeRPRk6g1EnBaPKpNRgCdne+5CEvYLnalxb6396tjw7e8HPsvC+OQ2EFFC
mMPd7iwHpwXuFxIdnrP4BKsRlst/Uhg2J3ed+lHQ3WVLm5dpL/g2+gjdrz1vcGC67vkaYBEXtCyG
iqCwsIXLgXEAhPNSxuq+eaH9bh8B+LNGwlDqpVFmJ6OTriEQ/YWmqw+zyMigKnUH7P8XtoSCv1yg
mB4ULrjyLqBGNmJriYWPProQgphWT+yZYgzDn5LvXda0oWU48dTpGudhkni9+Va4HlgOaRi9BuJy
+sVn8hB14jq3v4d0+zqg3TVcCRaQ9pyFOGtYfqydBbF+i0UPR693Akz2Lt6rmLHTFseJClet+dST
7Dv2Q/U37j2OZv7h2yANFNS1ZQFQKWunaZr0/6a0TVfzTylK0vl3oT67xFaYTBLHvO9uo5yS8URf
4d/ONSid5nIVjItnVE+CHIzsK5NdknRja6y/TtFwY7g/KcCmDFZ87gJrqT8McprX3gYNp68O+PI4
QFCxjk/yvxs51bPjW0WXO8VZY43yazEV/fr1+qYJaQJIEQ4s0U9bVBeR7ceYz1mBc1JEFdDZSdKY
rBqp8q81pRoz5wgPhzhccjpAYkS3h0UsmM96cZ0INd93Ha+1kbFzFjbTxWw4FQevqk/atzWrF5fz
V0LRtHHsTDL7c68Mm5wVxAd0bcnKbiqrur/k0iDVyFmU8RAcM0CvWxnQBSyxCo504nmMQzvQtwtl
NadSqh0Gqv7dX8E3NZFJn/xQICTG3hm4x+3phzgJp+SZi+nFKEcLlPGCIC4zHwFf6P9mqsy8CBPX
ltHshfMrlWHQee5DJcFrrUs5R17Kh8vACu0boM/z2R6/TGigQ6v6mq/nCtsLpXQF43UXi4skg52c
SwgSHDao7m4hTGRxbto3z8uDIxMJ/zenQjz6n/ps2HViWjznZutFAwDBAXhlIinaQYBeVywgxNC2
m0CBF47OT/JaL4kDyzC7U9o2mFc7lv6FRb3so7+37qhKds7AScX5RwmFaYQ25BFbeRgFVtEBp1kY
w0pnUz2BfrwMQN0epsxfmLulZoeFWbN0qmudFdl/sL+dNiqi3KRHBpKXiPscYqkRJO/Niw1h3cUP
NbdOxFROlQ4Cnqh9rWRSnTliN02XiPOd55XQV72lDdRS/uvIQX5NfXhMgL1N12drw2jrYCJNJy9O
2RzZmBfRFaut65mbPd09bAVRcmXS6JkiUAVokSNP882AE4O0ZPsm0BcWYbzn8sd+MOCd5AgH/c96
7JLaZ9G/Glh/sYNfwvyotWJqweuKh2g5mXjngGso9J9JLbmXdjCioqQiW2T1647YA5H075pFZHRs
DWj0BLjCFjmb21/124JX3pDGoHYi6jA4IdparOp/0w8WOs5wFfPoz45x+/e4UsqPJgWTXm9kcCAP
gCCy+5IzEg6daYS/ANgaYDccdEGGtVJQB1emS7/icuD5BPIiVQWfKlTR1yYGI1Ag34XgSV0z+s0n
MMdR79Ys/IkQQyfnDWNRIG+0Xg9WzRTxGfUepNNBMXSGrkzc8LQPrWX/H9H1vVGEGW5ssVh7wf6F
h8ApMNNidkBK3x/Qgfd7zeCC8V106CK/wYTHYIzIw/CXohf6OpvsgxO9XoXb9olXc5OjCL0Fhzd3
2xRLKZMXnsITSoE95Vsu/kAoBhazMYuSuqGCb/akQYst2wD5briMDk9rMhp/pJ32SkRcXJ2MBneE
gzx6P1FDRPQ+ufRWiJEBeH++xsighZ26BZ0/ThHwfAOjPUD1oIz0fSZFso9+2+8iejZ332alhMg0
smtJM+w4wZkFYgegewavsBf7FoHgJcwEdyTi46RhaFjVWsplePzdWe0RKVFNihwl27eqRlJnfHip
8B8P1Hg/3MOYjKtJ+u/TuAA1wjMX7diGqxmFYGtpL28UqYe9vQ5v+j7gMLFARhOSa/7wwIjlCtJ8
kpmURgdIfo1ooTxH5N9R2K2F/xDfXZLbnNN8vEac13YiZH+I6h5FFCej1pnb2jZzpxohM5Kb5IfV
euUgl60teVsGfRffHY7Ko6ffcEMEEB1XqOTdOyvxKmdgFAIrGBqvNmYKfnMtReKttVOJ1OaSp6Fc
c4c330LXDNVh8Lb33Cq7A5ejneHIsvLKDlGFHGr2pwYeHR7/iKzo1fgMiChccO63jKH1FwJo9RcI
AV7R0YuIxY4WlQeP8bv7N5cg/QkFOc0HTvUSwwR0zO3eRx3bOX6FGCqVtrnCW7CAkvWax9MT/SOj
uOfF3y0XLC3weQ+OROEvOigUL7txE651ONu4UtvF2k4CJ97mjBB7N/uIAjbFfVIVse1of2rUdfwg
sXgf4go+0QYICReVqJzPkzaCXsY38Ie60N1vBgCrpAbK6m9ktmYw2kkfPAyjlccMLjY5Mxm5W+gR
NCWzA7z5nVuo8549ZtbU52Na+b5J5+BnhLQnJo0c6N1nPttDO16BER2TYW5FvCV/JipzyDyiddT5
bYm/6DbdJN/N9X+xj4LNi92cwtQZxKX6LPlvonsS4l3sQ6OHCnqB4eHyTqAMptzSs+8KlALbO/eT
4MN+1NbDHt360uE9Kmtr49zvjGQDkkoNTbj3pzAAfE5BrY9xYY/VqIUtH+Oruwj/bb4GWKVWP/0t
srG5j6PvB7GtmPPs6Cr901hkZSTB1k4MAOXRiZfiN3L262DbpF0KGmoN7Y53hSQuZqojAuainJf+
USvYNuUFUc/bAj9XBy7ICQULHa0cGTl4otM8aJV7s6R6oAtS1DUoshoVwqNWPJSykAd6RuzkYwvH
wJ4GZ8H5mHxOaG08w7wsutR5HRmBPoAD2HfnscjVQQO4w4I2pSILfAPkzV4nnvyhsNEAEKoPNt7j
HO6PtBGsJUW7pV9nE9OAuVjTmF3ZTzo54nSs4R2mSMyPy5l9PvPEOngoL1L6sOUncd1OMl/Drqbh
xgKXPj6Ebzl/8Svhd93taIIhq2s2w2ev80t9csrkfyefQrL/3xlJ1FNZOtsgujSY/D29VB3HBtIl
+tcQG2XPwxLQ7YyIC6gnssxlAPpnSCVFdTALJwPEn1z4zpMb6NP4f8c+Ub8yYr7sQ53JmmsnyEhH
TSKKHWndHjDvhHG/osgbVDNySIJMQpxTzM3nz3jzUI/mviQqBCVJHzryFj1tnEWMc9ryoBUr8iXP
5SKvFiP6qeAwaJPpqOIw+iGB9km16p0VGTTPoeLllBfboUOBDgPrLQT+JGE+J/xkkn5PpeNLhgQQ
WoOBYnxMBGwCLdO+R5yAkWggjKS3dFLC9MUK/2G8IA1QYeTvO0tLKf1yd7dUoKJQdnADcqnBb8C6
5KemNuabltXKP5ifbRNANRpTxNA/iijnKq3i8wIdG4bYgHraI/lJwGXeBmMwk+i7MMTcTZTCeOY5
v4dDIbRXIPMT4iVuBFq4w9/fGQ6zW4dreEbBJ8lUVcQSM3OB48Hg/fYXk5EVC+0dY6l7OU1lfFqE
mInEA4z5Dvh+y316g6k463wfvWZYtYRw/Wrkr3kW4FQa+PBp9Qur1FBu3uaBpJWKT6arQx1gHUfS
Xsrf/4Z44IUC7UfeL630A5OtCwELEjZF9JuXWZDqB1fDHp2YffbvlRB70zHwlH/YSItTKoPAXsNi
5w3crVaPwKeIW+QBuUyYGQgovcZtoPmIltHsUMCkgOgELHFeFwQwrB2S8x8Gl65cbB0HD/4iYEc6
P82UE9GzEO0sfdeHpJDthG5Yhom5jB3vBNJ9LXTxUrqZBK07BxaPQCYMVYqQ51VmFszA74xI6Mv+
aSlpi0auOgrIIGKuzVwO20o8TMIH2lgiRzEygUgcw7u00OzG5RSGdUP2X3rkcNGrQagQrW+Qe3R5
7GbYgrvZw0krCooZknrmfURqjv57UmEwr2h2+0CMuJv+4i9OfDV2XLTgAQfTY5lRnwtACJaZOvCo
ymCdnhOYehOBSiT2IoljaWa0spHFPuRUCWullKG4yEbbacmtT2VP+iHLmMQUjJSfNcFw7N9dz1ie
tG/BEll8O2MbJGNne0qKJdPyh2m/X/gCdkV87xYmpG1g4W1J7B4eeJSNAFS4dGR4SCVMRQLsBgFX
CxnQiQc5d4xBPAdsI3yy88w8uAAtOt3hsd5e9U46cp6gzZzYb8hp0P2ZpVM4UkEiijDxnhxLThf6
OgApwe1W305xL42vRTdbASk9X5LOaO0L8NG5kSrE8m1WENsgfRaaKiRmYge8orAFzCoUNhjbbxfX
0Yhn3XZKmJL4wIo7DXpIq4RI696yY+Ry6M/U4FWbTmSMTMK4nBY2wrSpFmtfZf1AGScOUZp+Zyzu
d78CAcyQpWLUGJHRtI17k+uGAmPMqpB2JIxQ1DQMu2anrj/hXkXLc0jwiKFn9MDs2kM4/Rw4D9zT
cd0VJJVJvdOujCXHlXLxMHL51V/zFYY8nrcR+IRlBIjD6MtdWaobQ9U1mDloPkua74V0bXAH+DUT
JnewYDeiFkqANrfOYlbTDKxTixZFPLwUiXef2YJ+FV0bFdwjl/1GlGohyzanT07Ey0NwBHSQa2i0
msUgblW2ZqNvA6Vgvy/xr460J4VdzEOD0pGavUaaQUQC1ybDhHgfCgwZ0zW3ESxqoxNCmM457EWN
QZ3NLdcXdoMTaWyLhDDTW48rXNg4M4zQ2X+FIofWCKp5R7W+k5yrW75w+Ftzx39WZb9lelg+npXS
JGlGPIeL320cKfiW8m5FxLVliCeIiQSz1Q3PjQnygU89BtIDB0bbXxKnrsAujTV6zbA51/yjLcNA
mlNi/2CCfxpjO3si8x7D33ON0hNObFJGiGplhj5P1BQAXahma/BzSjVmbYiyCI7Q90ql6JjnEriG
0Z2YyfyOz3GVuARF3/cybNQWL3OHw2KD3iKmUJs8tnLkuCpJvAiwCP7pnA79PZL98Tjkmxhpdb/z
8cOnjlDmdt73zqNBjxpTtLfPTjdhr9fS1pgV+6M+KCLmIYTBC4VfMP0uLP+t5E7Gug1vj0U95uQw
MYFZUMyhoxQLVhxG6G5CEZWzA4O8sRYIiKWyareZBUMMiOiyNwj+29YS4Z0ARmhMEC8SVuWlLqsT
CCtoTRgTWYsb98LLFZ917dri5T3i7F/FDgi4PkmWhzeJxy+i0BnnMhISakO4s9Qa+mwz0ihEAmMF
zR4zpLI4y9IrLXbPtxEWACqOd/dAzgHxDiQ/EJ1zyA9SYRXhZM0xkhmAe0DMqKs0LIwa25Togqg4
/SUiAAx0DVLej2l3fRXQudIlNbBQhUcisT/gThuKN9Zfh9IsAkJJLaE4EjT+OFuyXbKPqy+Sq4D5
3v/KrdZRJXXqJpLtw+kVQIvWcIlZ/DaG/+xAe/vqszxxsfySDFwa6pXJQ3qZ1bHJJlEO2V5B8fCm
BeGZcormCPZ/VRJ5opgh/8TbJjENV5C0ZQdi+DvO0QaRdSwlBpcExmPiox0OGO/s3iMHeID+fK1f
Biszq0F+53/iFeGFpPWuPSEbIPJY2k3sXMP6d9fBf/uMnTOks7U9MQj4oG6/rpHEnEQxiS/v0Jdb
YCDT6P76Rx2TIPHYCJ4ZMUEGt4v48eJYapav537KQ/zepaT4KyC215+bBTLzaKkOcvoBFPPFMe60
y5KgasYqt4+BrvF2RWzBntenWZfKJ3OuM6PCjOfF+J4Zcw08cr5JsLjUqbYZjxrJmHk7fXAMo3YI
omh5WZK7Xz7oCnkFPPI2mkCizKa4Bpin4UihgtS3/kLnprFLQGS9D5naTo5++qCSSnOuv2cUl5gm
LW15SI/m18Sad4shcFZbH8I9unqL/mhYCJ14jF7ib+PAsCAYQ2moHwfRW11/p+QHodTsBbkoJ2kZ
8R5pwlIIfcAqIjULl3Fn5gWcq6ibpIKNViMZ6SI6X9hBJQmx+/56JkYXAi9Vvzt3AikT3Snsdwcm
ej7Z5pkWFMxN+rxY7eKaAW1NAAZxG0kYEfbJKbon8DG1pQxNTCYqJ4cG9YPP27b0cAsjwXmLhcJc
84li65jQLDNjkbiAA13jgxq/lSv9meyqYDOvhBgfNUdvWOcA+0I9vE12mXnYpsf2FafWds/2ZdhG
cjhYbwy7SkQHoNz6xpOEOABv6Dx/USl3bmZ+ScnTpXJqN3Vl735O756ZfUecvD+kUUWWbvAN9iYk
p+KJAaxzDihbNgYiZACxZvLdsCpqYXfXBJ2ENGA0Itc6iLIr93XDZsSdYPNhjD0dXm4NNZcwwI9b
9qQxJkdMipFTqAQy3aeX1QAeRwYBjk5ViH33jyhcsstnbcw04qmo98KUVlP8p+7u7/LLSgUg7m6z
Z6OVGAk9psMwbOmXu0/kKjbGLJXGkxytLyHtm1CRlDjZmWE88RyxAsg18LxzWOGNPtwlEGNIxq7k
NxMBHMmhXNV0QaEkkAUlAICFp0a7ZfUhM4hwhMH8xZ6VDA0Vo4oUvrjb1uxuKpHgtdjSHupizssB
sUUknlLRs7gjBuV0tVnLBjjLPtBRp+YDAzr5fbhHkLowooEKalX5I4EFCMdOeMQNrstogRaaoB4R
5hMLvBgaLh3MVnoMmEzxVktF5m764Ck+QRp3mqth9U8VRtHGJgjXjprnHC4Kd6kOoURHieUe0h49
dlnfADCml2JYo7W1sGXdUM6+sMCPsXiR4zjrh/S7np3c3uWj5pSAnFpweUCjLWbisk1D9r211TfM
7bkRcdKAdpAL8tiLCMq/+Z66UONZkiXSWBHdizYZbIEG+2QS5CdldTDRIi2s3j7yrb9Evr351qjN
jwN/yZfez5WvN2khTD4w4Q/qoN4VyE+pM+nlQ3XK0QuYgHR5POftSDKNNm0sXOpgTG8DPmuKDmvG
zAE8kywBUUMrClqJCn8HFPi23Dgvztw9FqTTELrXbq+k7GTDFy/I6IODn4QliIR4uqLgLUF6Un9V
qID8N8jmKjlrzC1blM9NVFvwvQktORY3y8aQcQpLG00HA8Le77w+u6OfgWKviSOgp8l4LhbzlRoV
C5RKVyrw0birWeWNwwyA3xnevOB88bend46M/HEmqtMm5mB0I9gjWpSeb+RnOzpyhFBK+0eV3iIx
jofSv0Tva36Q3g7yVjDbe9MtZzEnl5Q/utDu6ptJOnevtQHv4XiS/6RixkQ8/DV/cV4ESoaud04G
+R5a+k9L7PpJAMKmHkl7rw9vzaWdLOSP1ka3ubvPQqeJeLCQD8sCUJx+A9rvVyt4MCBdtV7HlNvP
H9V8MBUcdNLM+jQSXOT1jtsL2U9GGkxKT02RWgzMJitnMHU1m0MfIrQ+ZSG7HHKI+hskDK3fw7/E
2EK8xgjZZTX8m7qF1oQ1/zkSC6diksPbbDsFbnFf/lnBgh9o9vHlx6OWnKE1QXGaQ+W5yoUuKA6j
g9GPQjYew0G+H9ToTCGQB8jE7zpoJcuBO4QAtqlhpa2vvB17cDXgwOjyAKsDbilSTN2cC7QI/593
wxcVAbu4J7guDQao6tkTPG7vgmw+BQCWed/CAZMSfxTSK/sQ/k7+gVdOeUUSJfXin2wBjgezVBh3
GqxrZfkuCXb6dDAHR+51nznCa8RpHQIXxGS2fb/Vvhh4e0uwwJEe5iPK/XCI3fgYw9R7p+7KPbm/
OL9H0LHp69sLWmHXvfnbLFn47uPn2i8tJsqbgTIKkuPy/L1sxBRAaagFP2/p6AbKoCepM7Ublkol
xJAbLIQLR52n0S7ZN0k8ZedqLOUi8oHOYeQhXZsW4APF5pHFfAK/vvBkn+ceFZOZrNDnKuPPz3tP
mUoGGT97UkWWwiS9nWOI36eZBMQLP7o0v46STVO028+6Cd7JXripBC/UVtcO+Wjh/1afn5GR+Aeh
2hZyA/QHn66NRotLht9/wlmYYP0PPJsnZxazHN2q4C9X0T6pszkpfyRmEvhDCAd2Yb7ecOSNrDmK
OKyhzOrB3tNZXdTQ9336YtJ1XtUByIrQD8dN9M7IwTiXxz7q+/BWqcgJHu7xjtuUJlGBucw5t1Qa
NTVja80ndDVrfTyFr/AoNQeNiCzKf2qao+HARrn7x2dhtv+MFm+r19HcOzK2+CUNknQaoH0nQuq8
pDzMwjiIZfDK6mvgsBdDrfmS7tBnR2PbzRsyQbdB194BmdsWD4i7zkrx5kKBvOi53rJBd+QW26np
BJGSYcF59cPaaqeDJZ0BaMqBOIIC9zYl6dD9JusmIvvwnm0BDc+/g98n0NGJ2KG7iYCSJdheV3T1
c8BTbiS1pbK6KI67il8LgoiDfiMy6ai5z/hf6t+chj2huF+h11juUa9rt1u+PCEUConptxnkDai/
IOQfIxkYzm8ZAjqp6IKpHy540/rG2HWtQokyfqunbujhwRmZasPzVWgrOGov4XQ3UHqLtNDtGeAQ
f2dCiKgkH3htE19A+FNpbThozChoVHt8bEbJZLUux4p9awZy+OAsiJ6Ro+YMXybx/kgqYtPlNAY2
VshyIZ4iRfyZZAKw6CGkJ7cTOBQFQlmL4P7uzrzB/HdEZ9Ft+LTa3D/0M7CUEWNBAPgiWbGjPCV0
moddu8pvuM58+NETLtzq5rFrNX3mV05o+c9YHM0MD5C3SKi6oQ2wa5tf8PyAMlIcHlgwKQ/DNldC
e80Ild8acZ3fR6lwpG7xNmRXGWlXxknqIcKw5XGp02JlAXkleT20IS4pz81Hjo0pXvG3fN/e5w59
EjArKiXgUdLkP+UeW74AXDo2DRu9sgxvGb77wMEtcA+xsIH+6Br8bHFy+TnQfF1v1IVdTmcQBO2b
yR5MQdLd9iej+OrKSWoV3YesFDeXgRMZ9dtm4FkL+pa3nKqdtroYtBRlsSzpMxCtjuCElmlNVber
J+dnWjIFhp6V/NHXQmGKlJGGeBKobRK1K8g7rvGb8NiR/AyjWlaA+VlDtV4u2BfyMfSafCxiqE/f
rmXpLI+ST1VMZB0yERQ4eOtkLbsMq+ebq+Kqe+dHRlT4uSt19hSX+LbvL3LJWsjA1aKNFdNygiAQ
txUpx3nQ9+DE+5T0tO9Yfpzbub+Ev/si5dBL9sTnrpzLGXyg58a3zHo0CTTFsFCFrtq6vC0CuCcQ
UOgxODcY2dlCVgyKtSHMt0TsoEMl0xXkYRWrCchlbQznC76WxJsu7Uv1R3eceJPeXUW5ATkGgHRg
HjT4HZAivLVH8ED+7RKY/jRn49IppxwYcqX4rTOaWjYpooU+v1A+EIi+6y2w96IlQQARxvQQIr+y
xBES4SS4mE7/r168IJK5c9Ct8Grut1wSrNenQdoLyWjjwajkzUNQSBTrWSvHtwgSs/n9GCCtMwVR
yWMl2DljRVfUyAc1Tgsz+tvYl2wXxoVboVgJ4/4j8I14gvrhxh37x/lndPeFgNXiJKqhDYDsdCvK
eBSMZXteXlW2EutdTs+X73VUsny74i8pi6FsKNJUecR1qEzIzbvMyWR5j2Fzb0Zk+8rkE4kevD6s
KS83eCDj1Ao0eUTEKZH6WwR1V+w+Tbp4JFIK9gSu5iUtk1DpB8BJpcIMtohqwdmSLbzSRgT+x6K2
TSq0aVwKncwwXENojJVhRogL3udvfO+pGPWGCIf2ssdtj6ZUvLI7c10EK1mtU7NPe8Ki29myVufZ
G66AmWKkk7W+nPclczrwvMJ+krXnWYEI2/zLpg7VG6R9CkrDkBmGrOQOIDmcp0iSP8u2RFYarq7c
y57HN0BCF9C1ab+LPaEMu3u2DWluDhnaZcvyxoPfPzYWL4AILsBbDhdWJhdQxmcH7ra7wTIgIR+2
Q1DkjkFDLYQ4IPqbajRse1xYz5IkxW9WGvfAFXxENiq2ff7EkshSsKHVKJtX6kya/MHUk9dBPutO
dPcWjIBtPnk5Th//ZGcIO38wTMEEXdc/6DJliHTsWpJwfSFtH72iNrlgPRoWxC/ueurDpCDWCENL
LgYZOxBoF/O/2zLUAq4jw52DhsBGbfthJei69L5N+4kIpWqsnMELsfIlT376a7B2a43MO21fCO9Y
xwPH/M7sQtoGuFSYULYN2vJRZ5SqHg1CSobMb8+tnPiQUtvN5/AeLwlBVqHrFl3TTzvyeUhm87kY
nSlQ2aQQGhe+2KBXNono774GIp0dw0p8MvRRm84nJENqNEJR89GIT/B80/PHMe2uuaR9HSq0BFny
M7RScgPHVHnbo3HNt+RUTpShb38hcb2JhYwAxiMRrFxUgT/B24rSsKsSzzcuOUPY16Qfysuj+eQS
REwkXeeyaMgYz+g5kVJoKdSRicp/cXkqZvJaM7G7CfQUTdJjuC/vdhUAyX8oDPy/z0TAvij7hzLB
i3JUjtEMFbdR22MvOl4/TuqB7sLQt8TOjLr138eAZC24x0A6AoOU/VhqEpeCf1hoY96c5STXdEtb
fs7FffEnehir69fNeI3h34ScqYps9QYvIj9itoRVcOHFCtG9fU3FxdNICmJn9KJB7JHpk91xopZ7
ZEvO0z6k8bop5Hy5wlVjQZzDIbJ0RwIOj4UtNcKa1kdDFJhUlyuCjDYdwmdzkhbwl2GucZ0MmsCg
dBTrmOJoWPLh9mK8Tby3y4DVeNbIX4TQn0eJu1QR+klTSkMjyFjcOaaGYU5I5DQVa1QYjAW+twsN
Ncx8/AXt5is/htrQQoXKljsujGmi/bW3orAZq1pfehqi4ltnnbjRFaL4e6l4Ykb5R5iptdMZ4X4c
M1nn4w79skifk/baxw51XRQxQvzNT1SzTM7KLnzgeAs8vFOb0vci8LGLWj74KsmIu/uuDuMmGrV7
hDx4PyMluTKldniY+kABCW8PoAd2D1pfzX6eAwfhY8KuvDKaNlp480kSmY9lK8GmJF3TDBNt5XNF
szg/4dAdOiAYy3q0CfW0y9pWvMNqtTeTsByETeVBTEKP5VdorMmJbTuqcVG1YHRhng4BaNmUKOHB
9O7mavdcPEgtehU0ff90P+9ggAGdeLT320wfiUOvY3EO8xizq68A9DSeW7eI18Ffc4XEPWGd0ZOJ
/4S6IDlErFobUVJ3j+beRkvO7gPsutnWchixNElK+Mmj89Mk6D/gtiA3g4Aj9jpdpAk8xQGoNXe0
NTmeCPR4SwLEFq+KHYFD66H7dK8Xax6JtfMeYLnk+poPsO9COEPl09YszHmHNBCAyWqFnh4K+Uv1
ERtyakZSWTZv68tR6CbaySvjr0gQr/3cIr5/KFOixpsxVn0cgukbOj9iq5Ygo+qszGxw+MTPNt3i
T9fic38ghrRJzEdEKnpaebYbQwQG+ulDTDRDvTyV5qTPlsUzIOUOdeYyng6NEbMzrZneMw0rGpYe
3fafxlWBRxbBmJtylTR0gl/AezCb0qcnRjYJFAmd904tvILOfXBdZDaz3AP1WUsJD0mt7DldXiIp
AZguNPaJkDaLruQyUbQOiT4/jQnzTdITbrt4BgEiYxjUkJpd8UrM5gx9W6fMeSjumh+Cbfh1YLcH
y1Y2VO32n2pkfHUByZXnmZhsq/mYCBBHMD9Jo6bB11jbylZuyPo5OHVqdzyFyU0O5yEPYBNiWi3Q
Zsy/JwGbB+9PnjvEXzxBT0nZWSD6egJY22RM9bJZMkboFlCFI3jlj2nDsBrif7nJyP3LvDIm/s/Z
p2E+7IgubN9obE5RIRxDNg2rEaIRLsL6WRrg0nGn8CPzd5Tki/+aGUce0d2TICZWswFgpbgpSWlK
oR0+ulATD33X/qKKPtzgG5o5EJBaiXKtV959BfsaA7wNpssSZX4aowC2DZa4Azwarlo2+iB7dY+6
YCkez2PeBDIydwC/XLLzjrY7ABOMJZRiDmD2uuCmHbXfibCoQjwenat/znVLtrDhEUsVj6LpIEMM
PnMl6w/jwDkJhpWAYBnseXP6YT9T2MZ1CSFqVUBj2NuBs5GPy3dIOU5DqZX3Ro9rlLt/ACdaUzXO
dvZW1Gs5D0JXmkbjuqU95nNeiaHMQDFnghWGb5BAmrdyLV7rVBuatK908z0BtAKnmWCDOzGmpSm1
2fm0sRRutvnteRvRSsb1CLefnk1mb5pS5Heq4DnpqjpXHFm1Dvb4PM6ZYmP9TOXBA5EGVTECAqcZ
ovLPIPeKlOF5/wc2xcYyeQNmxMCKAhpPN2hAYyR+Ej0yP5A7WWiZ2KWzNHqTX03SVa9N0szTNSAy
Dg54A8oXQoeMUsGCRW/QzTQ77VPRpRbmuFlJyZX+w2IJjEQjBbtST6h9+a6hdaHMn9fqc20nstlm
B1DD0ww9DAP9VB1EvmSmAvcvrX8LaUHFSqznR3KQqlZhVZsT2LKU8hZ22c0ThyawrGxj8iZJWU3v
q1BhXXnVMd59x9bLinMehf1J7ZzrHaVEuJ7ICPYD9dQzsnQzsFAm3RzFT3syw3q575slEsx1uU/c
59hj+f6gVCqnD0poOhIHavxfFGCzgb5ZYjTG9ifvF9jDSvzq+G2OWbhMnErWjQxi8bx1wPQGF996
Ovg4HqIBrZ+Cm9mmcrxUKG+pFTEP37dPoEAmnVKgT6379j8lixUiElfIvzILjq8il/xTeCeQCkRC
R4Fk4y2s+/oINFTdRnmI4t+9rBpaMXXz7SxOL22bz+iTz/Y2pAMEwI4227pUJoMLJ9yqrsHbFmfD
61b3FeR9qUbp9ZCbQTIeGJlXjdBhvtDhu/nB2VOqsAZJJNHflleh4LI2QpoTpcWaM2gcPNki+dJQ
gl+CAerw9JNdWkljeXS+47P5tlXqfdj6cUJImGrWA76tsWwxYIzkE9yj5qKK417sL5vP6JJ+nTVb
w8vy+BzFV0q8+OTfX6d/BUwGCK84m4AV12GAQu5sz+JJ93/sTCrNn8O5PlP1plgiUOzTGeu5Yx5b
n6XChqqyxOqV+rD9Po3dZJCphJld3DC16P+YFne73rgpSINERe6fdHw2wyNVHdztPJyiKwZ75ba4
T042BZTA0Vm9cvrTd4/6H28yuEXLDbVpP9SOOt3X1G5DcwNz5eUtlmxo4Nziqja4aAso1KlbUWxU
QJyUKXqhq1KBuWcuDGEm/yNFZQlPeKXkjrvN9gxD/G+s1qGcK4kVNUh9pGnYfYsWU3EnO+MXkKyQ
cpW8Lwxf2mOpeMiKfiE92KN0W/PDZ8ry74b1UMX0lMoZ0dPlddL06rqQY595awyPKi3ObQQjgg0S
z9gjdnoy52RdkKL1MNGW24owX1ri0GTHZsz3ag3VVcI/jA1vJFZUb+qBRqm7KOelC1pOeuuJH4II
yYW6kVZWEBWzfwBXRKU+yTwZOKZfipUIi+dGMjbMXhCZ/7tjwqtrz9xwHPWIyChyqXDiM8lJxEu8
xiiEVRi61H5nhxQPhe+i51mN990si3DxMAyDEu4gWLYqD/gIMzPTacCLPxw3G2VNQ7x0bSy5aluN
3Yi689LUQLT2CjnqSqbV9VwZrTjeuCmIe7rnVgxDnOw6iBgPvxQB7QYMTHeXB+bE5EyY4odjXgAF
N4G8YkTDrrcJNMKsP/Eg2WWRFqSIa8E6l+y+QickarjPZhhj8YhhPbyIYOHafirr8AjkvVCNSkhj
MtFTXipuj7W9sEqYCNxQtqfCSYX/+6UAp0r/LFpom1lNnHrX530QaTVascAKm7gmOG2u26nsHUhh
AqUNHnsvhwP4YaYijm5n4fovZ2m47uSC3TKJSnobeaEHJlx8hgrNSZaOgwxI2WEy/mHSxWhDxfdU
TtNXwAH1v/Zb/rX5nLph7B5T4RINrUY2xKzhBPhr13Rwl2GEXk+rcU78i3PhWr2UD3xg0WETIcwq
ioQigtd1PxpNeHRTOJaOIGxNk0qIKIamR1syzO7Ocu81riZ1pjF1L/w3f3gpOorHW8+tPQkmIlT/
Jx1yscqX3C8z8gzJurqGImcwYgWs2jMZesky+Qq90gkfvyWsISXRDhId1NK6daicNBeZCtBvuPHv
WLBAKlypki4Y6ROFmNJP1YMM90Ql2aoXUxw9FMwF0GzEUZCKV2giGHXXI8Kk98daAVNTwuGVnrhq
wM3MDTzf2w5jS3PHTSNxWTGk27qnTEFJPa/Ijn65nYwEokyXeCQ/XVahpR1nkKi28hqWe6EBNEp5
4IMNB0T4l3UU3Z6kGsjgBrCxcrM6PgtJcELTFDj5qwFZBhcujpqTrhW7W6PzZ0itt5Ujh+eh+O37
Qppk9EGkyvz/M2KGdJdDBOd56rgq9qF8MBix7aYbGk5KW0fNbFwm8NLxKWPRQXwQbJdedOLYxber
/PGcGk2tYOT+xsj+rTSZn5Yh7YfPaMpjWSMzfTK1TU8crE+Rn5BjFYxlQFrKeU082kLUsT6OQDXF
6qyVNpMHBWNnTl73WxCuUR0IB91+quFMYAbIE1mpTJDBymM7WnYnt7V00twsidIpnaaCB5GBZk/z
vx3Adk6SFU64JayD2YyLGlJQohU6mdt0jQuN9QTY2XGjJ97gUFAN31hYsDDMqFWjZcS1+On0rjy+
mP3z1iT2VhUjtzYTUL01ltYr7J1mcYOKo7SwCZcb3r7mO8W/bV4FYmymArGvSRKTJch6HdUf5vxu
4MJByo/9esoGh5DYhkbkNOUTebXoSGxksee1c0QAiOwtOA7g40a5F2jVc2zCPRZHHYOdTPOq/2RZ
XQYy1lzn+mIr5/zkyu1ZUZy27pdLCcbBKcW0Mhfb0MH1EoaxvdC18s3AS8BrS11lxmA20hf1O4SR
rfbOJIQliv4OHaRKIRAG3fx76PAjeKDohhIersxds3cuHsvTr09YkpKz2XTt0gZxWzjCiQA4iwuL
7kHn3aA0uFuWiU2L/14YNcbJqzk6ppuh2kwKNl4GtPt71NQ9h7HagS/5oj/GoTE9AxPxSVT1Lshl
Kq3WimW0enqI+QBNGwrBOONA+t8AW1IuMs+MQw6nP1qgoKLXdFSMz3D47hlf/XzGSuq+YGb8xGWQ
4LMehB0CiHLTXoFUM5BpDIi1cHHrUI3MooyKvXdZo8azDwPhX2DKR0CBLI11On6YaFd9Ot2Qlc3b
gzyH/fQObWdxRG8nLF0g6CEsN/v+FHNiS/uzeYgJ+LD5zq5vJQ+IcpnAlRP2S2RBYCnq4z/TySri
iiYYDbAm9u+3rlU/SeT7R4zrfJZbQnBd1Bw+VSS9y8JOzbpRRq62rIoU69W/SfKx6EPYsZJE1cKw
lMS3X0ZeehztITB8/G+bhM325oypqMi46JlgHlmWwoNhnZNS7dYxOiGQZ/P9lbLTI/n0ovlOLl1c
CAA7c+xv6CS0UrBlfgHwWAeNYfWAdMXgcmV8erKCqrjkEiK3cgoJuxl2iEkF3m1uegoIfoEZYnEI
FDuc7gSmFrCpah03zd97dOGJXYo08XirkCVt7g5YdeeQM0gQz3LpTehM/rbHBlPLRT5BfYioNIlh
IN3D08Qf/Yiz53Hsu/wtALKfz8v5IuDfxojMouwAhOuJ1f97sezFh1fkucBJJiA3Cro9GSS/klRD
Qe8g1oX7+z/1rY94XppRCqjHv5XtcI4/ePwXS0JV4xRwasilwEUwf6f6eBWxoZ/8ZBTGI1ZqU4x8
5f/UlZoqV91tCPAKGwmlkJsbZ5UIrvbxbbMhkb0SMSBOwQMgJRBwn4CtHP8vk6k6LnxA2mm8wBIz
bIZr7lq7xp4KJgz2Pmlc3q31QJ26tgn3XT0o6WgC3m/2v2Sf0F4G/LiPMpekGDf6UhUpAyd4mea+
Pf9BJ2ryv9yrCZgSzoYgmPFGvI3vektrG/AGTKMFrJGJSqJsQgdrHduR9RiGrtlHQYx4fg9C87Wc
hx0fTlrgcBBGKqojDjHfec6ZBBnR8QPql0kFKDpdU/TuScxAeUC4iuSC26udAVYeSUG0N8kT4O5l
kF6I5KFkuJMXaXUCRjCPupeNHYyrXO7f8eWSurS7tVSdp8oqm3RSIIAsKeGy7dHwjwH9IDG+Tmjs
k6n4zXfOafwTf1s9oKsHeOGWx2+507BtS/sMTQfWBdIyr7OTOU9to7bp4ov5dj/i3DinLuEP+26y
/duoX1vJXryHsOkDvZijh16sqqaHfrCPf+sRdodmb/OzkAXSzNiXE5boFFVpgGgUaLwmPs6AreAL
WZ4Vv8OaEpWxfyHPGgRPEoqpYaW7wInFwFRcVjoQq2atRzWsuF03O/ZvMpfwSEkdBDpHrrGTPXzR
lNQhXjlNMws3/eVerdrcgwX3j4Q7mLYEGG0mtqa/spWmWjSTB7rvdEM2a8INKjEqspb5X2M908Nm
e4kj4kssuDmBFDezZ2z24MYqozp7S/+88bhAo0hNRaD/O9LjTcXJR4HluYqhCsD9uYsS2VDmSiR/
NtUnYnYFb7ex+IGJDKORPFUDLwyDIhensgY70IFHR86VDeP59YmFSxROqYDu5UrEXjgDVaBydHfT
5DsQ1IuSKCCI3L9jWlNG/4Y0BXbwoNUi2UuJM0XhkDiIDecMFeYBxYe1J9zR+4JzeM7trtTG1Rxb
h2lKOexrKMzbRvdupSRpWU2p3psm1+HMZoHdR2WEugl3iGoUr4zcJfYWGeTcAAEq5Kw8iZ5BSQHx
SGlhQ+8KHLO9khMUwKF6Bax9cSykVidxquYmZStUKu2uCSIQtuXUvOCFPMR1WVqozjRfctedFVp9
bUbG/C/wt973PRwDD1wn8Na0qYKfaL+dOzVCONCVJ9pgHxbOGLXhtKTnHo7VZUSWtteIM+ywV93y
DpnWlq7W2eWOrkYPcF/8RyQzDfacHuQymOgZTyg1VPNX/vXEnArB2qQV5gUgFAGw5xUfe4mbzkC7
ukwh+Mg7iNH98b9QpogW1MQRVhp+h+iWjmNitalDRyU/Fvhpq9mvmRq4SDRC0VBzB4PBimUR1FFL
TWsm7B4dvnpjrXUPv1GB6GJsGSmAVbd+azlATkBkoquprfwEi2Pe7aDrhOStNQDXST3hLurEcppZ
7fZF3fGd7kckqWyY2vvk9Kkvp4QLKj1mIbBIpaSucDfaMrvVeP0Gaj3jYyeuk3RKeDgiZwkTQQXU
g5qGcmE/s4ObIeIUM5FYqUf9PDjb3ZB3o+Cmf3SwSkU3/2ROd1tOBj+mxmhMW4CHS/WZxBTo2jqh
9Vk7R9qwnjkfo0KsZeLVUBcx3hqR9zf1NEE+C5W0nsI4WkNra0J6ZPMe0pfta9qJQucgbB9XcZ5j
FX/7j1SSID5kHziRF8mj1qgkyOiRnhUe0ejMZKxtWLUW1F4dPr02yAylKRvTGor98s09SDhaL9dg
aCQyQxilQCscqUSeA57mWjJzGYpRmM9bGomTnLuVqaIeqx7pbNQ+wDgd/pC+RQGGVutacW2pYIib
dJYGeV1UFAYwCBOmjUcgXRixShvdfDTosHx9HOzSRRj8Zimc3KGCyNiKCFRzF3KtZLKmqCisLN2g
Ut9veb7ta0Wwgw1ATTPH0ks4d3mjUdt87Rc3qKOB/lk3PK2DSQx0EqnQLJ38k0DoSN74eLnF9RSr
5hR5uXt39HdMCy0qx2px2u3YgTaSRssns8kPg3O7EXvjzXrOk2LeuM9G2oYCrk71sJnxvB+qStG1
CuGc8uwbdjYyZ+dUk+QjOU5zyTCAJjyHehcT3zxATEGNZ3qyNaxuTYgM4hjUgxJFBxa+xPVW2Nti
A2GHXOU/lqH7/FI2e2Z06VMHtPBFSPRtMj4hRUCza7xBZLx0Ytcc2pE4WqVKzJXq84tNNH85pbf9
SmhA+Kb7Fo3F4sxdXU3EpbYVlanlgO0kbdzXbEXT8w7CuHBxipVV+YT7tza6Cv75Cj3X6HO49tI/
Clvrjpdr3qyTt+mNy/WMmVcazxZi532DYtnvvWgUe3xgV8vBEZhpdHHUgfohXnoVOQL+LHmEmY8U
R+RVxC5MBYoOQidyj76+684jgB8VgmKsEoFEi62aNf1y6+JETsaXk1W7ovnWTjI9+UaXxlK6Cc/C
6iNGgXnyfu8ecVCAqDvSmbX7p2yJ+tGtiy5jpR24RQ7oyJcsVwom6Z2dt65f9yU6b0lnlmRcibe1
o0IzUH1dQ3HE3WGzpSU2D993DXZHlH7+k7Rw7GocC+Q75IajuHBT0xEsZN/nlStRaCM575e5u3aX
wuFakYYi2SzWa93dparJzaXjVqzjFemXP7dHlDTKQ408+2IfwNZtoxQtzpcBx0sKNwN8hRcOGR6n
YrCqq9cOwSNKCFkmCaxvJmijmGbqeO8guCIqxS9oYpM6AmGaVgZqTVE2VKFaNYLnMEd12lMg8iZL
N886o6L00fMweV/5mHxuQkajm4DKgWYSu3OlnrsH9KtXXNf+5DtSthMwnyx3Z2mWHHLHYUQWZk/T
k62d1oXPLZx5cqT5DoKNFBQLyc//UqwqAQm8sHpKYX1S6R+qmL0AVZz6lV8gZpubWjbeVoj5ZDoK
qH/JdQrdAPrO08hq8H+3UUQ3rcddzKYVroGATSIM/226oQVuULcp6HIgMCldBaKtfZ3uIhm7eoxW
XqcGCmohFdpjod8icHb06oxAho7l4zUdeQziQWc3bYtcZvs8EUWawOdKCtDsrTgEW8qtXTZJc+l5
02edXKf4wa5LOqXZ9wkd6Q77L+nvwCfvnClFj/b8MRVv3YDnC36gTJBnKklIMqFKnTKrJrEingZY
6+6rNaQlMUvy9xFbnywEA3SxaavSzb2gDKo9OWSKDNAoKmV4mS4edy2UX5OCEmltLEwDNVdEEKrb
XK+ArEnyPf9aPwVhWdN61AyHkMVFZDptYvwdBzhbgrUUeSN9xjDHnTpBAY7bIlq+lsTRbXRUhYB+
0lSIC1fRr6YQjIt1YXRfMSgyTqVSnWyKOxaO/mc2ZoCM6SeeD7sSOC8Cj1kmetDPKN9Cnc09TU7v
Z72V+RhwhVjvJu2s1lt01BmV/wGtlEjknEWWpT5tox4udCojGhs7J+hf2m2Yb6ynv5P+nWCA7RvX
u2bEcWFEsUT2UkL8PHGbaexFZX/LSMQc/ZUU3rx9oSwqS9PXkiaZFwOqd5PfG/v6RHbJUiRoH/x/
X4dFTqMCWkcdIttc8/3GIW5TTA4m35ucS44MJwjB3WfOjnij9IwlgwCqHyWk7FCQQpGLBB5GjKYf
cKDedOPzW5rhcCFdk4mizf41g8jHsgM0b7SS13gPc6NGIcCcslKQJSLuELneNR+USdY1nkvmcSAN
75LJIViHMohp0bW9QU/cm9S7FI3ZvOOEOCzhUD9SaVB0XZ7YP9+eGLnzpg7WBDv+vNQq58aTyeIC
Ywr1r0VU3Lcjo40os5P+EWFtTOUevjCHIdwVYOED787Tst4xSgWSNZWHuuyY5pqpy72wsL4fpAck
gFhD76ImTUbmnC0HG86Dq7cI9UWCsZcUWh+zGNtbMUSYISfb2ANnDVIIuggJH++NGqRR6La8CIkv
pF+sSmuvOB1Sfi5H0O7qnk/OMHYM/zYSa9xRzYUzi++nrkDgvgEKuWNIpEKsxjQ31WmOP7rAxJg8
aDS8n7UgEpsv2yIcB3NXzoR3dP4yISh0unvVIR9F5mNeNyVjuxUXQAcSV2ElNaG+wrSnDi9JlOYZ
NcPCreW93WZPTPHBY/pxjzFYwA8Q3zENkVALC4cOL07ib2Pj9g4hhSun9um/2ayZbGgvDNv3bQBV
zVoeCWs8T7fZcljQRiwYrpguoY/CdKT7dJhLybXbq9GHoB8SqRJioiiCtkCCjTRNqJobAeADoCis
mW8xcev+dh1UAlnGEU+2d8cfftq3X9ccygT01dCNkchEdWRWZg0YrTZAcXzX1g7Fq1o5gqNeenfP
OWuJV9NwJytYohtVXgSkyJ8+VcR2NQ4bSJo2WdekZOi5O+BbgDwHp/geYBUco9dWR2JfiEgKPy2e
v1kUMkSJQd3/zTGCR3mvnwA2eBP/1l2ps3Wkgu7ZY4fTXkVjrKal4qo1g7INENxCdsHXY5NBP7s5
BhXdaxoDdZiVDCJz6A5ERGBVDAOZauXcOaOTDv751numg1behPl9uu5X2q3JaXKCmCvbwwiX4B5w
VWgkaEj775HMJClEbRfx+buZv47alRAhIq4eTrcGhA3+KRqbYjxaf8TLPR+2FcTvSTo+4eGGSCco
uIRYqohb0IuoQEMTH7rdWN1U5ZfpyYlzyVAByIedcV1cCV30C26f5rAa5GwQRR0Jysf2dZkfxwQm
nBpt5sDrktAea/H6OdyaMp7po1s+4YxWLIqn8RkYmI+GCYw+Q19NDqRAzoVKusRBbm8QaZCW+Dnu
zHwiIufUiCYFRT0EmrDBveukVfOPMkryN6WvJJGJ78ruqQEgZxT3ST86Q/2gBLDJQEgHb1O2T2XJ
wAPw4teN079wnNi18Wmc/x8t+S45+tLysrI/jnnKu+cv+Ahe23j3L12ZRuWvnVlFk35zv8HMCAwE
HHtxDrUeJ+rM1c2EIOIFLWwkqiCISqROC8zvWnkm5lFuOVgTElC2m4ysdoxjLfyJAuG5QLkV576c
uahftGG3FKjV7olQcFNmID1O5B6FoSN7ABKyHCjciskDDWhkTbXWRPE2VLJvHg1ZzKtGI2DsBa+Y
kFMX9oNjVBSR0Juc0O03gXRkrDPUOZSuLkN739iRs49nQaeEdnFQ6Ww+zFVtcTUEdA/6TlLgF1sk
hKOelY8u/hiIAWPwkOZsYU5i0ZYEsDW2qLKUvC4rxkel1A0XxV0vl7qCa+XlGi5V6JO+iho5/qlc
JEbS2xMeZaYJmwwxA5ERS/fzs2KMCYDll97/83NgPhokXJLBr9CMBah0NNDU+Y2qrX3PeymY0Zec
hz2EjalZptmblUEJ1a4ZnWEOD98M2QMR/13xm6rurpcWB7LJgYorf7rtCwp6NnRh7ldSoTx7g8uw
lCSU5HcTXD2hpPQ4XRHKSdz6WnAkCMu/47/MQidLm7NIsvRBeOZ7zJX7z01r0cwsX2LzfzQDdYH8
xqy06gUwz2vMuINVhJGSl8brp9nj4xOj2rCK3UgH6DqA+s5Wz/eprA5DOmjpWQ6gxKB50L6vdpsL
K/fgeXTDGP8hM3+XURNBUfrt0cz8ShBvXOkrbxZMcNk57/Cki8epJm9WSgA/Lg3Lr6GZ9fTbveAD
BIjvCde+1Nyc/ZQgwAh+xnmSmn7rISUp3BOSAY5napghKRZqegNMz/xj9Z9qvPN/QLOfDdR9V75h
sCA6JjEuMQWwccWzTinZdud/w6aABIbtf6AkdwsG+uVd/WDuyeV5yRrnpLvA2yIeRMU7wJqhYQ2U
ag4eMgTxx9jjyL9Ucu8K5qiQYKA/cIOYMkTg2sNFZUbJtxEpvASjzHA7kpM4AJWUWkaS9ULSre1h
Ip6mK+oPc0LQ0Qpv0JJwszASwtjww0vH1f3kP1H/io6DHSXoyU8rjlEv87Dk5HdQQIma8gFiLEIi
uq4gJY/x4YGFC0X2HiOCenN+5OCPjOrbBwjE1rSORXtP+uRBRFR7c4353G+SLBW/XAmXlRBy+ri9
M9KzPDCQg0GT9guTwj4+fb1JLdpNB17gzLOkFS2pHWbYwX6vYQSpj8JtnPPCqXWsnrcMQgMXzzdF
m/jvmi3e3MmXM8QC7Qt5uznHHWXIFWEnWXLIVAhpomau8hIIedbYtqYWf9lY3bs47gFZQa3avgFe
arKjuYuFUZLAwaGNzTiDdadUCkSH9H08S/SkdCVEZcMAaSnwQKPi6qc+UYcm91rrG7TBkk3t4AP9
wgx4ua0BaanKDYI4bDdumaL2ZmIlKnh1TPLtCrxWdfTt1VnYW/OIq6ubrgtaGelcE9UZN4PFCuY3
Irg6EcaFxFFISAg4937Vhb2Xfe573r3q8kNkQpYVB3bY/xEWKl72WMaRMM66Ywry7s5Alqk2NwTo
MzhwFsSQ9LnFxSHbfvOxSzC8yOK/lIJRKmn4F6Od+VWCvyUT8hCyhrGgED2OJPJgSe62qfQ1mE3J
okSov2vP1lw1o26kGaYDMiNByzvC0JRky4boubIrSvkSheLhM3g7k3IroOjhIsbLI7lZetT6HUbr
1oolrGBDnHJu8/a64uHdJOVnP+OpV86YQJLlz8Eb9arr0dzj7tRmWvN++3AxNGTfDJXu0+CJlKda
ovJNv/sX/bzLTeHQHjFb5ta5x4dkvFpwhF2WrPJ/Uif82Ik40J8WIAwdHPua0DNAzdrgmsowXHTq
bhDq672oj29OcV1UZuiRK3PwJTEkIUi3yrPeKiPoK4+rHWTm3kOppJnpz8dHH1FCSZnJLrU9KI4g
RQcS3w1wNQB4JN2sWY4t9H2qsItQbxMJ9ctwGurKxB0VeJH+Ui1G1BpkXgbZimU5FH6knDLaAAzE
NQgKsPXt7D7YGbEYJexuVUQtSdUIFe7N2d05ioSKH9EmRKlf4arWaQNk8FG+HWoIbyYupoFIC8nX
2HYMBCN/B7+PtOl5IsIbM4QpOk4VzaDuKFj/P8dloXXvQtzeW5R1xIUfRGOqXvU/Me3FZp5IydGm
Xg1lZswLEUQQzdt2QZ0ZLBbF3/e+ZeRdRV+rzFAWj8M6nPI5Vo919AhLQy+6HJbTH54gBSz1bSG+
hYTM/4seFxBGqTcbxmXFEgV/+dVPh0FQfY2ESnSN1uYFOpzCv17aYwicaMNUZox/v2LuF+1rHs0O
ngVZZ9WA6QMs6JClncW8QuP/g4U8lYj6IgKiAX80jnTeEpgyntAybD2bUc44+WAyjyfKGSfYMt57
rwsI9W+I97j1AfugeKLggGfxJI/c9DyPjdj86TWApBffhlIwtHc/Fiaa3jjNaGmr2q086wUv3M2l
cKV1IeKtMnYZtKcKRAFVsqVL0XkcNMaIS7+Zj1B6NGDYo785A8gT3/Xt8o8+T/KFvpJMWTJOgb55
+IryZSYPOavkdZt/b3dC0+aKGn8OxpCvk6UmFlRSdFouSi+Hnoqj1XzGECPoy/87o+/YyWzen1UE
hnddq4MnhzJcaxejVUsaKq+CTebUCaUAzb4WVXMKBqLe5yhYasbwvzGW846LO3u7xcZoKI82w2UG
c6enJtPIGDEB4UYLC7BvblQnCX/MdV0oc0+F7uUjhoqF7EIbxLQlC2buAbeU5wIMhTBoJD2P4CT2
yxtheI7ccV8ipg2n1DBlVPqFWRadWmSWSEgpoCwkXfLmE/INT68WWOmGT7ookqCEiHMtsw9faQqG
yoXTl0iGUkCrQoabXGfhtIX8W8na9c+YQnHlnfAKrK99qf88odaEzf+da/wxavU/jydjakrcrl3e
iYmji2f7rDujlK9B1fYmUfgQyrk0BuoS3AzKHzagqcaueQEiI+4CHRK7Hpau7OptOH/2BISQneC5
jZiBiIqwmHYXLdJB68ubBidsLIhBamMm1qPg0DaJEWf9SwoakjugeFTfi0WfsbSA1eqM8BKe23Dy
o1nyDTAVc03fSkw4IA21tAZWGGxLAkPWF5ybXIP7HSJKqaoSiyp5Z8n5bjXmlQSGl738X5TM9T55
L/S79d0RSUu1eokkzVchGLviOYqYYbKhZfs2aflYC6xPRilla8XAPLltrnuZX8FjGwmBi7jtiAqx
PY/T6W3VpoJurJYK8rGcCsLUOjf71DPQp6TB+HxrDpo26+4kPeQDicLhTE84NF/DCZePZVALhWZA
BxiQvMVRgWEiWZ4Vw3YHKYSLhV82SPTeGGGSbvgi8s7qbyVhDkjB3DwFjsVDnKvtxHFJcawagfLv
mZDatUld6gepQtXTtKfg7DRKUVzA+s5gqnLtog8AcUEGSpi2CEAtl4cj/vc3LGP+vjXHVVAekbfu
TGEBbHn7WJN7A01poIreqxyTPEWeAeFyONyF3w0pVp8Nh/Q2jxxZYBYa15FbLs1dTTCy0DdiGgyQ
8D9+zEJSY8cpTuDe+8j3S3CgR3XwwGozlly+Mi5QA6DvQm7MTqzR3xDQ5GsaZzO7hnmpNBsDydvy
aJ/7pXj75wIe5/s7EivIUu7UPRtDKtWC1SiltMoEu+oyuVEUbkCCCXGf5EAt+Q9Cqz/N+241KmqT
L4BNTS68CAvEbHMQOJO9adkVFZMyJoUCm9oAcSh+PQUsdDv7o9mUlAx8mB4AGPN/tlmX6F4bRf00
TOnZBwDgv3D1c79X7eZRWu4U5nJorffba9U91bnnXwQc6UjHv+epY/j5unQ3fDpQ3y4MBmStfdjL
C01BYJZSgCZAuHuxeqkS+rKBMImZXprbVnHhRM0KoQxIvxSUbFAKw0kcGdydS9yPgRZ5IcmI0FBf
GpLrfCau2OvfTpSwaBblWLmVN71aNPNWWzQN/9hZN0dQ4HNgNIUjgLjsftXax21k1zUh/0cbbVWF
WyfH2k5V/epueDsvprV2cY+uUvwT4ViJQWa6JVTYHBCSpRUR64ODrBdzC/pZOsx/T/4VXj57YtGb
jlLNYumxdgEZYLglk+uc7bg8q0gNxWY4StbRMq4KIYhaJc7CME3CSGeabaDNJBJKm9AEdiFT2F9x
gCsvTKA4QkhWIkIHYy3U6DDpXpmYVCxlbzp3z4LUrZZ6XUxasCwDjkqnDh/CBA8Lo5raFkatP2Sy
dUBDWHaQetNUMNtHINg4q/6X0hsUU2tunCaSi8YPIX1eRe7QOMgLkV19THelGYu9teS11lXK3ND5
4l303mE3dxZrdhfVN1XUnt4RaZSmDbOzxk0TXEsNzREMghudXyI9DSqwx9++idk0hA6fuuMcEyYx
MI62SSfokT4ZfpfyyYL1SpNFecycBmGlQ4JL97TwTcER1UCyoRYy2Tn/EWMWp/Ha87YbwT5+HQG5
joG6qGQv99x0egOj98SBFbPdhdXlHUfXNw9TOuSiy8PM28ux2+zSTb0xRG+DUp5Hy1F6H92TNSaC
02gay8daoe/4sjELgScb8fAyl0pafRj2DQVmBscZQSQqIntgnjxMwu0VtHSBSQWfSiFzC3MsU5bA
B99qQySJxjXtfJtR6pi4q1Is0znBYfdArH5cpYblDx18kqYPRpxT6VLN6qJZq6IMRusR7jclP/qa
bvmbvu6/4Sbh3iG+11IHHrCB0vf+CfCo0v+A8GEMtfSoE+cADljvR1uwap/UhwbzBurIdr7+q1ke
6s5o8PLKwmbpJXkM7OIbq71B7DxzTybqEcFnkWjBsvT1MK4JB8uQ543DouHD6wR9ryJwMZ4gHHTx
MN8g+5Uj5s2IJI4dV2t/73eIvfzgtDeYt0p5UjoSeC0DwcujNGaJpSPlVDcp6H0iDSg1dm8IENQD
M2JbSjQYQ3qxcZkdQ2mox3hLZEYS+zmJSD4WgcxvEzq228QWr0MoKTstX5eKYW6E10he5Tj8xb9K
g81TWopqzvWWGfKeZJGyU26Oyu9sft4RGHTEC0tVGXcCVHddusdQpNtQ+ApErnOBJZODZ/kVmDAY
vSi66jhjsoF333DO/DIO/4ry8f0RC5AZ+46JzKOroA9sOZkZZCWl7OR4mM9OrGxgG1G7rkycmZbR
hJxdWa8vI1zN71VvlL0Id0ajfn3lFjgcL51S0Yuc3dXQd7RbldmI51gXlUxEEBAQ5DRWO06+3J3v
X5gDlOOpLokA1tE+wCnD65wFtYsAGLWYSrF/NwP+oWTxPQLXvzN0+M5KIHMp03WcBuOs215DxCdV
3ZZ2cY8EK2gNCAA/UbYFG+hDmyINGEvH6KpANkT8gaAdydoIwQwxcFfB166UxdSSjKnwOEMHsIej
icjWNonPUkq8EFWiEWOoh6B7+d/WonQl56nG42pbq97VA552DPVyUKOTyjAkKYTDIjZH88VoUSY8
BasTkEThL7qXzz1SUE6IQQKC1OLQyp6yYM02EsqwYrV+s0r79V/1M5kKlsQIDrbb6TcGsLX9OXoa
0jRkaTGIEwOhtCi1gbf3+/wdUxwmEc7U/DZM5vpJ/NZRcPHqJeyECnlhKs+IBt91kSyVteQfkmbb
EQ1Mvs++lIsC5kSx+lM/i8WOhDFH8DxEv3J4Jy5L9TPvtY0IFE4FbPD6/KiGkKKGsx7h4ISEHWSd
Mmd3PDf7/cAMTpP9caC6UmhRRjxtJpxpAUXGq8k4v1f69RAvUUFZ9UJbfm05MTXvkFo90vActEvS
hoaSzsQWK9spn/e12vy1/BjPBSottearkjWcuK/RfpfIM0Q/SSe9RPwT3w0NJJsbZVWA/DZz+vmv
LBrqJrZ58FwlsOnaElgoBPYTlzyY1i2to020om0KgjOsR7aAqRoGODI+UspPD0iPOvuOrJpvB48c
qymRH2EMa1fP6NH+gJPF4u2oMO8iYvxglYY9nnyKXas5rDrfzQE4Y/GNDkjurk8Il3ACfatiE4lr
9l8cwW3rukHgrgW+E20XAsddj61XLgP0xsTHkBIS7UejxtCeLUiLp3xJlIoE9+HtZSPZOZrCZM/+
50f3Reaze5QDgbsFsJVe3Qhs/lQ1bgjSjdMin39cCJzdhzBI17Z4OVPOoqWQAfVP5qXGFVCZl+BP
EWYxZBIz7O+6XiFXLZw9Q5hJ6NnaFaR78q2peP4hHgn4p2l/BSH30Qk6ZJyuFwzNHnizgrm8/Rx3
bhpj1z4IDn7rVtPdMfaGtTovNKh8qgtLShOr1KCru+XA1MZ3/6Igeq7+w85LZSyyLeC9gvqqswvk
MgenXOvjTB9dhxhS6TxXSHTnnMaBEfqk5YoozC9VnHRoyyiL5QX6vqs+J1Cc1I+BZHTN9j8VckkX
DXz6j2WCqozQ4haYsnlnRhblGrNT/HPBbADbCAjVSPVGuxQHoelJRxr95WuCM/3g8Jstf80h4dRj
2FrqErFGm45/W1gAG4VM0O/iMxfPkesPYwm+fbCfhVrAB5BqT7ACqpGoJyUhsJEQ3hXfiixieL64
jcqYveqAuNb9nFOFf8uXDlicE1CffLAqgMXXQQd9Lqo/G8jbj8y0ZPQNKbAF2PZt9lDnteFf8Qse
3UsAfb3YR05WmzN9qESj/1YYebiYdUAM/y1RXSpYsAFx95IFTQc40cUduvgI9BjLF3DGrmkwB/Ta
CEdZeITM+Jzi7wgIF8+g9HVawKrluuNMxzbt+enzkOkveFc/V2x9f+BD7Js8gcLiDeNpx9foDC7h
49seQHpVwwQLtq5McUSuDUk+Hr8FOL8yLwG9MijljZ1/pQF/cyxb4M2NBjVMAgnDI6/g5U4mfBB6
aoTz3pJsi6SclWMIssP4Sq/aLkJP+uiWIjKpx1eLUSzTcDrVMp8PWq8GQddQnjovkG+qGp0+kYuA
rxyWJSxkuE83dzHxqF0ov0aUwrFvpTA/ME3lDx6sNVXIayNnITh5+ZRnSZx/EVzmhH7N1F1djVxK
rnNGtLHH9bA8qgLOA0I06XHNwZiOj69dWyDgNsCRCme9ELh/iFtmxecEB+/SiMkfGrlssWp5Ggjx
vDxKMY0lkTxu089KH3uFybpmAMnJfe1eZjetfLq6JJvtFYcTHKRsJLoixzR9m+1Bn8NBBtAfwZOn
T5foT3fR3HU+ctoZYO5eZqQPspgAodnDHD90IwuK1vRSRwOuyDUJFwKbfdOfRQc+MDKr5jiNemd5
yY6epDOO8cJzaANguXOODS4zpCAWgGO6XE3i0RIVjT2rrL06KsA6YvcsNMj6doXsXWgXSxzp8XgL
XFSOEExi7+KBfKN8Htk4q/HSvULZS9ubFaGhFLTiWil7wOWuzOcTie+znzZ6iFv6Xjq9AiIUd/W2
sInTyYZLL9J4sCMfViHA5MQ6jtZAk+ip5hZsmw0hWg8dNLWP/VI/46Kp/Ka5lqz6dJy0ueTDH1q3
z6Jcvj6Fich1SApuJGpCMg5QNvJUx3AheBpzpkJdEYcjzTP/wZQRVWYuu2WK6fnQnLB4LPnjJzgA
PtjHiNCEzerKb3SjOCJOZt/VoBXZLeNpkRJZfQ6uY3s+LMA58/+XkRv5GDd0vYm91W+REjj0HAYA
Wr7oMcJ8gqGkHQpkH4z0iX9AXtFbndNJwVspFWLw6+Ssnrn7GtWgobs9AY2WZuhTuyBMz2hRMHiU
8UdzAQ6GMj9yH3gdyLxvzIcrXhQUm6tVTHXyxOwVOTxdpHDwPVVnHasVBDexPG3qiS4uyTKF+X6u
UCN32wXXMe8oPo8K5af5hTxCitgGdqIEjwTijtJGwQqlo4CxSHSCe2gza2D7xURJYYtWrUsWgah7
VRsy7qKqUcE+AdnKA+giIj54gTsNRlX+GoDY1hrj4lIo0LcwK4kDgo5LB2SB8dnAnhj9yYhC7vtF
0NcLmdfYvya6AlDsZ7mqvzYYndusuCxgsNihJ+wMWh3eDAb4XT4yELGxqnbUL7NhSyFQGk9N9Gcg
uZ3bkspNxFUknfi9d6vyozs/ABnO4Z5PrB8TggTpMVcw8/7FNO7rmUXxmWPHZtH0XEi/YXR4e8QU
iIi24UhyxEkOf4OrSYRXAlaXCTyienh3HidQDNMCLeWERkgPT0kJzF/mNg0kcSZuRlaaJKt5x/21
vYTLmRMEJy9g8qJG7oLthx/aoO0zOZlvp0KIGcUeSb1Y2Ph0jtjKNCeY/PJ/0KWdYDmd4lemM2uy
Q0njLJZgJQNKkfZRJOFX7/PS0MJQNj+d2Kn8wKtDFKCDwcp5Ki4lzLha+jKfmDg5hr+2jbvXxN8B
XWbNRkJz8UwdAgjDRcFOLJ5I5hQSGN5uYCeHaiX+VWyabXFi7SkpkDyQobmz6b21j95suWS/odVE
sqqjzsMy4+kvu5Ej5lLATEIzObg6vfgAV3lJ5seittjt/dsI1zcDpklj7F5XVa6d88HNCU7gTzUs
GvNZQqcOR9MM8zV+8oNPV2+kKEaNmEE/WC4/mwO7qbB034JlFBixKq++7R9fqcySfak8aZSskRUE
wvaP0cJfkEyy6tCMBhKwqUazgx6AsEDhL0ZNNnFj7fovBfyhNobMvp63nUKS/EieKfAbePkfvZG+
TJ/lr8Z/CS10ogf2LPyJLlLpE2SyeC6btVfLY5P5Bv18HqoChsBlCHEtmeZaqcqeF8LcDyqP3A7o
K9wpVnlltJfQgRj5KhRJ19nLxnA6YQzk86YqwwuFWAYKl1cIdsZ6TSNMQ8InPqkEgGCGxNKbO3of
dUvzc7bElbacDGuoOEOxB1ODcZfdJiY0rKGc5VdKgXD7MPTCnqO0otqanCwPxqc4iGQb+Ti5OK+y
kQOhsEQrhNRgmC8Y8X8hzzxfwjlpaexv2zNNDR7aHF/eSr1wHEXEUy+Hz56wRCl9cf+dox19u4oZ
aVDZjgnNP8QvtFPqeOFOLv5tBO3ITtClLm9uO+QA0zvfz5Dp7lhI60HqDZFeFX0NqG0rVxT96gRL
FCabOXQrnsy6g7jHM9cPlDr8vK+pi8Zt+zGCp3Cwfud1vcHDqb2afoCgHbX1oMCrtEIM8/HthinD
/GWP7MrtbkZ2e0HJAB0QCoSKl7fkS+zDJOaROKOwep7OgUKZdU/jVYqJp8EgAGVe41U2qcdRzu8h
qcmFQloPQqRdMTvOoEYuWZ08AeYqOnTBh7gqzNBveitl8xlm84tm2whnFCCemOmCGnqvgotrj3z0
lo/eLDqlS+kDvAuM3/O7BfHSnZeq45aKWkmPu/RKJDiZMWATi+jnMuNznRew0uJL+TgckZ4NEJbi
gNkj0yqjMedUO2sYUEROhIxSuLzWh0EgMsN6Gy2hNom3+UYKnDLeF8U07XIKusiqGxGkUIkZLcIS
lrpFJMbmGMX+v7IjxG2c22K3bwTdnV4sdPUapsJ9KLbhDxAgcteH0IYNftG3v4nNd+df7eXyQcXJ
B8XEgBnFGQ0MuMDNfuYjTZZ0lb/HkTrMciQiNKUNptf6bCMHwgi2IU5gPtNyskjLN0/bSyf9fCDV
j52gMKYr4NkUsDLnVXozG8A5lJ+fnrfAulHuMaey7reXIS9VLxkd64891NW6Qp9ls8siBicxlQKd
6cEVo+GsovYttU584hWskNienhHxdZ2+JfHenkv4fvLMFMsIn9n+h9ItJZNmVKiMoJafN/uclrKL
ZUqMnU/gbB0Kfwy6CMtL86YUqM9jh2OsRKu5CLN2jy4XOTAuUhQaCogXlpUbTTUpc5qpeK0ew85H
s9azQ9tPmjlim1c5lPmLajySFfvuYNw28ClJawbbJ/p3qYpcWrrRjjnEppsVfPWNbaELuWKYJG2u
+2Msn0w0vgvdqhkTaxZc+H7peuLCD+M+/Iv63e4DjIZZuvzvKRjhx9j8HBhoZ8o3bZra10pL7sn1
uLmA51/LiHhBePKZuHE4S3KYhXLjmJVTPflF52jCslloyBK5WEIr7YK+ycSkwse4dCN16cG3DBnY
2/YzYjlqDqW9E3JUEv+M9FpavlMFavfTt0xhP+mgJgVCAfBezA+nofycOod2i8PcxH6LyRzOMvkM
6xTQZ/6369UWaSBJ/lfhThP4nP5qjdqa8I15Ocjhr2RkpJwAhnEsb0pKqKRDsngtGswqeKsqEhD9
2m8bbQQX/jWWbCiNL3WO26H1llw0vAZNq7BOwV8UZThqSXuORSHc01A2HB1cjzq5RjU8zXPUiGOp
ZOYpVY9cY0j3EZkE2y9WZnyX0EOLb0icOkaIJ07pBcfEpLIKeddjDVjQV8RNgDnMfiLu6L9OG+sY
uqM1ab1yv4p1w2oYXM68RykJImavF7T5FinfkcrccSrWtK8AZXueXbNoiemMgJgSpl1rjlGsBi0C
3auJ8vncisNoTHvVXUWNE7rEHJKaaeUTAm0ZFVcQBc2C+IgEnNLDOyEiXvcFUqOGX//uZUpG2Ek3
j2kfd20NEBPEfui/x2b0iuSOsNJQ1gweJTvqI8suHO/cxyiH1//TSkXTfemqhwmQ9U4LHbxEs5NF
c4rMpXr3wWOzbPriuSLyCRJcyzkZyrK8A0nUgUYmYL1FuEVlmjbSKa33LSwDD+zsqu8iZZOrj8dR
PzDC0uU+KcjKGB6SfcO4R6CZ7+OFH1obIbXl5dpVjpR/e1+JBhnokVpJuQ/NREGbvyTBbGmkhJVb
sEveHdemHVZXyXdGEI60EuiCcd3UFzs/1DuJ87GkYQ4pN8xGj5gemXKsnhtDFfb8dSx+v0G1YmBh
sAYQFI/5mcIL6G0E3AIdYqRe84FE+UnHlNXhdTnuH0hpgWM5WdTbiarZvF8jzVdbGJd1mirpYOq+
qVYArqQK6/LnSvXOJc+dsKDSRQrzB4xed2/oSck5rxd80tizoHOrbmK2Uc60C6uN5CMoRbT0gLoF
MaB112Mdrdg4mYVV9BZ6ZAu9lBiiaSC6FTMXWGCSNowZNEgnrNM23KAdISqwjAnAiWGvG0bEwlYZ
MDXVkqcVK1/Wtjkw0mSO22o0PDoFf7RqV5LEppHWftfoaV1tVVoPH6nJVOW4KjyWn/lWAqBaRcPL
jqtF/qjI+OlqGsWFOH5/ccr2AVpCvGjyD5TBLK5twWxSeBZlPMz1q+lJ+YG/lwx82WCAa0Le5ZR/
18PryjUZVlXBb4XrkmBYHfdCy+2EbQ4Awv/RQ77/Cj/N2PsrDeVuAk/sJvurhbRDcgFe9AB78JRh
/v2/xmpp8QnaiNjpXUT7YewBePfJIxpufPgV4rZeUDo3zzuxSauv00PoHrveTp4Nm/+Pfe3Q94tu
Vt81kzb9K/Mj094nW6Idv3z2PtHzwcu0zc9O62EJzcOi35JIxqCnculavWj3JmCuaw6JYCjnlEvy
tOIT2+rrtjNVw9AoDtlJzZrw+oAF06moJfLGcrbSXErV0bTzbspb7c8SdcVQqJu3t0XbsInFO4cC
R46Sg1d1YkMKrfvMGbhnrFy5A2zovlPMqQR0JKG+sIkOMI9VJlFJZo/dC5s3OO8Lilfv3eox8A+0
rO4OlairXJUdOcZy62jXmrX7t+HaSYbJb9EeXvLr3Nk8O2n0USmD9vGM+IIkoVqygcr0uA/otGuV
Re2frVlS42WOc6nqj4Y9f98RJkZtZlhhPfc36jFIutD+tf766jNpO3Gp6fr3SpJzJQUyRGIk5tW9
NIczG+eIMOScq97V0Jo4yLE6dbLqhacdbkFD/p/GeDIw8r9ZJAD5tHUt6IV7C/tic3/r/Z9W/FIB
ZVF9ftWq3uyGsKPD6o98biFqAAb06fRElHmmjG47t5GLsOVyKLX4pb9w2BN0Xd/rqgfY54B3EIIw
ZYEpVY+w2SNdigZ0Xj++Kv2Kt8QRdUmGkx39nFQshP7nWH2+TKdbv8bpaBel1cIrnUfJD+Jc6XQa
DjED5nPMzzexAGpiaWNYb+BIHqqjh34Axp623/tnlWNCjIKS+pg6+NK1Mvz6ewcdqs/yiXg39KeX
w44y7FYxxekEc+tQSASQidPWFLDM5/oAI9Zs6MwHLnF+dQM6v4rzyDG+4Z03sVoBJrrk4D1EdLKX
6pRZkM85ndEAZsBS58pXwsmHwXAGe1pynjAyeiAMhsjWde38C7eS/1yQ1lp7VVB00RwAC8As7PqR
3nX1UZ58iKt1rOpH+NqlqmwMfMBR8MudOu+g9/fkA75gwiDACsJnDeF6ZJMDXkqqMJt+PEJvzcSJ
TTjYwzyQunxr4Z8puFjP7Svy73kW/SlI44uVrp22t10wAroHyqr1V5t2ZhobuCIb0FdtHtFq2CC+
WEH2jMxndee8WBOPZm3exbO2bUoTwMIdoxF0KrWUYJNyyVAd8LqC+ddQpPQM8Fv9p8ba13MV1dZB
fW5x2I7jwopOV70z92R08BVKTca6AXX4ciNUU/Urg3nkJj48mImMIMSqs6BJBdXrnMhIEXCtQ8GN
DorHeWBROUVTLxpLf9B5rR6LKE53yDPcNph9ZZxVpok/N+x82y9rKWkE4O07oZAJT5wtiSTp+nWQ
Ath8hRfQ+JrILoTvWLxyIeUDA9Ptd7uisiMO1HK//x5lN/4td9TdREWf9W47/aUvAD2Q8Ll8SqXC
kW6EiwlYFT9vsZOClk5BSSXg36c9jU4V9L4wQil1IQId5/FAdACktgTtMdtm6fu/hSNY0LvwmShV
vc27osywoHuuGiLvnfZD6yI8lxlURJXJ323ivVIplcqQP9n7qtx/AlJsZMlzQk1KUtLXbLNdHixm
QwNQS7gE/zLMBm0pj19hIXsQOowb08RLMM2ruveQ+02LP95rPH2LGqzjJ9m6tIMdBhoHQzrOYNpU
RqVnwGx+BThv5UxbVBsV2fdkTz+V1n/fXhmTlX20embHZ7KiiCiauT+gdHifBerg6msYWVoCtI8m
oOWqIzdNaF40W6jXgJLtaI0zaxu4ROVKWJVfq+SS3Zl6W26PPqML2egKwoUMehj75kj3E7xpC6co
+KY/u9SxKEqhltNB8pnZzIT1yDE1QRNBA0P8tPa6DfTm6Pxkz9EuCt/8u6ssvEpBmplpDf1xmNkp
qpf+YDjLy1AzlIshCTReLZ/azyLwYPoxK4HD2QOqEq3UoIRiEtmHF4YFvjZl6xf8sb1glYlQKcLJ
SuYlgmblYal5BA6HsJN5ODvmS8znovxgI+cnTbdlXJQnfnESUtz38xJN4GuzDpClLS2LLbdpCTVB
BXusBqz21GTfg9q3pbOyj1Xg643D4MF9m5m/yd7xDm2uSm3ZAGO6R5O27vo8FyTkHgV6r+aZxU4g
bCQJRy/nFIGMl98fCQ5744AKoJCijV8MCduem0bJFnmGOnFpv428GBq8A/AOCHLU3oHUtehrDUdL
d1k9i7jNCJEajEi8Chp4z1cmfvfCofPqP8maH1mKx6irraF7Q+hh32p83lYb1jcfH4R6Oc6LMtVF
KudPWObFKRtpYv4QD6qi6qzu+LMeiwoxBFCc/Bxg4gUkvo8lvT4beID2tLBFZeZMJB4mCrGXrXUZ
uxRFZ8pYDK43/D+whaXJlsDEypu1NL9v0igIcZpFCggEhIxEU2nAPbalUJpUZVzB1mRnHWKejUNK
foxlkGLi3dfXEzSZnu4kTp4jGUj/BHQixY0NcPK/UYP8+KiwB6b+Vb22kTafUgUR3ElVR0LlDsL+
OuDC0kPFlMdblwZz/ilWQ9liQumplFTCXO2Ng88dB3SLyMn4pantKC83kWiXEc/pLLe6lzyLLVlI
XUnE2AO4egW09eVoFIOb+DE0HYqwapK0QCzV5A1+M/LJ3VzmFKWs1XkInRXJcby47jr+UxE3viOT
lBAWR2WxWgRUKHYxdlgswfElznMizvSmheh45FaHVKk34i32493Kzc27vJoK8gwmcH6mKzwXiTrr
mBBTyOYPVzEmD8af4hXCsZayE62F6ihtplL4UxWiwdJtaVgkqwx2JKDF1VUS/OxEt8MYsDVmG92H
nXm+WTdPn3UNfdmGqCd841LHtSvOvFapLkiGJkhQeNQngaUor19VOZGXJJc195A6xUq+l/PjIJpv
d0n5huRu2THW/AsbnrfoNno9Fua1TnoRXet64ZeeKXbXalLh/fLHfvusqI2UPVGo4CqRVXoAQ3n3
1mUiv2XnVTeefE0v1OHz+OBOWeDWTPN0W6v7NoiyC8j2BwY32C7RJi3sRadxSuIQfBzWXY0k2zkZ
k1xvbFWUAcLpdFHi5YSMf6vVhhXNZBAyqfxGjekfYZiOaVWudM2CChgq8ut/6JTZF25DxsNANjN0
R/HBE8mn2bg6TJMdt8l6LQehtDpysYiGw3TlrM0liQ/8CMifFS0b/Z/YJtazO51jhv80AW1vby8A
ntUt+ALHmWtxeW/huxTc+5shb6EAY8l5YlT+f3xjiLZdjKJTpHc7RfRq84pSxU0GapHS298ihoms
gM/rdeIXauQeB+dn0g2WY7qpVamvTfC3GCf8kTMIbupaa60HaC8gFi/uKXRa7d2Gx5YwvJBHn8Hj
mMy98J1h0OxPtlzfoFUd2mHBC3ort9tQQ42fxwzI//yZjPr6AJKwXzl/WdGipIG1tqkgS/LB8T67
WYylj5PIwNyr7LaH5+RiYPqIYalXQPDKp4Ry5JPg9Bvz0l0yI321y7016Y+YwUbKdTQJYssh0P2k
nTSQFgX+2Fdb+adTWLbwYdrAkFmIPaGINQydpEYBtP25Qvy6tnAmFnpVNaslG+nKqKYbk8c0s1p5
EICqoem4QrbIeMin4c4tHmr4g7HY9pNFNkXfJ4e3zr71aXwcfFGdfMDx7Fy3Y8j/dP5qzcnUCULX
WR+BAf1CGVhylUo4ECSppVsiEh0N7o/j9Hi9gvCyF3Z6Ylpw4jgR+JJZIXdWpQXIcrWA//Cxgpae
Da+M1IHqq0W5s7/Hu+X5VCZ6Q6kqnCr0AEQqGRkdWYHkwNxurG7mILkQYCIbk63PVZkOR58rfCgV
MgfkqU3QhZKOL8rXwG/SJdGxMz6Vuhk2MpLW/aHxxOROImtjNwN5eBUkxYIEUaBWVOMaQYkqUuG7
UCeFYKog/MuJIevFULFNKO5YRXAMvKV6lzi8m21P/419UmcHJbtMxGCKLm7C+xOB/Ml/VX8U0/wP
mKdhhHg483OjvgrYvZLqCHCyEoEiF86ZBBRjsZb5LeNkh+FLqSr6uQViHySdOhJS115VFKVaQ4NR
sgpD1Ad0XrXjCkckGZzugOk5YuJPvZVK8Wpu5adyCJtFb8MWzBpHmb8iC9B9O/5HjKgSzjg1wETo
Y7gNr1EYalfSLaK9g+mbQGtxim39VpPiQgejXR52gVN/s3hU1REPJUCPcPE9wSA5yhZzSgo2AvAR
/elF30z8FX2l0lqZrrRyR/8uEe4ykDeCbBex0hQ+ovd3RX90FP2Ec/k87zW3Qp5TdcU9ieKMS5K8
li1UP1GIHjnAIrzBFF3CMv1CvrhbkLCFaA8zEM1aBcsph18TfzGNioFKd4Q7NLLk1ftCFn6Gdlsr
zXREJQb1Bgwo8sUuRa8ER8MEAGGH99+SB4YeM59Ck/2yfStgeQqWUWOX/2gs1kkOmd8VD1sGcWsn
iGyPR7pQGvu+2FLFqHZmVCY1kLvlsCEgeeFCpDd5BHEmfmkfNfHHmW0IVXQtOpmuvkx53fJ/mqJM
F3k0tx6SKQQ5Ttijlc8RiL/jfa7b0Hsgph5+T8n+WUtaIkBlOqlxh0ZtX9R+RycC2/tHUmeZe9+6
BAXp52qC3mK5wW1qK1FbB337G3ILASvEzvaD9dw8eGYW6whZFN+QyE/21+YOupeH7AOrzqcVILrE
/HzA/s82pQ/R4hw8dqmAnWygb12W7LE1h2GpQ9NyN3ldNY9DQVHP4Wt+KSTOsDJy9odwnWyNAqXk
wilDTRRdhtkB4hdZOWiLdP7abVfEAgoYDEAitdkSHceJB+wNaGG961HfxrjPMqlOXkKpk2LeFsT+
kI5hT1AyN7W2gp92PZ55OJLSs/hoyrAuEeqIPViLFFJH01UYkxyFb9LRQv2AB3dnl9h4ceO7+fAy
ZMsKptCwDRInmn12hLFsnWrOveipnw1GD+/mugnJEXQxikL+9DQanQGTE1AGdklu8WPUDEaq0mwc
5nxNEC2KnMctTvn3qDIALUpDipvjv25LvqbuZr5Tn8HawLPDdxvvEtsPmAPiXqe86UVWuq94cxGf
nmOcDXzj6z4Ue0zXgVfxnvSoqkBt18BV48Ck226BVJ+DRro610u83nZpzm5gZzr/BKTary8p/1fV
nGaStao0qQ0PTANtQ8Wbdn6HXopeb3W87UghMGyU+QlqgJ5o70SPuS3JEB1n1uycEWTkLzO2OX4D
hWUQUATLVL/gw2Npvn2HrtDpRkG5VvX1kPf6PCHtCmsgYDURN60B5+3gs3Mgn2bXWXkgrGb40UQW
KtwZqu+nTn4Y1QLdIZhUzghqLpwepXIMnvBe4Ur4A4EXp7as2dZldRYD+3eGlW2RJrW8hzx501uT
H2018EzF++WcVkQAQGGvIAJ4+rBDnEb4jUX/r1yc4CLgENf2uq8DNRmirH+RlOp12L1x1Fb4h1Nk
U/g6kQ231MmJlAZMCrruwOdJ8Wc+BqWPBMbaEOTsDIBt5DuFWUQ6AwLOREUwO1ZPF+hTfSTeBDrx
X+JzZdNXZMLsk4PLtlB7Lb2AvaadwqMDldFIU7mWJPgFTwlGlEQFj860oMjfAMCDqY9Q+4Hr0pwf
wJGQoT28yf2p82b4p01qya4qpLWmi3rwyNX3+A/G1aTG6gLRtzLsPxBrSg6DuJQj3HBThfWJb+0W
NcLMnfyKPdu1KdDs+RTGPdGr2xVi7F7Ih4qXbW6dSZ7vDLTSnUidJmuaUGlAGeE7AELdjYS8hqRY
v8sKw0pmAjfXTmnBHYnnZYpFOui/+0E2lqTr8DgSFMl4l6rmEprIQn1fXztPw8EW2rvQX13/gi25
kzEEYNvwPbRJgAiIgfVEvX5D0GCjXGCZhxRl3x62PIs8rUG33beh+ns17NNq/Gd4UXDQ6PVgO3Ln
+GysdtT4oJBFoPZqoAYTlbZF4+N7tO79k4S3DpTOroCREDp7x1b+nhzD3IuWa2zVUVNUrxkslJIE
BnVR7/QQXM3hoG0tbQIyt4i3DQ6RhRa2Job+KqL3MMyc67UK/gTKRm7mGtZegSTYH/iEGVt7eZxU
McCh3wYirh+ZmV5a4NGR2UqMDwyjVQjf9c/Sn5tgy+bfiXpzF4j4dbAJ3X0y8FK8odR39Yxa31Cd
YnsebqgAyGv/pp+KgzD/ZC+wcyc2pYg52gbSRLORqJEswpjNihla58r05iPtbl/6N8E2uObO6SS9
1rDf7O0iAMxORVn3V0B5yz5OxdtbqM/3gtl97VtSP8q0mmnWiFqFGJodIEW06IEp/Lf0ZCnPI71f
oNcV/LJczDAu02Dp8u0Puh9umZcwdoPXu3dPLeICr+UDC64NbT547QnHBrEJKrwTaz0t+Znrzvwx
WfR6oGvqnsJfgj+hYUvdHMvRsCsOie4s5YN5UxWYeZ5ptdCOhwGpxBrLsjPA20bJHiZm6nr8tl/O
HetkIlhCwprzfvgXG8ooAqiCORNGURv/mbFa8wGx2ep7L0UmYdkvc3+ENks5VRpg+IJ+updqUbto
wRekkxWJcXR5Uy4XmjxO0Y8mncT96hf/F+B1y2kJTAcCrKJO+Knq+HIJnuZwoGu9BDp+OSjtMvxe
/c7W+9yXTEKsBn3bvdFSC7Q8Y2iBjpJIzeJSROX2Y2c8lcEBZc+NKDsCebbznQQXhfa4OHAxwzFA
YMFcmiHQoY14Xw7AN1jiqgyD+qff/9sSDBpt/eNVulJqTO5DPBO4aWH5NUz1JDX3VjKLbuxQPydO
KoW4uFZLSHTUVL0OOHIgJeXXJPy6BG86GpG8dNjb6XyB0j8maRuCtdVPkzyO8ckc5nZMZb/Zmk9k
AQanGAPhUH22XMuSq1a+QhA8/85+awvO4fMNithT0j3lr5krao7/Yv1BotzaOXhM9FM1fqhNCX5U
dRGPW1PNNqBebmihcI3zqG9XFhfQOizT7MsI2ciGX8nog9uFO4JC8WDfpdYXFk8km6wAChLlUr+P
PyqjV2BlEHuaasOoAG4mgmKxi1l8sAVglFiXxI97Nn0T1IfBX4PHdV1UIC+Nj1RT99EHqLQJyU6f
+na0/mO5wQLs0VPqhbqgzsp8GTaRb76g7rWD9248Hg89mt+Jj6aD0uKN/2B8ZzUkbM37wDDTh+cH
qww3MoFKBVYm0vuMQL6xySvod3qpwF4GfkzE3axnuKx0DfL9t3oHsvtvOeFg3idiZTWgdjX6mJ61
gSpcghCIrSLvBmiQ/+x8AoSsc+4X6lh1Ay8NOMT4rb3WoX/c98PwfGhVNvBXFGxssqifLmvr1qPP
IOdSvCcfUhsN1M/2ceZIQ/2RG3V/BRdmUeBzwaNu8HVSZ1KSKjhshc1r4RkrEZVMWKEyWple+YO/
u/NEIwY4f4SFCxd0uOsBStg1AGQCuI6gHTv0aU2uYa5RpKEDpO3TX37rXRxBCSbbnInOhuqn7Qo5
ncY4ZAEuPqk7cdPFENcLAQA2Rt5wHusBUY8Halp72O5j1yqcvwtoU/8839JAae/WAKHO/EXjOD8Y
BEbcTPRH2rP7FsXUkPfCOgoULkXqfmTXjL4ufW4wWPBqKAMaEhSh20Ixf88UxGi4xOmI+q14X8NV
+J5HmBZ3k341svu2zTWapLwhzIzU6G2t8TVVP78JuC4H2jXo4slfkVJ3+MzbgTMaRw5mLkpdrZAF
Ns8TESBqoCAs4veMOEo4MZLsTLbdF/FVZytaRKk1eZNNDZArdgw6csi4q7k9xp6Ce7ccMERcYxQx
oND/8q54owjsW5XSdUvpvLMbfGJ03P4TexQqjt41R/KCwNOeeMHZRmLrR4FjLo4oriJtankPTIHv
ExWS4wS6H5NbzQpp7lkI++D9qv++xEc7OfQvH3RJBDqd7REdgelZflbHu1NCIiZpUT9AMPkFodnO
XTJiTrTWBFkc4VPaDSQ+09NlVVJSQiwEfqXzbVKiia8UezAJm3lZsr+QfbzM7ROO5jfwIv6g1lp8
Tgp/jgLHW+cjz4qwZyFexFBjRPSYhI3PkFngHYdjtPQC+79ssK3RgaMuTS+EsJauvGpsSMCNsKr2
+mdfy/VeJIlC9kIiaPGCB5EPftvpXQJpHyFlJLgJwGhgH86NVRayamWGh1zdCxt7ZLD8minCXNSE
mir5pXM/uOFgOLkEbTlprnTqlxfvqH3/q3XvGGXqvEHDJFWQTldSt+r3wYDJ1caaIlaSiWu+Z0aC
3Xc9BgrBApaJ4s7LNEdLEUC3b55Q2YEZBAlz7n1kCQwM83dwQHfX8HGa+OuoEMGkT8GDq8O1rbVQ
0oZ0uPnihb7HpMIYZ5StsGy7ptd2PGRx4QkimTPm5DahzVvoUBpt3vDmK403a5zlJjhOOHRi8wOZ
r2V+o/M9SR+mi9gQ795cILlcvMoD9XRPLYklHnW4oA4R7+D4FrmKQKH7cqqHaWDj0BmLs0nqFZnf
IJBb3br5eA3ZAlCKIc+9/WujFVMTwF83tMUB2agsDM85l3IVyV5KVJKoGw9HjKi+jnOMUkkKsZJj
3hONK7DcgU2BpKeT2rGv3KTZN7+Dwcej3f9STmIUACyIr4G1hSQtP094K3fKyBPQd2SY9t0eAbTO
1xegLty3QYLs9yMco8AHj9YnJfxKOY1USMRuc38Z18+dY6LGSNrfXYdexICNz/TguEBBlsS+PIQN
0AlP6dKDPfdjIyPpBSVdQKPhB/8kz7N36Bn1aqBdk1s7QflRXM2aUQHXbwGxeZev/N4yz13L0sNv
NaHUEWbzJ+99o4BpPPA893qdpff/MOqotx5SaXY+AB5PbD8CxMhP4ft//WlmOJScmbDuk/VSubUO
wkPQbRr/pVybT4lLUQdo2RA7t03JbjyVyxJfEvqhSA0D+odnPzMNTNRzomASJMhNIxT0izeFDNNz
f6F3XZRjIbwio6gSpSG8/pTPGIJHC1HF83fSi5Zo3KLnTZtNQwS2oJMirA9x+eiCT5kRFgTZB449
5cYa63E/y6uR8kfyt3iaKSRTBAayIZ0ohj//RIoJ1ErppuwD5OBv0pIxfHK/6X0Ij5r4lo8mZ9f8
r1nE9AlE6m2tXkryCgcp2l6aWNdM2g2yfPAa7rU+zze00vBPzJpmDbLJh/R+2jTBX6bKVh5JlNE6
oGmGUd+KKXd1wFACKUqLMYSdMnRJ/dMqAz++Sqn1mDR/88JumND7Qd1+LLyhIJY9Sn2VuucC4yDJ
2qHvtb7OLqmyUXQLxG3gd/VSUxHqn4mnZUD1DQX0NDQuVwLy8XyVkMg30SVDe+J0EGj5NcR3bqqY
M3EyvUziiNLniVae3YcFJDyhjI7j+De/cZjPxZdg/G5idh+3ip5xzUL/dYZyAz9iTPl+tueyy4R/
ZixpUkNmkxGPxFbfpJsSmz/F/wotDRuYM6k5a9OwKpFD9aqlvb23XXvqCJ0x0KSbN4seXXYRwM9r
VRsbCw5J30jxSJ+nPzOSxqECK+EBdJ6Xc5zFpg4oKKqG3OB/26VZm1tQxcC+ogQQAqsqzUaUdwes
Nt836RqHoysmOYjmC4XB8jRMxZ1kCYJHhqV7g8CN3hyYZoi7b/5uztwdDJpMACQnFAUetra+w1na
ADa6ynlH0CyraHSj/crp0ZjyNGMxw7PVumWcKAHrQyEJ7HdXuOKgz7Jh4Tr7d51KTnezEzoYHM/4
JNb6f8CBRldV0mEvSpTcH+/DoMfvEluAVLKCv3zE9n69AITTEZZrvk6YtL1d375Ut8DwnBBH41dA
dsCfL1YGP3nlyWGhWhPMY9o4Zrxdw4f/B3a7B1cci3RVOrajBPe4JncsNdBr07mkOEjGYWyEL2PE
0D7icZJrgSXo+6kPRtFW2txO+vjOOA9lp3x3igVPwbpJitzEtcmSm4Rww9yChNaDuIHivsuHqFu5
2FJMOYpQUUbTlUNRaqlllBe/EnS3NdzjAgPGbrzbZdF1xJ1IR34gBGvO1vdyEr7ICjzzI8Li1153
0n8sTnWX0eWDzJexs1JvjVtUzV0Cmqte3RdFTrvZOTMubhK2ZucnOcZ0Kp3gPNwgjV1kw8QhFo8z
FVL1vnzQFaO8HmuXMU6NeoCSUFBpdPOtIXnIVo420YVzfoOawKuWungOPnVXeQG6aK+vyuaF1SGt
kjRSchHRDCzR3oDW6ecme3FefY1+MlIpMYM5wvahNP0iccQGgaM08uH5f+WfDyxz5k9LU5AMj+9v
4SEjWctblxZsusPJwj5reJwdBWk5k4eVtLwVs4T46P2LbvocCc+7qY9XguaZjkilAjaR34OkptDY
+16uQ2XyfrDWj9AnXhVrtt//aofxJuSpdEFURwZ+MU4AOXQjU2kaUFo2O3cWMspsVZ17Hx9w5il2
4IgaaUppd+o4si/D0god6DzufF7UB744TCZ0EvVLc3Xx3ajLNUqqzbBigpKnzwY+bDzFADpLaNmN
R0jlWlenBIbG3EZa4eCShesPMG29liZnx1a6YIKbjXdbHLjMMXnBir88BdaUpBGYm4v917GVmIRp
ebGi1enTZCcc8LXd2fNrz+UbKKPVFtZ5DlS3Tf2zprCMbfq/G4YFCVAJEcsOdsksa/FbAAUBhyjt
Tlq5g/XVAdFYgp4HJnzqsZNjA7XkroOuTNz9mgTgOgbTnGEawIPitMWajJ0fbpCdRuJeJgbMN2aT
F/M3KGM/M9b4HvJ6RCVYCd7HW94a8juAO7AqQZ87Fi5KdzbrfJn4V070v/sWwt2JMl+5RajecrWA
99a+qVN2vnUsAnC7U/pELP3yHAwuRa71eSdeWLJL2rTCt++rCwmkpjpW9WLYtFHo7kgCZKWDkcOU
4vmaG6mnUxz2SqW9AWqAkGfnbhbuuyUYwhjSH+dmd+3sI3P5vLfuQrJCiu3mU1gfTHke/Cyqz3o4
osv+3MXsLv8xT8gMBSZ1es9rspjT4mu9T0D74MJBr2yZQUXjBufi4TG7VeK7WkAZyHPI8Dvs+U8G
p8bPh0kxCj20/vNnswlIMknNY2UQhI5X25hTqB+z+1Wx6UyDQ3VZQj2JRAfgf5N3ystxxtscYtA+
019aMl9hgeJqAFUXutOh2iOL0n6RwZg4VhmD3nZfefdpUaLruBPRyLruk6LffLCCa6J4qU2Nshgf
loa2+ktfCBvJ1XYnqsefbIu1U0AQGtePzNBjQAzyhHHXnWqj+4h2XgB+vLlTVUyL1rGdv1/j1Jjn
BkMpEkqsjFlY/8Xq+pMX9z4IuJG1d6s+wtL/8fX+Na4vE47rZxT0n3yVXy8E4AzYoyXTchM8p/Sn
W1zIVGlxWAImc7zaijvq89xTGmg0KnLBe0FUKmVVwnjZFxTOVti3DMtjNSRYpgZ3PNZNMbwHIlMK
ZPDlWCRVl+F5ZhS9+R27frQA84cr/D3b4xwihz3Lvdv25Lm2Q5fHXXoumo9NyHwIcjRdjWAoL7ze
k3MRWE4ApGv6pxkdFn+esoF3vFA4O9nmNxmc82Bil+EPw48YXBI75O5whgs269R1c/1V4BjqiGph
i9cFnaJcvry/cIMLVfYp79XyQ2YyFVdXqVp4XFM67W5nQP467aBMH5T/poUCHSJ33xFZmIO96BMX
WWGDiX8k7oEyUeuN6VkdFHBc0lqVt7WQI5CAMfPd6BvlFci5kJJqzpJRhzmMpf/KJel8qtaMJ3ge
FUHGA2Qp22UDvtVkKBJ8mj4gR72LOOVLk2tCUFX71NYrBtUZqq0FMflJZ5m+USw1/o+9Zs6c1mzw
qicbrQsFuIcfEkYPvaG8KL8STkUvMf9J7cwH6rMa0LloFl4NLW2PjqtA9ZWfzhnzYioQArRaTuk/
EwoiINgQqj7L9AV8SHPIifq7t3HZS9wDw9cZ6xj8KTwClMgtSuJ35/K/KML3HN9mjOLl/LbCX46l
eYvZMkd16KXR9kATO2Pj0/P0HyBEDwvgsx26pyoq9y968D+xzYE6KjsO7PXZW3RYYXppVBKJzZWe
AmXM7Ocm8hy7/Eajlt4epFz16I/eLH9SY24q4LzBpc+2Wnco2V8wgJZWEirmdMsVzFJDy8KLPMur
AV15ex38AvKYYlmdmAZZW/PQvqPj9BVB0s22sz6XqyJx4wXiec3eo1urSBC/rf29MzpV/0xFsYmS
fX/Myp+oe5Yfe+YKx8k80QnF1EUhkPDt8FktZc/W8i7vFELFln62e6PC05Qg85IZ9CVKDUyEbyLK
w2JvngNZ1JwGrPAGBcm+a/0l0gqzsESfilMEUmpIRzKbwot0FEatu+kFI/hBCwHfO3bdHs7gEPYl
n80tCVV1wkKuCwj62nka2R0W9oE31VBzq2PhlPIkQKMdCv1TDBLeFz3vEKqlEUB74oP4MR7zHilp
HIuvJogfnctYfHFSxEr9PoG6JvZ019fO3s62+j/4prmCq55anwFIjkFWe2R4eB0HGhh5PaO/e6AY
njvdemJL8VqF/HT78HfnknrqAYws36zx5w0XqodzHDnWzPCBLcpdavVu/pyRbUoMUTFWkeEHscvv
4ark4Lxe1e1zaIVlTR/+ae9kGVAZ/nbVl5BKWeCzj5SuWWpdiktF4wzzGpjyAJO4KXfWIzT3UwLf
cIrF4Get+lVjC8p79nIyAgtAbcMottAgTnN8oL+DgsSXcLWFtP3PkNaXCafBpsLCQqFaKihXUm6d
fnJanjaPIXv8zWTxLPkqEHgnyDzE4SRHV92vodl9tRmm7LjYyq9Ex8uoF0juWEGTqAcnOvBMeHnb
ZPIJmrQnGXUv50Zkcy8jdOP5LYPzEdzyVwJNEDBn7P4+5iUzWJPXcFsCiCAiL9geT5ix71EFVT9Q
7FhLLE/h5tW7yFiWaDxDXinzQhBYIs3RUgBXiWM8vHBA8rSG+vzNq4mtULefi5C6NnHso+FZtl48
zCRF9JYw5cI7BPzmZGIkPKe3RKplgq+5pjasI2ez+COuBlZYXa7NZKvNhsjL3E0yiBRS7ivNTNLp
PNOSbZM5e+ovgtK1y7qZW2sMTxoboDyGq7LuoHloSSLvYYF2au/jCDKAu6EWeQ6rO5mY0/LEddxY
f8tpKJ7ChqaJX0ITXvn4xZT955JqvmSgSFi7Hn8Gt9gCbY+VHCbRNVOKtu4b32CTLjmj9LIej4lJ
e1GcLdpN5ZpvCLmTkg0TPkNwkuVoQrMrUlejPBiCafgEDuOUO2OYAxgWVl9ZNJpL+3FDa/SJF9kS
toytw8l50qw0AyW274f/mVi2dqfTUABuqCHJK4fD8o70kJXp8SSnGJ5YISMwP0hE9KOgizeJDAjJ
lIw4RSP8emYRPxsNpbXNcMh4dTAzMq3X3ZoWl+tAlKvZQ1A8PHeTM5UZy0D/WcLDkxLVruVIcotH
Vnvdsyf1OJjq90cEdtVqtdJuX6H9lPQwEHXy6goXObIqFU+q8yXaWc4muNo+cZHk2A7gBQW5mJXj
fUHFrRLliWn7CQB4i32DOn0sVq8+IPIDnkHKpXgRAGLHwsObm61kKZVLFNCbkDriYvoIUdzfyhVt
u9Ort3CMZuoc+2U4jeGpIa0WbfjNcmDCMwgM0lx8NHmrN9SQjEUGnIVHQyb6lpC2uZlzjkCsgujo
Tynp8uCRXsvOdCo3umUMedyluhbqafW1TriRRTPbfs2edMuNFK7nSLe6y3+rgeNJOOewJJxzoVtr
bn5BVRoU9YW/RN6gpQXbDE6t7Ek7oaPaBzJHt1kwUYqdTcsYzDOihnz1t/oPv+4dR/0tSTwRNy3L
7M19Oy1Yb8ca0NDBCsRxszGz1ymdmhvMQ71sWBj4rArDbeDkfZwjFMzulLNibMKVlpOvweWO46tB
Kvz2ePr9vw4YLcIQ5IehGqw5tfjYWdUW++AuT51vaQtY9MBRIlWH+NYEeqghPkMUcQRdS3jFmG/t
2+Aw3RrcUw8slGZKgOTJyZoZvCDzlj341ibBzCr3qip3j5fI9cmizHszJDW5bH+PExM6t032zzpa
l/FUWMeE6M0awzHrRADSUwsJ9ojDHu4Ek6QHXafiX0qVgzkUzGKCapubv+MI+apepW56Ypc4dSB6
+75QllZi5A5JnBoeV08qn5vLWwadidSYPJDfi8wzY0XbRBtPipm/3eUE4HnpnMDslMEeMPq7q1tR
IqAmOhley4+yWCdncV0Q7FjhUUsb5nTX0IwuPvqNGIXc1KbAQTMVQ6spGS3wZuZ35S63dEoh1KKN
0GQxpHhweoceZwKjdxn0utCg0eQxgBlIMuGC5UwOfd78rycfe6egeFAC+TgSkTZpu+pozh2S4ODd
sCossEOHFcnjR+4eTdm/h4tdiScYpup8dRAu3TCElZc+u/8fDY+2aBQ/vZT4Wm2/BR8evnV3OhNq
x6memPdWbKcLIFzxaRNgogIQrlhfk5c1+2KaakZH3LsujIlbX/m70t8QOzGcNutqfGzjuknrusex
ZqVWRUYuQAh6EIY2s8H84HgvigetwctvML9OeoJ2+HSA1Tc6SLPxZzgffPcETCdkKuFUDhNEZc3D
V0IvxnPZozQiFSX6kbLB28gD2EVWjE8YPJrfxWOpiCP8CM/rs350/KlQHBJKqIxDGYuXJ0pRgInV
XytWuNQ3lEnbZ7gcZXbHSShf6yq1LSa73aRGVBrY02JJ9IOD9faGvE1WlwNz5dbuF1BzZ8KnoKJL
Ycb3G+OFleQMQBp+new91ELS9xXSRIiWl8BNzfxseGZgwWPWWarBc43SDXK+jyfdy5dFhgCJ8viI
NVyqARvRl4gy9UQaOeehc28CRP3t6N4hLWajZr9Zp3lTeChO5mcghvG0BOGN9VWO9uxFDn1lJdvL
PyHFs0W6KgmpXUb1sPbUwj7iGJ+0LjmqhbtXdjjldPyw0n3vJnLFcvUqGq2DbvsKpk+MFbG5h5PP
ijDStgT3NHdHiptBs2H5tiB4eNSoqKbo7kx54y1KVQYUH4ArThmIAQ0iBvzt0uBmaLMfgPAcRw7B
yQlIwjJpd3jlAU3cla2Yedgs/Cs72etdmylYyusoIdRgnTr/Tstva9ikDSsvJ2Ey/EI+SGSDCRK1
FvDTXrg8Tizm1xXN/1TtzAS8Xj8zs2qrDIGiHkfwCOXPmVcSXBvjQphVk5gocuSNVYKnv6b5DGVS
de2x6hz2ONm6xUdNJyiTXcAb6H0Ok5cFQYw0YpaNsnf9nvJpBWPI4fQuIds7Wx8OkjiF128uFOF7
Yjgq7Hs0tzK9yF8EoqS9ym1MhF9ou02T6Tmw4F2kpqN+JwC2zPr6D66v6ruysLIn+Q0HIC6lPNxQ
nyG/QphRmdhdO443/v11ENEsFgO0+ASjpTZRIi8SGX0duouzvcrW3rwb+FBtMkXTIzC+YUVlaCQP
pz/IIixzU+LOMd7UGa/j231UfjvMG0Oh8vj/pRPJbewlviQCJwYDQKzn4wWbjzEjQ7En0eN5mdKc
pXGzvma4/Xsh5VsckuvF+xQQzRGSbAV8rYXkXy+UX3NB4KePYuV4RjO2R/6vhJ+pOBEE8IpJYUNn
nrdsZ4JMA3uBtWMAEQifJ3toKkHEeSYukqJM+jZsIdcEYYlla37YMfHYngn7Ui7uBKxz6TBqSy1c
0kX+Q9y2HLsrdM+rE23uqnqNAGNPLJ7QZLn+MLWBJyiOxurySa4MbFsIagJytBoy8p+u2ip3YUar
yu1AmZsSAWhCaFyYVbdPuWCWr1IUVkok12ZYC0805Fr2bRU3skY2OMOt8fIXVCIWS2LX3N2gViTu
C91MJDKCO5eKyBcPVmfSvHrnhQMQXkeV5u/yJY2yn94Rc+JU/t1Hus0eIkMdgtm2tLEaBbJDelBg
e/laC9XFRtbJwej/brfOMRx0cqVcPTWDgIy/oJ8J4QSQxH4ldTR48niZxqjVTJM1aSNi6p4lT2U4
2Yf+4AP08qEZ/dbQMTKIZ3ZzRrODz2Wgy80K6M3E18M6n+tW6MbpYHWBaY1RPl6VkpmDlj9tHjc7
PP/IxAO1rbMrYGUFhGKM+YDlBtxeC9rJG9OlHDBpIhrhsCmCpP3b1clRTES9PncN45WZ3fnEhJ9J
rP6J3oV6tc9xo6499EgGE2W7e4V8euGNGrqo4dfqlgCUVH5k/DFg1pvEHAxM2A1o8/j9/zzNwtOX
Fmk1UFOknzI9sCJrpM67CZGy/ZMdQTwP2Qic3acNJBkS+2MH71DORSzquYPEi/WTFWMiL0ecE5p0
n1VgephZh2hkIt6C9292gHlhhtP4dKK1kFoF2S2eIQeCCRNIq5BCS/b7Himhwxvx6xmAVcj7STXX
bG0TKuPTmnvulyJCTxKQKbG9tTdJsmJOwAcXqS76zdzLEg0Ej/aTz2mrUV9LSq6LhB2Ww/SrfJhv
vCoNCHdPnI15HIPubLKV5GEQymYK1PYWg7YLObNAYUevQfvpVm1npHXyRV5WQx3sCXHF1wFers0/
hO3YFOIqbC6QY1NGQf8Bi4/9hHtQisjE2p7mhIC+6GONuPHepeiU4gijxD/7tkwJ5zs/oijo3g9L
QrNgjem1bmkQ2ARIH8LShvzcKcWQSzMOVUWzN/5651MdeW6YG7W9r/VaakO/kNTsd1/Wb4iAcRWE
dqBzzVcBYfl9rW4PFsWuN83dO19/sMC2svoA6UhfKk/I9mAY9hUTgQYV0sh78z33gdselZ2TX9IZ
qR14pSWdBCvZE4dXjNiwjkbbidI32tJfaeCnF3HNjoBpNhjWcnzWJ6I3bhh9fUrvG3s/4JvzLUta
AfMKDbWKaB5xJxdyG8OlNKJb1jGgBhfHLdgsukySZFOpdNB4sVebL1K0sgAi5SSAysX34QdKFbwV
IR8rmdqqStYT6nJZ7p7ep8wcwZmtEZmaX+PPuKYcUnBgonw/2tOE38QCZRnbjL5OHe7rCqdpC4aW
M0OhlIwhp/PAk+L8nYdvkazRnm6p8eNSfrzpJb3nfmbusmPLrvh5MaBTup491fNr3E+Z5cjERm3T
0UlPlx0CgtfVzPNR+wVRShxu6Fa5lw1PVkGyj/+Z7dyIPl8BWZPbFXDCjxTgsl0usvzzBUjrMiP0
EMv5D/FzyGBpJn9oKsi0T/A1yBZvn00ahvdnpqRlaKvCEhpW0SQV/ZM+aXM08glRxHuhflPco4LF
094TL/qScymn3Ur2XLw2B84VgQ5QSZ5Tw3/TXiF7gX9uS0JB6WJGXS2H8sJyngY5PRygbNEI6gF7
KKy8W6uCiIwq6t8WLS11xkbLfkSPCIonqP5u5cz1CeWFb3cRwwwxGPtvoJ7hzdwnvvDVOAOyKsja
0WJsmPPQs0R7AFLCWIYbJgQkH9QDUVDFmxIqDUeLbFd88Q9iBsMN1srDp//QYqwamJPuEUnmuBdl
8ZAYR/Edag7N+iFZqkEDH/7SoFHqcnbjh1mP48hivmapaWKZopzSAhpoDqA1SCdzVwJtiB6KT+9s
yHP2gizdlvNZ3Wzld1N9BBAWZSz2RTNyOAPLtGXIezacyPLylWe0IYvbfATFBdCN7XycBAJJp/sc
QjsiN1MgC971S0ESCYN69xoi5X+4awk6Bo0rIU7nOI3X4d/amXmhza3h3higDoJeJCTJ7vjhZogg
rT3pGMe1siXKw9bDYYimUDUwDgd1L0IEj+aYqGLInByuoAioTVXQUQSJeXtwc4q73F2W4rIbXQVr
fzCU8hM5teVYtkHkWrjJ4VJvodBZYuQjrtOf6GpLJZ985HcjXrbuFhZoAb1wW1UV2sICik9emJVq
iH9+HHm0ZPw2yEEyJFA9jqFTSPu6ZKKVWAOZjlVOUFAax45rIGycjr8/ctDww0zh0L16CAx1SNWn
KQARr8OtsoZGFZltUclpDwj3psJED02NV46v/0LmsurM11d4OMeI2kb/0sM8Wk1e8ZkbhXOs1ChY
M4wOhSWGUXtPxwLQ2UhKJCHX/1nvGxOMtPi21eg7a2prKBH0KT+EZvL/Sa3NGrG2ZrP1j0KNvX7M
NbaqS8vDswpAwU+EXWXx2RhLXT+4kfwCnf964bJWAX21AM1rCkQXU3yNWaSBxzb0zKZnBETc81L7
hIwUm6Kn3Wnd7kX/Y2tptVuejBFfoI1mJMEL0wnQnkeWN7K8vyNDAgSCQi/pEkJfCGnlDFTl7N8q
Cg6nXvhx4ZMr4oQ9ahmDviRQTWYcQSSF+huAr20C4WrIrHEPTgrOZJx59lSwre3o05ML22Ym5K81
a06lJa1Lvoar6zMBq2fs3EVnRxJMRz6TdWdZS+QzOqQYvFbPjRdCswc2vdQWmXxIU0CWSKrZeV8E
qNSbsg0MEIFmKTfz38RXfZTaLEK9iJSfROXGnqdPegm7Wkf8t4LjThn0SC9g8500UvDE/NwcuwSQ
+m+9pz+ZQIQgKKfIWlUrIZskSqJ351gnMmtvboJr6ZFFPtqinZA8p34anoLoEFFqMY1LRI393cVi
i0lamLPEp1bI0vhauY5L3AJjBPPdsF0D21lUq0fY4PFJVt1wSDPsF1pjz3+7IHuKl44GOLKhS6NB
1RXs556s2a4CbhX2fY4e6F/DKzkDpqSms+nSuW5ix36nq7s7PFNMPP7RqTrakjKTyg1Yklcu5p5G
aVv72+CISENZqnox7YMlHjUqKqqk4jZXU0feOKzgxPTHqubDQi4k3h32zkObpLKMqqE3lLrryKLl
kEt6/k4t9blpKmml0b1h4vO2maFbnQx0xtvJriK3BArgT7m3QH9KBNoq77HMRGZpYIl0nhT+ZPGl
doDBY6Htx24PDfe+56suOyu0cwFUVoP3LU0oRNQatj1OJlEuDFk0vfmi1DqE/dt+Zzqp8IV1Yy5T
ASP727LTuO6YI4aKQB9PJGMls/RZVRMsJaY4rAkSH7sj7xW9L2BdbAMjCNfeJ712WzVeLCQfKzu2
o08ErTwKVoobKDwVm2ug+JCc4+CK7vgvoN2HfPaypxP/YiZy78zA6sOnUNmMRKkQj2P6L8Yyw2Z2
XnzZW3GNbeWVOoFZsTZt06rj78f+oDmtBzFGF64TM38MghgRoCAvTdBgdTQklNTf9Ixbh98tv/nA
zYJa5Me6om8yf5O9PKl15LVBnRgBvuS/ygxuSv5n57RONyv8xnr9K8ILqhq4L9lbjVL+WIQCaFmH
x+lPrl7ufZbzDmo9UgSp4Pc001Yn3rHv0IdiEk3fUxLVhxIn1EvU+o22A65yGNmnTaZwSEH1uCI0
WG85tYltzr/gVxoMW7o64VAx5GTGiNn2ansI+y3vr8yEmZjFRd1gncLy08+1HCQFlEePjeu+9RAu
2ANgnnNzVg8ZL76zGHrHLlPzohiAyHx1DkclN3/YKSgnhTUv36QW2dLK8Rld0BEpSVTVuAZkkYlQ
NzsWe14I/QXFf61+5vdZPHNlqq3hPH7sexQg+rHY/UGsLIHWBGOPJMQMa3HLaN4UWUG9UZ0GADiW
yG0iSsQn1dlkzF9GbUuS5/EtK157JfNKG70BMeyNKhxqFJsaRPLitJEzy505LITbjp6KY8fODR/D
a/7GZ7OdafsTpn9xuYA1liMFl6f17cGYeI9L3FSNNTrJtdVp06fFZQs0q6ClGS3THWVJeJ7o5Iu9
m3uURF/as9QOcd6Tpv3TOdAykjMEjnqM9Gic5G7fVxVZ4dDjYxfCQFxTxu4Rl625V0OSBPmNLwYN
uaAWCben9u7WOgSvgd7kPiAJCcLMWWmjvHLaHqY5K+NquSDjxJ74dNxXvNpNjxjFmsWIv+m2zyG5
l2A1Tq8bLVZNoW0dv0L2XSBAXGGXU8s+ydKLiKjWN4cNf+hMfWOcNMaGlcEIcILSCVmBe4HboT6f
/unM+XmA7O81gxOoWLNDkURWRjSN6WNdcLwsg2iNQV+BkoKA+Hjfcn/DBeHTD7O0wFWIteDsR5Qt
+k2eC6O8O8VgAi7F0m+NryrC2zfI7S5IixR177UTtxNojy7Ho/HcJ/VtlTcrevfu2431hOdOGith
kIh4huhPKiCUO/7pF+qnUZzsH/9yMRSL+XexZ+yl0lmdV4MpkGet840Nx0PadYqjnDi6CjSJeDiC
3GOdMKiKAa13TnfJWXV/RhJfdg9LwgRBN3FtRlkRfft7xgMrn4/WVPJYMxDzh8FwGCT3GE+o7IFC
dzhMtcZ0/+k0Pv/xACYPXuRgf1J6qYusUXAcLIwUJFM55KOMSYsi1vI5+tgT+1U4N9VQRL1tQueX
ZpY22jlQ8TanhHYblcACKsoxWZSrW5RuEaoDAV2rjqpx/lH9PYLYWRdyVx/LJlH43vH0RBvEIn7B
P4Pgr6Wabke+qw+ira2qnN6MoER0zTHCLTgCqJo1HzY7N9HKJDQ7qyWy/FbIGThHqhZKfON2/548
Mbaoys4KOfHhof43q0a7mD8jmDDwh2S9+o9Ial8HXsqO5geApIzf2iFmq0oWmi8vFLYsznrTMF/U
JzncjqNEkzoBwzZgwSQnblgIJpTudwUP472k1UtP/SJUsSus8Zx/tBWQBGd19kh76SCCJB+DnS4D
HZl9uPVqO18S8SZAzPZCrqhZxbb2eNQDvcx2RnLv4IFY+aMI/9DfLCtVdRjaE5PIiNV2myWb1ZXs
lLRNx+LyuVpRm9D4gqkuu5okeW85gXnrEc7B4iyTnF6quyAHEzX1p2JNVUt++KLQjbOsVvnu1oXj
mmhj8URxS1jR7HabNAD9aSIZ9xO6CuE/fFgDIclzg3Wsa1JmQLgGTFCf0gppCBSxQsh/pb5SMBTz
mfhH7Biobby41Rblpyo94jHf5B6RUxCIzakECoEc0VLd3j4ToOS0ywW7Rjla8+OMkHCibysjpnW8
1EhmoCBhqYY4KFXvxcr5zU8s6S9UvrqK8gwzkgHQC3sB2wcpcu9fPWVlFFRLOQqreW8O4nf7ud5D
LekleKRUeFT4fUvG4v2YpyCZXMWIcmdqZ+wFqkQ9hcsz8TD6hYZPjXDehkgcyJH6Vk61QsxFJ4aN
hUUTmatj381CYwSsmyGwJYDQP56fTK48L5eyWzt8pohRmPB6krXvEj5nYk3myHS2gmdHMfssScuX
LPyf6sim+Wu2aQFBvhbwyQHOxpLsrplNrRmvYIl16Ps6n/KFGrNIvVVNhnRxArsJ7nqlRgJZO+xx
GIsY8XLFCtUXezwzJ2Jw762QoISpK0ovok7id8Jc4OVPOt9i25OznsufdXW1km/26xeEyuxdCQi9
baOy0lG5KkcDstJmZJWbo6F5wOBvWF/xlL0D9f2r6qaJvTmOJCSCFhEhWSAROuZbLDmZAWqMF8TL
DLJOuHcF+iZdglpOlV3kjm0TgA+KR++XOS13LWOnJnvCfh7OZkiT+5klcVgjUjRJ9IzVeYTgNGEh
XIqSCdkv7tYIlwB+gUMQDRfhILq3P2UOt/bBTMybCoSIeX+fTOUAEr95LAEOacSlZ44ZEy6RD3cR
jo/DfIBGfviNigaV5Nw8ErB7xfnBK1rq+x374U6/6zS5Lv85fOLIbk3pAIzihtXygVsMpBd3MvgE
5XD62wQqSc4cdxv8AcRKskNwjf+Im01g8iGwakxbVOzSDMFrIdaQMBq5DxCpf2OiLPNpFKYoMxPN
Zq+4kcxYyVMPTEaUkyzlid6tv5KRNP/sKCXvyLiFpevX6/8Osk4UPIuwGbjZPI06VjtfX9X43zcS
4ODCyPzJPRTAGME6OjP9qKd2eP0vudeNfTAHmJZNXOiRGRY4CvpRBgwBv/ETUOkczQNFFCkF0Hil
UiNBQfr9xHuqUhgc9uWNNEyE6dOBZc78qf6PvzI3Oh0vXUG48/kObU5gYmqxhFYOSwSe7pv8mc7L
/s/qLClLM3+ayj84j49jNRSDCS2QCzvcqqIHq7g95bFgeZFTeSJc9wFhUC29q/mYJ078yjl7DgTK
bpNZ7BVR09wDhCKqKFh6GvVlWQraiNHTMMHMpCyaVmuNt+Sx68X+oeHufNIbHFHl5bhTsub4o0b9
oBYWTceo6Sv62DPXT8/AC7CqYroZchwmUwGaSk3s0lznYoe62QN7+Svp03md6Dk9qRGYpb86HnbC
nhywOXjarojZ0C4TuRxVfOMwNo/EiU3ES1G7LldVqFJXSpQA63U4Lewo+AB517x626py0993zpdv
wRxVbbWmfq9031QaB2jy0ekjhL46VWguJY7ZkrZ46metDKomNByk5CkstOo7yN1niFK4kgUj1h2u
E/EMqjKe8Uk/SI6jwXYtjw/BNN86yEAThSKY5P/oBk79lZzTVkMs0ryqGtKvoG6HEYMg/Mb7C5xh
+hqOYe9mfkRu6FGXgZ3BFHS2BrXwiRiHH9UOOleSWB3/pJPKnlhFzDhMHtQSpWudaAyyekNbV7mi
9VHd9FtTSi8ahowGEi0ZCHfJjIPoZDkSizgOb4rpUStrUBSkx8GyJP7AOrxWZX6VgEx4lSLRnRta
nBt0a4Ua0WSLY4YZUKCrC1s83YClJ4l6cODomvu6SiODNtAn5Tmivjz2h/zyWsxo3jUbzjQ5pRfY
9MSXE+c+x0sgSUFw4tGqW3ElL9mF7O1vZmfwDGK3jzdXrkgqYdtRIK6V7eixAkP6eeg3DBNjvNJJ
wOLRrDn67BIEGP+mNtarkHbq2C1GQOaMCGV6F7p8EJIMWuBnsAbegaGwXtKwm2l+PUWBIgW9yRH7
wR2TgdZ+h6Cl91GziO+YmIFw+4M+tUycsJo9acgY5ctOtH7/DPMeOpn3WQiSpxjLtK3guUFkuRXV
nkubJXOsaI+kZnyllnfFcAHK4ELhyA04jmymDQNJaqSes2oRNtIJB4hoAhmvs/oTJcCUDkEPHmsR
ucBUIphApaPR6j/FwvEAtVeq5tNu8k3//Fi78nv/AckvRljGUa0uTjfCpddl/ABNIHBXW41R0CGY
+hWiB2LDIhB0IF49FHQTh+p0bes4coC1L+Usp3yH3llNuS6Jx3OtiA01kOC6ksbSVEL8v0s3AiiX
Jeii6wjhZxCRfo92wB99CSvF3bUSJ3mPjhWRjeG4+s/yX1Kqsjfs3ZVbNQ9gqPiXX1I07TWnt6zR
Th3xbqPtaBBsbQD9tJHem6LyJUertNhBIDxloYugpf5mUIeR6n4FVWXCCPjmilYb0/Q7cmRiz2wm
8F0+1RCxkpAD1PtWIEAc1s2YZ5io2nEQYte1XDp3MwsE0sy9iuwoQdctodENvUAGFL5kh16My3Gt
tnrQCCZaZYPwu/QXSRxxN6u/8FlSmvBKPiTjiDnm3PPAw1bLDop1KrN/tM/2pJkvZkEf1MbTLtOz
aC58RA7JWUqmeea5wLV30sJKgy2eoxj68HdirvEoaNUbkLByHj/+EHRbu1eY817cUq3ctVznQsMD
KkqqgKdNesCIKjOPnvoeBcBCaOr8VcrRcoY8Hrcdh9m2B4MSc1flp+qh0Q62ZH36ZxeAtYKdZcAt
t06ns7/XlqK9I3gaNbzVIGK/0bUcVqmKNxwZIcygUSIVYbH/zRd+evkPzKzmZYjVZCLNhEypjXq2
WQ9KRbZj2obiKgfdUaxZSLb1xj6piVDOlZzqJ8KVj4P8kLSV1ktC3rEvaaIG2PlpNXOOcqYCtQXt
21ROjtYYTNlSWl5e6u/AJB1I2i+gpoqu6cTpkGpCZRI2XJiXisYUITD8AvaWQ5MlVjTBxWR5UczU
Chaqh39ew4ax/IvKfN8Eh/qSuUbQPGiqHlzGxWkGv2lHUQsLmqaiyOOPE1r37XfquQMMElW0QnL8
hp3dEo1gCEfVmy/7zoshzUHSZE+WWseR9L5FpLfSd7Ns83cnt+KtxjX/nY5dW6ZL1Mge5dATI+pQ
jxp+n1YdRkoiGg39ddoHXPf/83EMq/NLkmOykIjMYBexo+CqxE3GzDwFR7+LgaRljV+GrZrof2N4
j67eQsURy9LueHeMWCFb/9dSv/5qJ5wh6B6Xsdm5wKUhOPhbEeEZft2scQqknnmQwQQ7GvNvZvnu
BRn2rXqhpEF7bOp3EIq0CUV7Q61vCXhpONA6G41tDe69sPCvhseioBebvskW9EtSNmkOh4NgphVN
jdlk5upWwLd+laE4peZjuapEkKtFrqIWL/MQxq98i2oIP7qth+DMwSA2XAmo5ZLhYj32jt5WoA2F
7DozJdgNXF3svdhGSBLv+ay3Hw5FBt/ELZBQcYiyUGiGW7HQvmw9+ai7DhoaLGn7sGuNPgGnuK9e
IDkkOzCdyi3JgGBnQQLTDU0fUSu8xyfyutDoTRU19kmbQ2ZavjfmwRWrCcqNZxl3jBBphhYS093Z
Sl6XbnFpRbYTpakC54B3Ce7pJ1AxAi/KZ7dmT/F7uhwTTvd2WxDATVelXZ8QEgCIwx3M2XZp6zr6
QCdZ5G62wbx4tvzmMGRYuvEzMLrwyoM9HpcCTrungTcgyaQt2D2z+9QVfGYRwQKpp2mRlATNIwap
4ylyUfyTxA30B0bY0ldHN+v6V5raOu+tIk0+LrsxoxhlPVFrqlqhkjMxknhG30u5dAqX2bX/Hjew
xnUrhaMtFXJDbDKoYz7ONUjtZOaiguagyGoGiWRIkOrFd6oHtyAGo65c44d1bXEpdjetVU0dRqW5
bbWYX2aYbuO8UL1T7q1HtEqpTyZAtp5cQ4hnOw49MicXLUW81td2ahCGhsF376Iq3Dj8ivV53WD5
o2BvvmrHV2yHsUPYjb0SxVrvBBVexTOI4O1o/3dUE6BsRwM5qvVxrQpUs/R2aRaC3er0glDQJ5Ff
pzUDRMBSzEvU9sFqRU3LurVrrPA7Tl55+XHfEUGcUYvT+8yxKMxTGPQo1G2vkYl5K1wM+25wZJl8
3i7CwhIcnQnQfK+ClApJsoO9kh1MLnHDdo5ADPN+ThzjE2pw8+MjH7eR3dXQ4a7eugjDnoeMkJVC
mfiYeLZdlcOawuXktxLzCId4EoOLDLQrEYm4vt7jvZPAdoBQPs4JpKmZglen8EGwhQhJ5Zpafhaz
dVkVZ9HQMgeJirXuxrysD73WYOyLYbNMFRv2Mq4ZRAkTIZsQjr36Bs3PQwvmT5z+L0Xh8QpOtaX4
xW4H0MgzRTsLVvHi4OcSLLnXuxudYag2Gf2ftIq80XuDrx+7tcc50DST6nZsijclvpAJsY8Rr37C
TbPi3j5kms5vI6N9J3cR8ee+q8tBgp8RKb6Dy0ErXodtwZPboVoqh0etf0MCOAEzSoLkATQCJYLc
xpe2beKI1r8fn/tydT3qxoooAAC0eGvk/LgcWWuG8LMfsXl07n6FYdGnBWcXe29hK7jVIjp8lOKZ
J6azv23FWgergAmsuoryYhNyr/4BU7GzBGZfEopMAihqKl2/FLsxqGbk2rb/53rfDdNPB7wsHf2p
pw0oJhuqBbqVP2Scml1UqBqkIlGZB4cn15lgdWG7FNYq1HZ8XtM2yG3QJKvMjdibmCx7k3TCIsBg
1n1TmpLJ8vcOBL/xUhPyvXM41ie2TjNaVfDG9l1YIrFP0Jb4XmWF4btbqtOG2YNu8rTeTDBqdYKb
EiDUAKAAnW2h+DsiC2TyVkCECgYuposd+46nRsJAIkEHWBF3e04gShAoHA8oB01bzQy5N7cjRUgm
E1BMUhmxKwsnmB3Ri15as8d0TM3z8LtCPlqzB34JiVg0D4dTrxLR7SY/kdYyxb12OHHBraRaPKqH
05f6D7MvXbgYtRYXiDn0yXyT0wVQnEtfWwOlGx4x1lm2Rz9l7nKjdD5cdjFC1MmhABZSJc18atJ6
vkTbfJoQseFEQMX/JkFS/R/7kHjHitwVaUaVbf5bZGAJF1sgXljzYEPabPttIkFBm+fqJesiT0Om
FzRwcfXKzxab9hSw+9YzK45Vf8F1iQiLCbGxS2Ta2PHXnigKUZpKr3mOlZfG5o9ai9npOh+Gz/Ni
XPP5fDVYFZgACpBb9WmHdFlUyU+HZLd7B7hNwU+3RZavR07Hpt2xkgjx9NlIEparWv+KXqYIjasp
Gnwu8dJkXdqYqKfgiojNg8iblK3h5ETE67frqsO85GtOyNnm/yNuRgt6fqcBVKvJBYlfTggTBHlr
STSvtSoFhRXbk4EaTWgNXzCyl0DhOXSN6juDvWJ+MELP+f4CsuzdODwbkBo1K8HkVChE/oyWJJSW
O0a/2ONxQ1bMC/CFTYLLmZJBzYPjhPuLvNiGBaIHxmQUrOvTdFNKGtKGtGtjAR3FiKLrPgzqp2N9
6JfsL7LdnWrCn7SkW7SOFDyPW1rCzm0kFlxPNbSGb5dbcfgbzqom7/0oFNRHkSg1ZSXTyEYq8Wop
+cKV7KgBeMnWTChAQ/XAU3tCJkra9683Iv9Hth56oy6wx1eniWVXfOmWBnGM5N3RklLTt4Lc8t8l
9CArAu/9Ly3aEeRvyKhpZirEcUG3MiVb2uUemJn1BIm8GDUb4Ov1QdSR0i+4odx3bKyAvVhxsg85
WqincjTCpWCeEKtU5LgOJmBmcAzkPPmtUo3MXVn9SOJLmT40FxUhVbCJcAMabnEm8P/HCDDcheWR
gZy4sYwKny+P33oFVjBNqTFod5cOJsyhl0Nv9WnmjfUM6VFHHpu5r/9MLDIFdzrpGY4YX9E+7RL2
1c+8dhM3/XnP9s5MW9kQ4B5KEVnqbpgvCttoxx/3RsT42PhfaIdIQu/QpoenK1CM5UmfaXKphvwa
5NSDlRwjaJ9cjTeZ6N3CUc4j7392y3GUtQoNF/nOCGo3DJsbgZvEvift3cf93Z35yA+/tbY+/jNL
88x9gXObgy4SWsaqqBOl+Vr5yw7utxRpfFsSomIMmqw7MlevobR324Bnx3AIFKTY+bHFh5dgT5OA
j7BE3Mk0/ClnUz05Aa/Mjxr9twYpmXp8rQ3kNiu9Px7C8aIiSvRELKOtZLUECOIMGuAJ9ROhgKK2
hkC3I5x2eddGFod9wHD+auakHGsxrIxIU9Ds5IEsZQpz6mIHmRWlcXV30gDZBrdoB+3Q5poX3DEa
SWbQeUAYdl71KT2ti6uM0+PHw5W4fFrSgfXlpglh8TS9HEK1tKgfsl8pnvLpWOg9a0/88SeTkRQ/
NNysTwcyZEYRLpZ43CkXYYZ86jH/FUREpGT4R0QdyIfWjiqmC7QPHOag9hy8OlArc3dGuI/9QwA4
x/uP1rZzvS2UshtYDzxdhPzJhO0maU6CpXAYQPBKaJUIJwv4O/f1iby/y1LQnarLx5QS8CMQruW4
wMwEeZUv6D5aOAR5VSl1tI1iLoY9Q6c/Jd6qMrho8LAsZy9HP1/A1Kx580KAQMz4fU5RqKNMgwFJ
QYVWXKX/fKA1L//M/fk/2tkmGuFrAZhWy21z7j7HKXMSpaO3BcMwBfqSz1n/BVloQihhzODFh4JS
4SeNYxyL4OY4eHteNBv+AtdbfBzwmke8a/Y3XxSTmfAStvwKzjMu0KcQLb7jH0zK+jNeKKbFOQrz
HHekVNHPlfKoZIlkATi0iGUZ6G4zY9gdi9KTMk4Lu0YVoLBK3GRl6XEHIiQSb46OwPRv0d0hY2fT
wugAUKsh3P3XzsaNivuP+DmsV82xQ9AWnsZZfZhkI5h0LF0hbsvQ3BaaUkBg/mXastf+6Sz85Dc7
oubhoU7LUKkUysYWBWE9jdPIor5aaMozJBpFwBzJB40iEalJ/us8c4BnRpYIKrog0Y7BPpyiGuHi
ciejI3vlTAZVMinxWm8maetkcsxPzJko0W694VBjGm/R95/tu8uKHB/oy9U48fRX0EtR1AVOnWZR
S5mbF+2BrLb1vhLNhBAsSobAAnPnJpUVm84il9AJ0yzXpIaGhRXYpwQ6MA1u8O4RfdRQiAHy+V4w
3Uhu8cHf/+TbVOUONYliP0g4zJ41ipMbT1aG9WNmzgAVayKFJhF1l739KNdPIEEZAgol67YFqN4Y
KYorfegnjuOV/ZjlO+Z6M7j8J0bFzlgLg8LXiYqGTkclZuCGo6XfJqsSgXueYALdBzHRTR+yq+/n
dzWSueXpLEsDmlcSHQZ1WSMoUP5NMh4RqWHTC3vzQX4fTZ4nCes5iWpNYOLewYRPr/+JPIhM4iCw
apXQ5Vz+1vQ4nMZS/MDWh7qkj1Qf0sv64uL9m/fzfmsRo4F2rivJf2uaWqQDKYO15mHd6gZXfUwh
fzM/vWs7opH3uI1YpC2bKlyKW9ixDlaah493x5N/ySo4oyeqrBhaxhRqg1bAXQEtaWNM/2UY4J+2
zZ/23JmmfpKgfZVB9jTsm+zPEzXRqeOZ1FuCkTSu5ofDALpasmsglcay9Q/0SEoIG6lG3i9tThQE
JHEmQDDquITub43XdCghzR5NZdT4UCdVferVyqUf7ZcMEbWnsn5IFcM4o0wJnHqXSyCIrYs0vpi4
hj0T8GBIaSh5wmfot1KZuTDl3WDTlUAF/9qWazYUN/hViNMYmyrqU5pJBMard0S+gsAOf04bY05I
+5toRwLeRhlT4Ccq+rEu0ZmLN4nEF7+XnwK0uor62orSDhMceGggc64bnwxIBQW7XHFBzHNWtR9+
BY3wUi9qmjHIbPx0jGMeEjGVlSUcta3MaftugrA8dUHwMIt49CaBIHmTW0i1V3Nr+vn72mZKE5uz
Cf1rUUd7S9/SMv7DcidiCXNTz3sn909TVaARqvCEF/nitXCv3cDmKv0DhA63WZu/8mUJCn93RiU6
uysJ22RZ7QtzyDlFDO2SX9LpW2vPpxOpO4IaE764S3HXJwbWxJHUbrCvVaOirNbXaavirP/RUqz0
q3Mkn6BwFfGPOliD1BAED3Ki4JpetABYX6XDeqzyuT5+FX1c8UrX20jrBO1sx+h8yBNSAaJD6vMd
bn32290aPlDfWsKhEYpOOhghGg52fGK+bDKQCTQIS0OZhwmgjm4wL9eGcXtSsd3Dmca74HB+i9WP
F1TpovYBQV1YthTMnq7IKQwFFp2QmnaLQpLmLThxtmILDLhgQgRbIf2a15gfrWIBuonEiFRKnsmo
tAsAx9Xxuo0aW6YV10yFpUpUtSg5b/aHmqenY6tgjnhWSRdHU8w2TZCHKlL4E5AW5bLKBSTGl0JT
02wWk9TR4das6x2mumIxuWSvfHUmkZ8Kgg9Qq85N/kGSyvTQm7yHgBOcJOW8wrZtXAfaqTak+gt1
Na863+Evj/FhmnZ1J2nBW7AmoK/hIY3kwqT7yrQaz8DfGtuC8tDMtU4T8BOInX7ijh/YvcEzQA6R
jsSqCpfCgZX7hPrnxmarBcxwxpPT+ssQS2+/WuISFN3ZqtUAtcc2S/ghOhFCNFVYuVC3IybhfTtl
tJKX8hANhTfcfpU1XiXix+KDccQ/nhFJkLLOnvcnuf7R1NyzNJ+gLyprHNvJpY+rDDHbl5J1f5kC
kebK36nGv39UTJ14Tp5v9nxrQqJ4cIQl43phqtHvTYQfJPmFcynFFndLuBHdC7r2XGZsQKEPhSDQ
L1AAfFR5NrSBSsDx/JwTdp2osz32vU6PlagKaySC054rGAWjfDZx45M18AZqDWGLQKPuPLDN3F9f
JdrapAYoCSRtf0r+MpL50eF8RuUZqIgJOCWFYVpfUQ4SDDyzb3wILexJJxX2hTUvT+sNIf4JNwPj
qs4qMKBGrJ9cbkO/vehbspX0NveQLL3dPWIMtwn7si2YG/0cwS8I9HDbKVNQwwREq9CY6ikO4lUi
363qV6XSH5ErpclHS5yISSrHsWg2li4XBExdxNaR9T2vDRoUZIXi/oYG5fcWxhNKwOpzsQKXRl08
8+fNUVORCo6lF0Df8DHSHU0gA+7ONBLvkSYmu7jp7gWzLSItZYNnVaI+awCQiVXN9VB5RL8yf0Of
EG+mbhfcTp1qgeYJjUS2861dicM/QtSKAjm3gMlF19Q0MIQWDc2S+qETlHAcPCVmUtAK/F2Gou0B
GjgVWiUAsJ9MGlI2phExcdOB+Fua1YW8hgOk4kiEjmSxhokUjaZOUiNVdQ4XBjqLs5XJYTaBm/sv
AZ6+Dt+eWTEpLtCMftUW6V5hFmBA+EEERiSQODoe7BGUxmayunOpuqGqDNF99xHI2yVONp3A3CkG
5o6lv+7gG2olKjHzfdmk3tYIGyFNk2Oj/gH8Kt0rE9bVttz+FxnJ7h9ZAG/dVzgTkXeSlxDA7KBI
+SD2Jxl1v7FZ5UnnsxuKLOkIr8e1InwiuRcvAqbfyUW8BU0aql8a/YDo93vfn718fQiiA5d8T4FV
a6x5yQBQZ+TO0hF638zWmR5CojvTleF21mPeUdAIgBQYbWcToBHdgCFxe7LqRS1fxAKGp/tlTn7m
hSWieiqgK+NjVohkNKx7lRqNmB1bWesVoo1rA3gsrzCojyUxt1WY1FdLsNzHYQxhFvAFdTlNGfUn
uEXSlxjfnP2A510Wm2kQZYor36GTHTol93NsxGgeI4O/mmBt6Gm2qIgO5QXVJ0NFS+MeEvG+KiDQ
tOaK/nGzFH6eaqo5bbPQ0TeFeUGNO4iPNhC2QIe+NTj+mj6edDVBXfumqPgH82VQWnXQeLYqZlj7
JAiEF8XNgcnzUnmMY8jCmLQMLJNXTwHShe47K0CNVSGLgHofzkpeLD99T1OfdRXxqDMnTkWtZUcl
6AMyISU/Ag1dDezz0d5cLX+ZelPL7jIK+bTrGbNbzyRb/xs2vE9caqM02hx78HB2kdbTcL5lAfHt
cv3KLK6vnM0FlFlrrIVL1sks5tnddbM3RzpYg03QADGw3adWvpFdJHO0rCx+rWOfbIUC+ZZ6XDFk
p3SG40d4e7QDR/WdEGvmoolor6cwyyR8mRG6g5kThPUoX0rJdCzJ0kQ2mQDz1O8ngW/M6hqLHG4+
JjZ/uBJOi0e/U0jFI77WcLKWZrdjK6g8UxKOeOI8TCrmPd7YGLcDfs8si4OtVG1zvbO7nP4XTaC3
nODv+hKY6DhizcLblssGvlytO9QmNdx6sFuKoNtuBSQiIlU5J7D6JDvSzTXxrOJOO/Qe5edOOIwj
rnkrhBK6/3dbVGs+Ima1F3sqXMLpFnkHMIpgVOKJJW9vkqTabDNcoxt2UKXNN4vclfNUutCRTeQj
kfLeiJOLqUDQF6v2ibcGEVVbI5NU6KVcq5R26jXmVblTCAv91Y4ND5wL/oaghHN/CAT1XhslCAdc
SIOA8MRpU2qUky9iLkD87RKiA7Cgr8C0P4ttDMihdi91BI+pitzFJT2t+urXpVaLnLNPmb8v61uf
5KIjwDvdnRBLL+rIAx6F0PqrJcp+VJteRKXSB8bz/6CTtixqrGNqngpyEHFVFV93WKT5x2sMaG/v
7TG8iBIM4Qjq5Wyb4sAQ7oe1sMeveCnWnsskqtBsgDDxC60qfh/8+ys8xlztQK0QM9ZtaI7DvA3w
UfdYgyae0aNuI4Ks1NAlMQTHd0I/oyRtiMyl42xcESkl2MHCwSDdl6xkYuwOntclgP56c1ff9FMO
bAXya9dO/m0KR4ljOKq13NgNIvIGYk+9+NeRQBYrOoHr83z0g2E76BRLtAYIMilt49heUrXHGvgH
URf55HJ+75qAdq9yoEirZQHivZKaZy6cuT0abIk6lsAZ7sbiB17zbI/8vI/hDfFfkk0u0T68BElP
uubu5giUXu4se+cQwWLLJZr0C4YZNrFxGuZAi3bQKS38lYZBHYesp3SAfw6she5DibPuAEv9b9r5
NRVV/mAhbbR3Y0JnCcbBeLG0GXJsVmUKS0AdsZl7dgNXe4yA0/xOClZWU3kQ4Fo4NQIZGg0/hZqU
Yb7170Zsg6OSfAXMAoSlr9+3KWzhz3gh3nDYJtJ4BtFXh1rfyz5YVWH9Nsq0By48TvAyN8/OnO0q
8o85Diek3Nrf8kcU41cq5QTcjoNn3pEbLa7C4H4x5JTCFGlxcBpW6FM0jVAtf43wz03JJYeasUuy
T52Zrf8KBsw7ntKV7c4xR+1gtZeEAcjaL7W8ajTjQHTvmTkOys6w5i96E6NXoPyTW23xSvdU2goM
BIWwHxCCBEnzhfapwKg3eCtE09OyLU1jR95vwQsqtdzUgjpXVG5IfxcM2A0G+j4Ipi4RUQn/vmxS
c2WwSg3e/eK0R1Gdf/6QUgs5HdUBIYchgsux3xUsiblOf9vuUlOa2pDKiiaYza1dNrnszy/dw1nG
rp140sAKqcde95DpKZWvqx0ZerBHHIHwVJqKGG5OFyVbGqG9zXiAqleNgh3T4h94W5DL/TiY5evA
Jyald/25rPyeHsdVK+FaxwhrsPwGc4eFbSanPO7MLo5fHUM9gSxnR30fpDvSD7qollBiNeqRKhwV
wpKGyKVxLZn4RqPnqXpEpfL1KV0TFVbFpeBz+e87grrj8q8Aixy2GXFd6Ox3y9Xa38WKPWxDAtZQ
u6zprcFS18j0fbA+Hv5LbDm9HvSn27I9ClnwiP59Al99ndwGnLacgnA0llUnApCsZ7fAhgvZovwU
Yjj4q5glXS27oOUPXgrjbZ4fLJspbaLr8NPa1aqV3bglSrOAokzKYTw7+MwfbmmFxQHr3rbLWkQQ
jhlueMF7xD7WtzsiXuFYs9ziwZsL3jtMUHzWVOYb3Z8ohEc/5PlgZKSSzWmQf/fB9mg/uIWxRrcU
pBm/rAfkw4sLBo16wYOtlGvf65HuESpQAWmdKDnYSPWnxcNN3RYMwZ2njHJ1yrj2DC0RUexGi4Fs
+gzquw7hlc5unUhD1UqXy3EMRk/mr+d5uGswn7/91fxKc5qGxpCdxzbAqWjVReTYIvoyGw4bQkSG
ZGQkLix4nc9YKRepTfcNq0hZujYQwex/aO6tsfeDTGMLaTQnpbZD/buLaFHpOGcNxDAr8TXLFot5
l9dn+T4GtdE/lOJQ6Oawypg5IARMRwLhOnA0Xttah8MXd8CQLIqx2jo/zjDWGAogOmNYVgYVONz7
vTDds6RoEZzb+fEPdCpz1EI4Yv6jaTHRGEQyRwyFOY2GQOa7OPFlpr5qcbEQzot0Ekh9KTxGx7jB
osjLcEImIEd8cAFvjIwp8h8fO21KEB6/jjDkyVP8M5sMQwZMmXhQL3TtdI3g7mGr+Ul5C/LKh6AA
wRtXo5Z8wHEYasnp4PjbF2S5AKmGWQFNueuWASuwZ1q415BBFUJxDaJAKIf+IRK3TSL3WzMH2etf
eDZ1V+5vECi4o72zpPbHkFVITqhMkR188L2HHV7HRsS/SwjfDYx0VOvVpVGSp8uLUldsYUcSptKw
DdWB0fsGLbhm4Xf39m1/QxEiY08MXBtWHUWUpQbE2WzVy48npmqUTkCb7vo8Qs8hyWC59hgr6Ruf
kbFpif8/4f2ckJz061kUi3ovcsQw73pQaDocJBUH5IFIGk9QLTOuzgbGjrkrv5w9mx40PbnEVWNI
+PHBBxianvB5Y5BCVJg7ZCR2ETunph2z+WDhJeRTnZ7dEPbh94jATZYGIK5syutz63TRXdlNPfox
TlAERtCFGZS5xUbGHoMRiM2BFLnStrIjbM31RXU9V2GExUauoIsQwVkKKHiUDXUGulNbvAWRtR7p
veBvE2nSr+22ltVqnhktVEuYOnvG0WeaN3v4UXCzHCPsC+LCducn6yUm9297D2ZCLqylkXqhM+JJ
Wtl+5xWwdBJTXmWN1nPtj+NJ6ATA2O7g6kIP8jKeZCLNVwswJJJTeRvCh4S4orjCrL+PrdNVTKZu
Ti1lln0SW6152q+mEN6QXoL4sEUn7O9Ko4alpUhsK8UYJ75L9NOlu4RXwIVIApWylaQtuHKiqV4q
gypWnCB30BxbPjDMC027Qwh6+/2UkzPjUiG0HpixJtu838G1nr/7eXMBdXxQmfdSAhRK9EWmIZJ2
8G23azKsSzS4C0ESN2y5IfEkfESbEq/ycdk/Y+waznO5dk3PLVMbuBA/vFppPQGCeYZ9AZRVV9EF
Z1TlLJ8XSIHoZEGuYwq+XZyxN/12GAFbZiKrwTw7PhsKtvmCcpTfCxre9RpJ7qi8xauY+jCPiCP/
y/bWXpzhOsEr7DrvNkWpVfGFX+XrJiHyxNo8hxIA5XM0iCojNxZUyOLkBWtYwzgrobans4FIbYCw
qGBXy4zeP6AAMBjPYpFd4QkOj0yfnrU+kLcPE3yOTQPPIgY7iwh3wEo4bGOc+9brT3rQSf/zsyxp
zN9F5Tb+GafCZzRzO2OceByyK6JgB5gIKPR5kKhhb3038egNgMZE/1p4HduGe7zXmdqEcP9XzsXu
uw3I38NyHOwwpHH87t2rklIu99o31JcPC3+AQ9aWBKUqkEspGcRmQkDLIrEc2IMFbuCzzBMU0GMG
Lr8+sAoqQvz3aACG1AOCNag+OK4ZU3TwBRB59gLhKdp7aBGAslnPVchxbBc++3rRr3eAurruW+xh
oW2zjAEGSD2NUmUDxItz4kJ8lpnp7aTVkWGPri5StNcKaK/1zuXGnivsjmo2xdMlZ9taxtK9UJb+
nakyiWS8AffVrAPM/7SYD6Uiv/j8lFnMIH0DxlpY84Mz0JCJ8a/gE+mGIpKCXA3/83WSJLfG6WHf
fmnka5eAAQMBaOapeaXaZmLNvs0DT/TyP8CGQDdb2UcjX/fANuKg6wWqdYthqYgAkBbP4biPRwTp
bbZ1j7yEc4Sr8dO03idhGigOZ9PruS52kKcplCrldXB+w9GOsIJQvZ6VdTejhZlZch9EwwjW5hQs
iyGq3w8ECN4gwoCBgstE2tgs/Cd95aWU4jt23Oe8nikKmozBkqw3fNiB3H8isGcWz94WESNIRe17
BFxn3dTaMmTBpuhzPszOhsC8VxezAyf3wSWYnC1aX+CIXGj/0ZhMhMEB48PyRYwEZVDZAvaUxBOB
yiAPFD4jYHwNhgY059aZdeBFfgRI925sblUONVk7tMGmRZFGjroOgfzmM4nBt3K3OAvBQJdPTK3t
jVttU/+rjV62rsqkiqroiGS7PZfxli3HJRQ/oIeVpfWgHtXO4mu47rgnH7i5J5O/b2Z+5M4nZNVs
PIz8CCPpedeaZYMKIVfTzc5PRxGF+3L3Bcw0akVO6HovgiGpiS1bgDE8GCIPen2H+0h8R50wrTDz
4tOKoDSm80sT30kQaGk0OIULfK2oMSvAAEl+5qlsk5oFRhvj6Cstpg49Wew7EMBEYzJZP+w7xICS
mn22GOcdJYjn1bFDXe9Iz4tpuaD/R/wDlXatgABHa2wpicO2TWYoNjDcKAq7+cJb2CvJecZUk1xP
m/z7bXrwtBU70mP2IUxFcfJaJJjV5QHW+lqV3JQ23EnJlvmZnh3no2OLO5WfljcFYl5sP0s5kYKD
4o/EYvr283/TrIY3wV80G6IDqM6O1mGU5covHsY0QN6jJcnI9oP3fY2lX55HfVov8ZZfQktAsLxJ
wKovhxPlF0hzFcP5w6VoWjvupFl5LSiM+rEBdoz/UhR1pkYeZe5WHf75W7GhtchpRsurnjqREWvS
Lbo6kuE3dPVyQCcV02uHzlsmTIC0i38POwLm+kl6ZHVLJYUowvvcGWNv0tgMrWIyzwQv80c3PeX0
j7pEZc/RveMN10LYDVg+tx/kx/02fCV8zVpfH35mHQ5R1oqUL6WbZb3ImgCFcivb56SuS6xF45sz
ccj3XFdrWu8Y7ANFbY9D+zp3MNPoII35Jbpy6zHBzsrkK2k8Vh+lPCAnRS6RfdTtVCbQo6kUUXpX
93VDCDRYfyYaSMr0pcweH2Z4K/ZJTycNSN1jmjp+ZpV6Q90/Z/j7bBd2SQz3Lu5hFEfpD0QJXRuz
DFnlCf54iwib+0c2paxG5HUtpC4CcBam0WzdFtPAk8VAiQqcj+bQe/UjLHqgwE0Rg0Fk+wQIHvsd
oYfN5Ie4dQ+G8W1RmG2dweX82NyfuFZXSRGyizGq1nts9pLA8XSFe/AxrNHFZiOcARSQyedVmq0Y
D5gKFBRPQ0c5UOT4ndkUWBntsW/QU3EaeeVqiDmYrOKbwb2AejXgPuPQ7axeEJivNSWffmIOZmcw
BrFrSRuSXgktKua8fu+UHV1a1PqcNHMgIgtBZAqPrlgbZMOSoDEyIcALdU3CNksK0LFKRTaP8tpT
iDbgzrcHfXDwLM40ozBgZe3x4BpG+CPtPWWTIaO40N8XnnB3zArh92Z+prenbToebbBYtHhQz3t0
exEytdWqkfcPN5aWDGAq+6acLc2wXwh2tshwc8ZI1wrDNR/KPulcKgHwPQgA1d1+5DdicTmVCFv0
uooEjgya2Bd7G65OLu0KFNF4yJE6y4rzPMtZr/YsPa10C2qb+gB7ohMXzIY97ZPf63rtZVfIGPPr
W5iUBydZ0m67L3FB6wU07PZxEKt1XfAn/j401cr9iMCYIfb48No4OTrP+m5A1ENI1Cz/4HxhBhUl
I86emrDPp/GTsNWddzvhloYS4Be2Kmxzq8EbKZtPaTfRR+fjHwHRAgSFdSiXbZEQmPun6vpKjjN9
jl65YBeo57J+6dal9pOpW6NhggwZmfbaD81+sGzk9QznNfK6TsXrDm1ctdMMJ59KzOTNFDDf79vm
hJhQZV/+8gAPk2WqqtNvJGA9LH2be1hFDZnbXo8SvUCTHLMZlEGLuxGalRIEwbheScvwWrdSNOuC
7dVnWyzgr+CzwsgTqVndLEgDMCm01tU9aPXn2heC5STdGGN6R9xz8OjdgrZ9dgk553j+hgHtX3B4
5uLI2hXgrzV5vrS29CFXBpZcx3lLxWpeUAQF+L3RbgYz9ZJorX5OtEdRmdZlgOawaW7WPKYN8jBA
8jDui/tmjEr4gWbwyXn75uvia1WM1WgvQDugFfC0Tam+GMQ08gHfe1jcSj0OmmEMY21Ld/eXlqB7
lk1Olhw1JnU9mqwVPC3sfGbvnEBm4IOpJ4mdIbmHt+HtXGxjXJOM2goeDNvsIi5/ULwXD1yXH1dB
BeP4R03OyAJaY+KiDKqckHnGB9UrvAmwkrYTvSuPWBxd1l9TRm8KuGltUIFKh/HzXF2jgeKgSiSs
Jq3SR78qIrz6xlR4OzlcJXkjyQjfvsr9uzvdgQpTVY4XGhfqCY1Yam9Ju8VzdS4Ue4vNMJqBUv/5
/k+nGzO+9AcHdo6zX9iPgSPf1gJp7RVtiSSIgV4f/zgRIzm0mEX1EgyPiovLZxfmpIJ7rzYogmiW
Fd6ZpZtZ91G3m/9shxQU5I+MkcYnJJGPjk7FP3hnLFDMhV177ZbNSB2oiWbPnbRqc8LGrrzT0EU7
EKhrS+15IRmAGD+8RlQ6u18an5AD3l/LYJWYafGbH5CGjX69OZf5o/lo/ca9er5nHWF1Cw5ywn/2
WPgfqn6r4EtxVab9a7FB82EtaJDCXG+t5szVyMghPbx3FF+EP0JkOGs/f86fqDNc7XbPuERtvhGS
XQ8KO0fP2r/+to+yr6HLn1pyqLBBD6xvxTCL7/slbX/VVSbO7tYeWfSo2s8ULYHjXfGe2Gpyk5RL
/NA7lAqvG4pPpLdemOv72pyDWVbtfFgll36oJCkBdkL0eVxR23WY4YiD0ogMEzeBIUYupt6CDYaH
krtUB5a2wumAGta14LWe4KG5elpk1FKA1baqoCcrHCc66CgKlx0IQNjcveNOfQd1lnMHg01ahbGD
CHZPYcy8ueCIbkJ9mly4ZMwu8uwp4cCw1+yMph9JNLoOflRnXyDQB2UpisD3hVo+7ymQRUADEWm3
7W1IRZzFLyP/+CxTSd72gU+B/pbQ/iC1GdsVTc9cp6SUnq8XfQXulJ2SnNzKVpkdsBhB8yME0+3y
ImWbrZFSIOUuKOMxd4YQu4Wk0ojRKtTd9fCbXj6wKTQ0TZ6Zam9LNPbH8YOkaAVdEBbq+FETe6Ex
siQuyx9hopUHmxXO+hD2sJl28UV1qwAOuID9LhTfMBEQcmFnq/tbb0ri+Rzv2SMz0RGCt+cDG52p
qUWIjTaYv/Pdhxi1Gm9jq2Ke1SGuVv4LVl9tcO49GqAvRfeDNXlcqCRyGYEa7VEe07HGCjj2Yk9D
sYT8KYLu07n8ecOQaSTIEUwymuyqyoNeufnjS5GGW1Fgw+UZg8VbOXR7JS574npxksoY5++BUCn1
LkyUOqvZstA9YbBBG1c0Scbj++iJOaW8yQoCSFjKdVlvwjoICv65hU8uXJTRzAExpgxhL6i3/YHY
CB7PNShDZcYnFgkh7AtiNKEmZdi78TH3mvEFIPUQ4jT8FitxtqoBl2EWJpYQWv7Y5PD5s/KhN3rw
TaPOiXLwNNgKlHsNe3/TYmbe5tcqxrk7xBjJzGyDV6ZapQKJSkhNnGQQIrAJ2QKxzHtxLHCRDKZJ
CuCbYD43t2Q/Kn9niaQrjk7Rp8ca5tXV2XwBXksi8LSNN5wANG2IjlTWRcDtyJ7QwjF62QR9v49n
ytYAGifEZErbhRqwgFbYFcp7BNYWahdnReoiRiv9B9EItoKscL7X9sgmEVod6A9TplynM13k2Hwa
Kk8OpCjcLsL1qZMI5oQHQ5vyu+8CZKBxTvgsGEn/ICkQmdLMhLfzgdVkPrjsJiHAHKuAtM/1Q/Tb
pgc/B79kylOgVdddGRqLQHmtec4BWLxUFv3FRL/3RPXDFH6SEp19o5z9qJWHOvvmEPdva/ojrL51
iLAF0N5VbsBi5tySVjUpcjGDTuhuJUfCAd+vEfJ7rCnwNHQq6T1ODXnkFS0Dp83VihMT+aIMJYaH
Oujsr5NP2/gr6yzR4DE7o9YJWQhcO8p+ep/xbvCcw8jRTW7CjuYAfiDH0vNfLTVuEHYTDdlJslxH
oLeiSrPhVZYVlbD4dSby8Cl2nJ+kdIA876wI28TdAdX7l1BXu5VVcxYO0bN/4Plh+iBBlEEp8nv8
aub/O6+7PaDa2lTcKo2rbVFU9H7OPmNGjdVApFmUL6VBbWWd/SGoWC9GKZ5Na1Pm0zk9bs4oddNQ
GeNqCvdu1rtK6tpzLh0rKXBB2FuCoL+vPCYBbmw7Mh3jLG0Kv+eGxn/av2WqTCW3G7ugCoPa+rmh
i+2Ie37CmHwp6GhZfVrjeXWi+hf0alHl0G7YCH9kyPNRde5Nba8kzQ19PUPWeRQEyq1XobJntYLX
k7jRfHuy2G7Fg+7Krw+Usr9pZgoknXdYlfuJ+WtcJ2R4C6WIe9NDvfSAIniGQJb5Va6oAHd7xes8
ZZ/9hPXkz4FscSyPHkyargRGsBoHILEv27d67KlV+lzx8H0Zk+Gt4UaNSr1pEgHbR1Bj5kg/opDd
MmSLhDd1Xizgh4LrTW0SjrddaDVP75cXokMDcQsjrJqyiESV71giYc++sZSl4CdePdglF6szcsm6
7xytkkZveAXwOIBLnmGs73H7gUFvFAlmnTrVefBK2kODC/sXG4NsVT7JJnnE1N447ySvkNrkSp8o
+3o4IuCCqHcvZ4GYLVgQpPgAKOWg1qaRyoh1RZbptZsegNIlOrmR/RaKSPjnfq2GQ14ZINHdgCdN
TN7Otnq8QBISQOUoUb0xYqbmPFUqqGMeq3j+H2tLlFyf3lrg1bass8Q7dYJ0scAZDzjf/L+ty9p/
b+bCbuGUw3arYsBeIPjEjBk5O4Zz6Oj49fpV7hiwKWdiKEg9gdmDf7lYUaa9jDz802KS4DkGuMQz
jCsZpMqKTekKw5Ol6uRj0pBVq33DA1Bnn5G8CN4VuJXdM2xmiHW+WIhHwXy5zw82A4OnFOGPzmWf
SzclB7RcvlaClrz8uD7yx0JktN0zh4MKhg+sY6wodbgFBeGvyW2c07whNh7Q2AqLjPaWThhypJcs
kTwSRvZlp0f/yZ4m1JUBmmWQRd7LniBSWRWY8BYjSks9kEk1GTEVuJafJvEdShQihrmGsQeCclfk
cID1wBY7Q1d7YiTl/2o5OqD7lH1NSJXGSLzkdRUXGJwUMUPHLx06f9YAMUE0Mpxnz0jkc+HeLOJn
ymvKZOJB2aQMMm5ig+0zkEGoWbM2/jXApYmfV+EdBJPq2/UtlsbhgSgaLUsNFhX1GlN8eFuGXVZ8
uupT0mxaAlsLijTmqMeH+n98fmQGDzrottIs6L7rnZx4yBVktfFY/93DbA5QnqOrSP74sqmKK0kX
soPbKHBxq2MlrgDZfovzDYs4cqBcrohNoeinoho162ut1RaVYl2p+oLaezWvdayXK1B6FwIGP7oV
0YtwDLmv/i5BLFzmuaMdgeLsCmRCmYf1IMDcSebeBkGqcQCw2LjtvmJDhVEN6kCbTR4/EOgROUfQ
k5iSJ+xw2v5hYuHxT50+mb0Ygxl9WcTbuYCsb4K6TDG8gOVGTXddly8Ag8j6sugIXVUh8llAlPHy
8vCtTr0N3DBu72D6/vKV197lquqWSiraUNd3dezUbBRu8IPED4MkGW8EMdDSz7ZUrlQ3LB4wYdi7
Xbrbi6Dt1OviYw9arYxanJkGX5qJRlkbciMnTwvU9a7SUbeeMMRD+YE4Py1blE2d4Eh7QDAjh+4J
m1Bkj0Al+wxi1Y46YbVsRYTR0rdxrd4YoVzy5ywlbGLEueInBEWuoDJMxRMRYnscU6y2v3X6kZ1l
2RK59DPLsQvNG4cyRNyszMKs9+HxKw/ZY9df6vQspXtX3t3J/4d/oFTzVniZQhvElpJdeBu7lF+v
g+WOi2m+lYPbDgiSStVbcXLHuDV8Htsy4bKyF8plSHVgCAhS0M45bNK6SjZzqug3NeTMmOz4JaK4
kWOL6DGovgO7+Zy+k2/pLMCwtk0wR8d+TrFbnr2+hE4JDvIS41Z6cvtra1RfPdXOk5/wMWYvg1eG
dPIyqcLZGfxWXYrmJSJ7z7hJbxeVjkezsIo1E+v6MNcL2U1BYZcFfUnkGZu3jaebfbZHfAFUbZF/
R5YEDZ9aU3YyOhSg3HXMm0AKWiiwlHyjfErlmr4iiN1ZyqvT1w3Jai8yrZ68HB4tQWJ++2H1R4G9
xLTeUl7DEU0g19kIGEQ1V1ygPjVZ2A96dDgXHuIuIgqICsgTp8kPwQxJBLC0/qzC9ACUduAwWJpw
gPlRlnrKpSYtQLoscy38KndeYajdPyn3VAvBAJTZK+tk2XZPi9Hiyd+ws9m5yZU/q8SrJkUnARSF
/N69i2JnAH7wOGDwZ5eMhCJDYs8FBEb925BPgLRi/KP966qdarD2UPcOVLrG8t5NI7prgOyV5A4Q
sI+O/B0ezBgl3ybHn3vDuE+LUmomxhGYykns3POYnMRcKtAFBXVdmwIk+4jCSkjYLxbFHpiUVQy+
9eOlWMXtdhhBon2y1qiFW/nh0xEMR+95cwRIiVakY4mXuyQm3pom0YUKn3quytThcP1oXbvYNPtU
fNMEumWU0kZ443Of1stsvtLqJeUyjadXIPs2cwPxLY8Q8EuRU74yb/YaXMPAEctP8ZSqRCJihp4t
rP2oqoVpEPHOUzTK7D23rOtFRZSbjWscaEKp66yd7nuBzP/nUP1gMLtq5Jf9lXS0AuNwnJ93Wv2E
dusXePNtdD7ucl5CEwj8Ty/lD/2shxtB+imEAOfRV0S4YbXwlVtS8lMsjHSqj5xUv3nEEn5JlU9j
RS5kEWRpEyCejGnImg7hA6K5eqA1EzmV/FBWlXmtggxZqGAzok14Uh/4bx7UQA057Au9uAAeZI7B
Dn6qRolwxRZ/QUl4TfCUEI+m8r5cgPWSfK80XXFe5Jr/zSJG/fxKvaFNmVLtJVG5rXNHQswyyYbJ
2r4gkIajdqHPf3w3Vn+p3BA+QvX7cvlBaZ/JCcNL8pjBYpzL20kbRCcz9KAZYnx+Wsdl344BA2to
YyrAfhiNZ+XPdBgwE0YrDcw/oVMjMA7LdVfrP04rpqcgWhgshE4coBIZq00F5mc3jt4Bz6gT7fY7
fcg7utUXdMlAEIrL3BmcZQJKBasqz1JyKmUFpPgLsn4HsY6kTWJhE5Kxvc0LbIaS7Sq/ymLLI+ew
b3sTiEI5Le+JmxlyTDNUpULWaeQqVHzCN13IhZklfdoMWGGO2n6n86RNpADtCcFu5cQuvjgaNqRn
4etBCNG47bgFcJs4SXkv0ISaqXOuMGWNIrPizXF5K1OOu6E/Qk7lMpFLxOEkqFyeyB2GpsFgXdc5
bkcBG+MyvuBQeMYRVGDFTZr661cApKXuljsqcQgDM2RwNVING0RbVndkUSlxIlASlLNwhGFVOhe1
+R2vvkKvSnGrFyUm/c2Ua10tj98fReOPq6J1VpmiIa1cytD0BvxEEKfK+WrEvG+k6lDub+4WS4Ar
zBaaaYRG+IZUdzNVMubjQlj06+D4Q25G8wxIpIfn02oQYvpmWymPb8Un6L1yRtPq4EP4G0lBJ78E
glfdMAn/xXIa1VaZVN0B/GbMrPIxqbqvkfMv1ZFMkcbsEW9iAM2YVXVZ5WYlVz9y9PumOcDYkf2G
DQBRZNPVH0TOJ3aWJiBuzX6Cw9lPGltAlpl6ugRzh6HooHsHtYORbnZ/A17POIWieOCDTrjWpXIX
mDAvHJtiC3q3/gUZzfFx3OLJXsY8CfAEnn57XN+eYMdRNSc5wvXRjGT9pdvW5ZnkCPfeoBviciIj
EMurKE2IkuSbnEfwNc4PO5w+WmLLHPwjNcSnLTAq/25mduba7Zywdo6wgeq4OJKK/eXp7VR9S5Xk
beWnaMpQPBVPx5RVNXA8FocxTkChg0LnjxMe2dZOJLERpY4A3hFYHmtUg8AdxVJZ1ephdyRn6cFp
/nf0igLwrWmKsLrZfxzZHgQXG0wvXxfN2dOSwS6l0HR63UXqT5QerE7Xndq6f4cSSI7cUEGuwrwe
PRUm7UXXxYCWiLgcWacJk+cq5WcovjHfK/JHo3ARRWJoAV2ERhNzLwhSVRW2GFZAvktCxCe1dDT1
oytSiZFRt4MXQxsjMQi7t1hDNiFOddxmuxlPyXOYmbRk+tLRzrfVzN4gNpGpEwZfArAehvazqCOz
Zts/W5v4wm09JZLDs4pF7R3SfbQBU0yr/xq0lUFmDYUTdTMQ+P3hYxEkBYe9hk6IWMJGXA3Hpsbv
Vr1Xh/3wtC4T3w0rH7Xoy7Dta+0755ipBg2ld/lip27Bbim7/d60Ie0dnj4dNIEapfy1kwmH39nB
pDlKmnwRr27UhHHEPDdM5PrT7uCO7XfZ42UuqKLCgNFTSjatrKsd6+ZyZocGDY6Enwj1HeTsDZDk
PAKnweMSeW4Lhv3vjk8uNDGBtPg/iNI4v1JmD9Qir+6vlojY0auhysrfRGY9NsbFKE5Gwsr5804z
V79uYetPR0206AuZLYCT7i58aVb7n9banBBKmM09Zz++AZcmDjCcNaCQPVFyGZ7u/rWGX9zWUH0h
9gtZklm+k1QLhbk4PJ0tfssy0CYA+f10hZeIYX9zsH7El2y1nPBTxdo6NcrOExWUcqD58N5hpw3f
RHT4fJQxhNOMkya0M/1dgYgDuOhC/xO2P1Hkm18ZiodLYUpLFc/lfpEeatHdm8WnpifvvBnuPX6u
6ID3KtU2iRr0xC/uI4IBUwSp2MVz8/TM6FhLShU2C9LcIr6pqLY3FqNw7EoHni5HXoVNrN9N1V1C
yeUIoVIbzbUr/JLGeY4GyoSMPUBuLDM8i9E7lRBUiBu3EAPkew+tYzXzEW9cJcT7zW3zZE/UPSF3
iHrSSiiyY0ic7g4h4N2DAT5IoVs4XkHQY3NJ/RlWXf7Ba3CfnURreQuabwKFPt1Z2z7tV5G8DUNU
6677EKLmvyc84hpCtAUqb/Y4GD1Ygz1sqdKDr9DTnxkd+saxqgHTmq5y1KRoRSdTjQsoJcDUVfY4
7d69jPE24O+SloLN3fv+0L85+vNfca9hlpLDcfXnW+KTrrErQQ3OkffGrj8goM0qmQqDKSm+f0pe
ff9ODuzugqPm8GT6tJHI/Pj+r789wfyHsBCNuA19WNA7oUS+br984zpGONgv+rfWmJ99/KSNwhfs
oCrbOAx7yEc5zgGNSmtUbdiJpRPC6cU3qS7ShviiLLCnF6YuP5v85NvguUv+PDC9LpfA0soMJvbz
vHYGiX9xSanOPNRQshq/qRgKwcvkTIdAIvK5WgL4K4DhCNwaVkKuA99kPfXSHmD2FDFh7oyuRLNq
Wh2g58xcrjDpcaD7W/2I5+ABw1S1cLqAeCBiDY8rJlfLacvvz6UEuGNNEieRO7RrMCHdqJCmVQmp
S+pAFB3nAphTADxe4OdLK2cy4VEbC3MdfVjbGpiGNFZemWtxUlR6ChyH7DbUxTW/sY68F/rjtS/b
qJseLmQg9rSR4BX2uXTMgFM4VatD73NjWMTPANuYb/EHC5tcTFLVuMFwh25/VwE8aef+qkEbS6a0
ng1PZkD3Adcg1lZzqJ2AmWns7UAug5DI3RtlaRal81pfj3XRb1YpgJnSZWEKlFIt972DWtXR5IW0
BOG5zZUWHXQ1DHO6JCP1Ndr6oFuU3GMdZrcwYKvrOjYg5/SV2IONXYEPUfo5iWSdWdESAc5yzXj1
6xolfzw1QR55LkPIEEtMHmxULrBDkWimNHjyW9ltpoE2PhGoZYL64iwjciBJd4WrR3lqt2u/nL0g
uzLDPjLCbKlHPhMDmoUEqCWz3zJx+7T2qamoa9OMtPzUSaQZaRpCRgSJ06hdrfvESKFezfeqjxfn
zq3zzbGBGqMMD07O5Aev69NuBWIFbbkYpPQfU5fuB+iyvFxn1lTtmzALDvtGY7lJqlDnoncEOsEf
EHTAbLE4HQWy9i99jHgrmHsyxwAlhVnhKXUVscBiEbgCB2Loal/LHB4Xtupw2sb63KV5B4uKRu/8
ZHJjUQxB9dVHHDHz9wkTCuXIJ+D9U0Yin1kd93B55dHvyN9Ag/GTicofI1ysr9Nv0VJ3GkxOHevf
xxB3SQrJ7gZHe6Z5X0TfXqZ4UjLcRmfMU8vsSsurB8dhtRul/ADUR0fpsF4d0F2uzGlADNdfS6lb
z8V4q+hQb2pZ6KcIoV4E88dc4DcSjv17Aw1ulSdh2UZsE4Qal/1sOl4gx/v0ULMxZ0t9uSVcQzUe
iOOC8+xfZcQKZKxUQPPj88feD7fY10yckRZUEUtTndxZmJ7Z6/xI+r0cEsv7ZVApngccb1hgyFXI
H5VFdUnvB3Jxm8sADjSnU8Ls0vJ/F8RtW5p5nZ1X9/PiNIdlvgoQtDWpKu6fCtYvLqrVq4XHs8VU
qRJQOCdtTljBUVfQOEbM6k+OTeGgk6AvtsY7gouVE9bKTPEwU8Fgf9WTjdgc8xa1hHC6xQ9A9Va+
UGmjFuUiYZKOEM1TjSBERLByUEvfBZ1u2op3vPfVl9TmmCrRStj+Judqn+nl26HGoPaygjDh0Vfp
Z2EChOgdT8QZQ8rOA3WwWlWvqQYuw4B0S/rMVDzzab8r2A1abpKvt8lL1zcNWdILTVyzbF03tP1I
0HtzZMtpt36fuVv0tNImLeUKEBJSyVfAEn+aO/PfLqxG9J+s5djANFoku+LLdiss4I/WhMj+rHsJ
ZS1EILDTSY2Tea+aiV9XDwXDDZP+nm82xRg+STer4VRuAUo6qBquIfU7pzewE5gJslSC2XN3PO/E
puTCQbrTFF6Q+tAyUhTg7GRr4KXgIjXBRAPUZ2bllbv9bDA0Wt4axoRZnIgPnOjDJtqgXgFvwRs6
JXkndu+flKxh1d5xlizhatSrINmlSVEhwfPJ5d+OEgGcuH6/qRI5QvRHAmpWR1SnozBABrN0waZo
Lvrg0/DT5VzLridy4wvjl7gsdzdAAj0FFH/50BGUC24509mXUjG/ZoHHKSHhS7pWpVb9HAsBX6J4
SQ9eoOO0CtJ/wiJO38ZmRIf/iwbxOKQl7VBkEBOJ1z5wtZ9C8aEb1a3UDICgtmfI1ymcN94mrOeN
z0XXnItdq6ektBZElXLhYw+fnuW8kH9oEC1/FKsPcp5rza7kee6DY0B1npDyW/2iqmyIZ9qGZIjD
IDN7H/hbo1ANrYtgqITPGjOIQcJCwSqnWgn4M1Vb68v5U6Kk5HP98s96chrwpHgs+SAyscKj8Eu6
iV9voK6MJrvyw+oV5ow5vDXETCT+2xaqF1n/0i6EE/vGRU9bXhC7s3LLGEotg30Nuq00N+f+oVKV
wlojuIKKxxG/ciOjqIqLyebuH3pUKFPmSzQEwSvQguwyiJEfVT1qw3JqGx9QqHuOdBaZUa8yFPvd
wnK+xFjqAwCXgjKd09idWku9Oi05kNEyFe3xdJzQy9RXMVDFJI8AxzwdgCHcWoglwshGjuFsdu29
LdqK4j6r6FtTqTp66+pyAKqjphrCHAny0DG3ZvjgZNoAxfGfMNDVUPPRXkZCOokUmpUYxKNrAehe
2GxoXP71bJK7vedYNTiG6nGWpvKoZ2NXTwZivXkCEtXzB5I/EFDPSSydIaz4Z6ONTL1avt18Dx2l
TePWttEBhunLbUu1Dw5yMo/IKa+PtLkXQHE4X6sY153keIPUIXnI9dBgPgTOYAbaaDX0erpWxO71
stqinVKSWrunHTsmxKZWGs58bG+EcqNpmCIP8XoJWnxvlo6pixB+MHveaRfMJbT3PlkTNV9FCAGx
zS8iJ59oDAq2Eyk/8hb8SoyYQYa3TG/LiIyVgB0cwcLu5QDml6nhkBMj4HWvgJZhkIYWwFyCKV2S
i7kmKZo5G6+iktnYpOLzZfNFb8advL2SbFEVrNehxZ0yiw8iZXDKsjPVDrupDDkKUpIT1zPxQL9m
tiDijEPVinvExidbz8ifMQWsY6MmD2tG979gaL42ruCTCkoancHq1G4bRyZ8c9fxNVxdhUCIidK5
5KzG9SzVhiW1EK6EHPh4h+KlXtwEqIHeFOBwZ6nabKuYK55F1ok+Fxkzjej4KlVyBlw5DR+JwuTs
orirf9yGx3s66dL29xTZmqYiAvkixE+f1W1eEwP9huEfg8DBaNtS23reodedbMYLOp0gujotniLg
zYTwYmaLG42+kFB/AN5hDLCy+HjQk6UCRjHAFeAV7burSOziaLe1z6TxV1r8CfAYs17aqkr+Rn0j
o4PXMg0llhFosDNofPRi6Pfz98g5s0LX1S0KG6em3JMGvlgP0RcrVCy/sL3Bwk9kRwxRte0yTavl
ylV0Luw7LdfiwSzZ8y7kpfFefdDoJ6bof9PmDTqRCS9Fvdau2+EagPRQPZOoUIDk0lqkQlwfCjOE
Ln4ZVmB4WPvOnlGku7UeIBvBX5/BLUgEhAJs9Q9n9Rk3futx8pLfkXqz6sGlm/9Sd03w3j9jLcU8
h/r93ioB2lIuj2YYXw0lk0mvSY7+4a5jwai9IsdqoaVXnu1qVGTyiENiR+5xvCIizDavektK9Kgv
SaJBjsJi9RMacnXzaXCgErghQ3QXFnjMrJKZLvzqJHrf7HfMnuRshMWRSw8onOOrYYvnxlBscLYw
ADaLEFF/ftcXPckx0bhFabca3U4qTLQIBDQuK3pa1c61RcarpGbk2Vx0SP5KXplaKcF9ZbFBfrnK
g6hyAsuFS1EyQqYz5fMjRSC7sJLbgF3zId/WdGcfC1VMwtyrut41eclIUXOi9/+dqB0+bibz51X1
67dYncgOjauvx76g9UM8Yw7Uoz45SQvJAM1ks9urZdY7s+xVqTbomg+BoG1BZcFmS55BcmXJna7U
cHmVJHsdr/tux3vAGE+Jg8a43yVjrhH/+slNB9ZAn3rOZKoIfssl2TOe4SjVG77x4ACDh4TcW/Dg
FiAu8xg/owdg9JBdk1O3KbPEiufq7XORhwVZWw49JZVAozLnyyO29RH9dohFSFPsOTiRdGk5LLwk
L0lwgF6k+Kqh6u/srWiBZDrOz6mqMWPeut4MppiZ6ACa+mileJA6Il5hLLFR/XNWb4dRMJhTHhqW
FdyvijIqCSpVtdc4yNFtFPG8FZNRNY6iGtAXoSksXuUryoS6ClDbRaFIb9lKfhaPzojwhf3Cwnsm
SjejvhuVVGsG1NhgMwt0eg1ydK/FW7Vv9jnPjF+WHmQPY/p1FWSjRc9QF0Imh+sWImmCfx9amkO2
0OTkDbDrmjKJpnN115B/yf32DDoDF4NQhXLMvToQ1gFGUQOGlIFzeiiOpBoUSs7ZaolFqDW1CNl9
tDNJqvUG7eZp/p2E3/qbh/HLMU48dzH5YkeOwYtGDB1jxsqeHBb9sFFtYU+VCsKL0p6XH9XV68Rc
i6dfGQQ2nVTA1SivPkVfhq1qOdb2g65CyO5dQW5KWjxd/I53lNugBfyHoCrDMXAvnFIJWd/mgDsJ
3kPgIAeMZb+lDGx7txFEuRtt5XQs/iOH9bdM6Ie/cT8zF1RbPci9eh3+QbZcOPk0BWP8mZ1iXzEn
uAspeW+maVEFoFPPr5ZkGVWSb27bVibWOVVayZOzfGjUxpjmXukGtpPCyLk3Z8xSHmY5rgvqvtXP
hkAmZdSqvLK78+3e0N/Fpu1dA/rCbvInPC3TRgt4qMzT9br9cCqpQE4q0xThMtDIRDDkOgw64Ck2
gsnvLKrqbh/Fo9op49ti6mhjTMPJyH1Ek34jpRfCwDeC9v4KKlNpWSSZo5AgAa55BKBwCm32aXw8
PUssX7g+RQRrVrbtAF0KyEmAZmXWIUAu8onpXgcb460VaKhyNWT7hTQrXKx0S2cVzOPKxwP78UCc
E+fXuxHAIjs3C4+wtefsLmrQtrsXXzYMPLwhnadO4cxKj575/avtKh4qOMaGnDIVFvjiBHzv9kWi
QMRDO0dvFZQv+UKDKxc9l28IxJ3vc2kYAc0KgRYzJ7Bou34oFbiuZqE2QPHVdb+iJ2JgeiVm3TOG
4iWpnxoMV/oA4SLxy0JNOB8UcgVqLyKyXHUK20kt2opYcPNV2MfJ0BlM5oT/6hipwhn4QIi50OeS
qRyVh4Dw7z2dV12tqtRWa+RS9q5ErXzgW4cYGBVCni/Wv3JpHq7WqX761dVYY9dEVnnByURvrLTi
ruaTrk2jufIDW4WTNfg6t5YnJDAoHAOw1GlmhFrFxvKiJmRnz74JqzBB2TiB7rD0FQPDsXRe8ARP
D3w739Y7TepOTypO3+5n5qOq+c/VdfcmrkpTdk9/Xsj1HtBBCVVUlRWfNnLep4wstLAg28rK09M9
VljIdWlGdwIdQopPUS3iCNZjUrA6Ewo6mVNRmQecUvybw7XzVKEcR8mru9T0O70utQ11usX63ODv
JD1GI5BHL3vKnBR+L5IEUhqVLHn9q4KoNKROecL133Kt9k4zWO2fX5p97cnnAFqaf5wULNaqCiNp
i8quAYJTS+jar7h4QI2bifU4Im6lsZ2cQtmuFEsobEEiLs6bfl2/hErbD1ujQa+GJZpooY9Czxga
ZHIZgEvXZjYP8pRoj11zPbCfRdtvDTjJ0VEixx1xY7USENCHAKI3t7iOki5ZOzUPExvFqsZChKEX
mBhGTHNPG8xzURxWhiNSMvjyhLSPqkzMUAV0I5/qJsIXJad+qoejAA90D8HKWzJu89iJWyjlTlqF
q/QyhEfK3TpAANa5kwg/OF68QAmf/Udlq+eimcIVj+uXVT92wcAB44VsJZdMuF+6OXcHkkJSz+XH
pM92BCq8vG4fUMH5dhrkU6GfIdtPv8WxkNA4hK9ZZ4+tJKJheWGw/rGW85s8mTZs4boTw9tCXrWr
L5IFVpNGsrDtk1MzrNSvtP0po1dQ5j6tH8SlSaeuymBCNkPNo3v46qTip1/mqf4Utc2jMMX/3/9Z
lo51eC5I2kJHeKNEh0AWU3dg6jqgxy2l5GCk2mno3ANBgp2CqfBmXOkEO+MGaGQL7UfWGaE8Dlzi
91hWo1IgcJrwy2QbaDMW8b2Sclj77DS/J3DjViTex66jLmZNK+Netop2yaVz7hHKmY8IFzbY6ScI
swId6xf16gjJGupLVZou3YX0+iCS7zuMGl6BZib+5edrp4Ki9BQNiRqq4Ic9Q6gsSoZrAE+LCYrx
x7mr6/4KKHqdyk7nj/HClV9bvFa8WeT3ZMICoaXhQiJ2a30fP93bnK+D6oGKlkXSEV5IiZzwDWdH
MxNeRu5TtTTRITcYvuJKH8OtG401EqWa/5/CTbSdEAs5DFJLCCwlLgNDQM2JkohfHRRqS1Txu8i1
I/QejdRWmReMg0REbagwvyZlkgcjPBxiUcDRJ6rhs/rNOEvJYs332zPu3V9ilsu52KhTirLyhL2e
9/+mYRhL9Qhujh4Frh9vPcFYq3K0SrO4DtmvsOtyqJJpcrcQh0J5EmIPLkTokEKpnzDY7eln6yqI
cD/5ziV9JXPOc8qV5f1f3Zt0ieBVQaBQVTh1lFNMMyUtOTTUiRgYJdfYzGqH8azphztEhikpeGIK
Z+aA3WwH1pfGjdq+vgse935DHYYm3fV2Xko+WNDHLJen9ejoHSR6AX/Jalmng9FFIcO+rpRrNhnJ
ZJB3YWxqkl/jI4eAPj7PVYJ9jqdSh4ngMpJ2kNnFv5gqzhwXpcXs67veZMICLZr1DNWT8wV2Atmg
XslsN0paeFJ2Fa52dvEV7Kp2B4TlP+R4m20ufmoKtqsn4u2Ih45dK4gHdBYOWTMJ/HfC9hYPC1GC
M3wxdyHJnx2AI1C9lNk8pAeiV3t5ELO91nr8KXXOcfnRpVLZQ6J5MjHtxxcAnRIWL8wjEe3tZy3a
6ukm6aL1qhGQnNQuHnKmYXfr9rUdAIdLLJk8zBchiWAnWdvH+S7ILXjk7u8wDQ748uGlfGds7dxu
yjczlYYbnvcTiMGLPInV1UCljum7sMwH7r/4M+1f8mcqxO6f9kFuT+hZ60W7IQSfxIIvIDQdUIKq
dN3eV0KH6otQE5X/KPu0xBLxmq4QkQmVeMWCXpzG8xphWGgnTQ7RO7fRdhfdm/1kpVjgdZON7e/6
lg7BKFpjr45FP/pt4uTp5KxqibausUc3yiduSp6aru2Lm8wXc4lQvSx0ovkJzhFV2w677iKuL3/J
asfxJQ7ZfWOxAahRQHEyLr0AiFJsDbNpXEK6dg3TpKXgqGI1DIaG2xQgF1tAgByyPb7FXkJWSkGn
2Y4vJ3uusbKyIvzgc7UxaRP8tWcgQvffRaK1cILxBZBlc/wZ4pMaeN9VJbyJKWNUUCGgwmTK/FIX
bWk843VB5DRjlQ7SyUq1eNdcj26cJOOVjj+ZS6Af4QSxREDzm6yvtd2qyR5Pt0mYY+nyTEaIMu8E
g0axlb2eIbFLr4VP+p9heWZt9oJZdQMJ82ZdNwta22GVfUN2r8XQqXi0G59NduSq4Nx9pwrZeoAV
DxJ0HXtYQtRU5rDPulZ19Ntu0ll6vYM9VhWuU4AE+GDyq4nBHHPbKkUt/FiVMmwjL6+5C+nH1//g
Tj0Sw1g3EgMpJCIxiwFovmLMPLSOofVkuNi4kFAeJTYNch5GCTfYnqbdTddfvRYa9/RhVHUUSyGl
T9Btj/IU7A6dAK6cwVPsRBdjH3+IAuaEQ6kSvYb42LcCZWX+aWVrHARZldWtbDfs0os19oFKkazi
aBtHqe4GFKr4Qnwd0ks+IPVi/rsOoA5EqlIn/1FIjjskwAvGmO80FoktQllpQHuwagA9vdtbusrG
Tx3WPH9FkK18kqP5pjG5+22Uz/xYKeVdSts3y6Wkl6ipkJ/uR0vslLXrkXNw7VW7onsBCX9HHAvD
8zipp7qq4NQrP/qtnUCEvR/DsNysjtbr1nxxeRCu8sykPuoUsQQcU0LWfcwQwHC8Rz0IXGNL2Fcr
UNlcUjz5pHF5h6QY+6zZ1w5dM1oWdqV4isVLkCVt7V4jimXp48X2RiKbSIrx+EnbsIS9agtttBfX
o7uH+241Axfe9XWe28p0wa99fQx38+AqDIq2Rw+cWzamYf2hN/pRWwUHrae8Cpxp8r0p4s8P/ni+
Vu+mWN4NC9O7CnrCwgTySyEskZr1RIWmfg0Dxz24STLUH1Q91FoJgHoa904HhpOK5MTpkYK170Hp
iPQUIypnuvA6oRAXb2+GbdLuJcoxmSE8BeXTFfwWrhdUuxKI1tRYFdQEk2CptOKPAPfz9OIiMhU5
kqkm0rjphyCCzmzl1h9GSeztJM4lJiplAOiw1C5E3GwZLucYyc4jkUVI/MqkHGyQGfzZy21/NK8L
NTK5keupftzENR/PkOp7HSa9zqQVUylQ7MMfzBSbdKja8sB25OBviWZLzcY6O8HEC+SYejIhAT8v
wd4U8pLPpa+nxpBD9p2qQBKcCw2DuFSWzMBep4BPOdY9Gmyl2xRHi9PPWZsuDguJx6mt6Ma4BNio
jOnQEBHZ5AVyCrqfoJ2I8DX6E5HOu23H9n+sa4dj4+jA5u5qG45INdAVboBl3JHhR3lbWkaBlzYM
sXkONpeJG/Jo/5oTdJEnmFwwJGk05QEdwLBiVO94sq7grPswkhvuomqYS241fC9si994277qh5Ho
RtBdEz4Wj+FkRWpTrpHJBrxCEQy1MIeK362M7v9mfJGUfaJY6N+P7iLc4UZ5QoqQuk/HJT5nbXZF
s75oYFbqcApZXP7kw6b2fnYNgh6h1Tgyts3Fsmk+tLi2COfcZhMzQFt0fudQTM2g+WGtK1/Wei5c
Tjl/P0JK6uFnAi9bfXRf/DYYyQfZ6iuDBVTDxF6CJEsQvu8vXv1tJ01yS9BXwk/7QJyGLg3J7zTK
wS/J33TJuPVQJxnWdTSFjS91jKWAkGTLxQWW0HOX4YiW+jl78fpYhu1U77ANCQ9tun7yzwAWWLAP
jEAa0br3h7VHuaY8ubogoBZk1LCYkqAgHU7Kt3xAxNcWyROjH6nNak6RAOMhiS2lfJbNeMnUjpmp
k9sNZinz8dkBJhfzcI6Zjr1/UnmAKGMZuxcpN83aiI5zpMlQcUFi3J+OM/j7DD4dA5d3QoEZh8s1
2LpEzpRwUgcxOcCoBh1p6Oi+pVMYruBFFBNM6rzjR6XOsnWWd55bgSIU8tLyZUOorcGpuCHXfHff
zLtYek7P9ut1C//Pkg6z759Ms1TP/u0mOdqDCF/5/Pkd/UqJv3uN6MDrC+PfP/NTMB8N3JJVSPOO
MgXvJtcwN6WW2DZ/oduE3IBik4O2YkZ4q0EgPjvCp0cT+UO+yRreT/dKULhmPPu3KWaDPzGrFa3q
bUUqqs47KFyEgrS9wtL23I+wc58AzrX+MKscutKfznd19IOYPPCC6ReWVUw4ZS+KZdWQ0oiG3nKz
mquZ9ZqrjQVRrLJRUMf24cxf2tFJTTU7TB69K8Hxw7tjT9V2ZqAqpW9/VYsg/XA1OW0nNPaXHQpi
Ffyvg6A/jQNgxSSRyrTIH8wNL+CGk0onBjMygQVp2THyY39h5LT/HFJw9oO8mGGQ8z/wgUMhnqLM
0EJlIAazUCYnyDoXNPnsOlulipvYLw0xHM9jQqopJ2KbUw1/p5wbdpBmKvDVfGfVhZ5KmkdIAfx5
3IT/2S5y2dF7olmcvvDOln9pzLKUAggPdLREDmHRGLYKs/Alffwrvq5sGQH2eqJtNI/VtcpHaQAF
glTwz6JImLoPHCbTj741OTdY50DoTXZpYF7JfefYdHWV3u73Zcbn9eym8tkwLkdNanjoFAjsgBbv
h8hqlOXtpeMW9p5d11RWXoi2FJ6tsajMQujLgxk2ausZ3Y5VZSKTmjsYFm/1cspiYdYRv9ASSOLU
zHE8/X4R2DGIwKzO9RHf6qpIjqFP27nY19Z5PU4DnbHBw7Qxj9dJE5HrYEu2OhF98u0EnW2aZUFb
rQBEjNpVaKM7GWWmyx8DacX4XYPNLV1aAP5s+zrftoMStL5jld8ifqCyt5VhKqiIUzbuX+Rrm0B5
/8+TSnhuZ9PFT+aBA4fP7fM5L5h74OiVjBRVQ19vrM/hVOUW5FM+Jkz4LPEH/kQJjOpi62A1CypD
7m1hnOfBmS7j4aByq2YXRtBZ3mAtvZewSn4LpBuuE1y3shTEVRHXv903qWJ0qZo3DfbCFOygBFVq
oiyqoUlWFmrZXYqW96+LTSEw6TxojAQPp4yEcfPM+QEtM8MmIY+8LHKqA0kMf6bd1U2K4WqGAYmY
5yOcwOeUh04jOyj2uxAgXkcCZH3mnTd0KlJNQzW/AJzJRSxdp5jdhYOMF0tQ2Jjd9SNgG+2lsOMR
kaxEyV46abSFKSEDSY7epfJniJ7WigO53jyp+Ms7UcVtyaF7DBwTBiynBar4XH0GTHI6ZIjGZMso
VzdfaKFd+EhD8l3PeqgZFfu5pe+4xSscRJPA9p6wLKJURsyu7zCF4akmeNMD+DQfrPgNViSFcs8L
s4NuGSbLoReYiIEEz8AHXss336C9AYvVnNs4PT0fyfvoLQW2qTA3SKvYegfut4Qte56972ujnsck
bsQ4P37foL2pnWzVXeEuCqJl5w2zTxVIONnoU0x1kBKp0r5LSmCoqM3DRff3obt0r3mXm90hum9Z
L1dD6SqSkId62VfU+kMtuRj3S92HVOFHRkOeqn8tkH6vfSLHkGbttxeqtiWSdeHnbq4Gqw3AsvfK
ftSuIcJH1KbMAMRjmtTK9pzDZgj24LP9mKr7WlgXBuaMXh9CasUXs3mhJvBJrdJmdMcrtRAdJBQ9
frQoSOX8pAxkFOl0CCCnVh2AgEJELDQORoJE3DT0MZI9YqabwppgpICzmdEqGQLTBAjJonRCsHzH
Co/XuOEt0RkIPNxjUdHaA6lvJV+sLUudZoAnqxWbhVj5ISCT3/NcYcMtaQeLslKVn/Kl2fBtFx1M
QLtqtELbW4/oMDrjRPCThkWOgC1sxElwF23Pdin8Lod4Nq733wVEWWLoQpRWB2Ylf1hTzRPvu78v
j4B10Co59yIiFyscgMSw31CSZrzO6yjZWkPoVmGsUCFjjmpVtul9R1bx/kvheMqMpA9toq2wDFgI
UZdpjm+XgpVSj1W+Qkzb6Tg+Dv3lkkBnnS7x5M2PZKvIVb1ZT1kVKJWquiaN+d4W4L+2/J1LfJQI
DBGPlgymRHS2nvgwFkV2gGneTHyhTZLQT3ebX+J795EP2C4ugoSfhQyFkT7S5uYmQnF8r3nKF+C6
HyhVTIUynfNWYMPHexHyLZKL3/7vHi+k9IIjj86bX+UaWf64C9QgwCm2jOURx5CkO5i9R1W+cULn
VI9HxriVesr3IW2ZSXDSyXVjiaThSJzqCXNS6TYds3rakv/mrcCVAcn5PUG0+hLxyLqN8ieOylc8
WMT8En99SmEU5v/hBz+jvBCPcK+yPvl+8oPUFTiK66HAg9GxXhr3REQQlzAqjSjeSsI1uu4fWcBT
1UhwVuwnJaRLG10JdrJx28SYYja7j0OQpsn1f28pEZ+wtETQSJ8q3yLowEuzBYTPhl3fAgmgOgDX
SUHIIMkKupSwVzm9OAzJXeceIOqTqv+xx+/h3q2krOtqwktGLp32Tg1U5xpQUpYKDQ2cvBJ2eLCY
6n5qRn5TSomBIp8b1QKEIzkCfI3Dpitdfmq1GCD400lo8jHBvdkcB7Ju10ettRq1nYU2KL2obOWq
zphVuEorIlwMhssooaSZ3kjya4JvCx479IMYsAhV37EI6R1/vnQyw+uaCVk8wC4z58GAVzQYJe87
cRy5PNTRdMitT72V4qtp2ErnSQvPWfUhrKEVv1ySVwvo2Ok5syqXJw/i4MgEl5+JvB5t/agnyqFz
mRNcYftU8k1vxuKQJOcpzYHOBzzdINXs7us8kn8Y+NrDwqW+xkeJdcgQT+87nGk70mBVpuTFJ6EU
cWd+kVmydL3WcnlREaQUJwOxDp8JS0dxkZDBAwWfx3ukwP+gVohLuOnuwk6hqRXc4uOK7o8+qgQS
GpLvoVZWVbEo9DN0z47cVZ+90qLmr+6k1b8LXzQIt+qiRkscaLeEEtQG1VsV6vhQVpviuyW/SMzw
AQ/h/apJzVU/DNBgUUKWP9mCeXjyW+dpMgBq2gHxjFC5YHp/OFFioUTMimNsF81ZQZ9xfNsdhcjy
GV7BHzWhnVvgZDA7DGQxh1cBquFNMX5N8jpQG1h7iYG9uhvvCM09wP1RNHh1jEx/5k43CeC06KLh
9rdnVoP4F8cqkEWR37A+HrcAPlAplbH9h+PTcTqfcvpBkJzGkX2QTz8cUHFDIlWLvpsyQW9NZXXG
hs6AHnws+T70WUKwDZC2sdxvdiXoQ8R92C8u/LcITACvgGYbx2IP5fZ1L9bHqfFtUrRTzMeYWOA2
0N+5dEiG99dZdArntQ90rX1PaDDZ3iYq1AQUqpfAlmbD98znXPTVhzUJrnzmySEK3/aQ6vhjtRce
E8JYKM0JmmMNfcG051ziL3tgP+zCoARuwbnvFBv1LuM3woBlZsXHm2HunGHsi6+2JIz/WU1wRfDu
fukFT3Js6yx09oVxLJQSYSbNZVceXVOjr2bqagITo8CM2rgzJzmjml7Z2SsAhJbMh8j2FH39k0nz
xDlOb2whpwJ758m7ZJCH1989AJSAOAUsgJXDt3vf7avD8jmV3nr52dcBds5qlilbv3frIEog9/Uh
p6zeOG/JUfHGp9ZWeFkMXA9AESnGXZFexwZkGHbCx5be0HVWJnNDCZi9p7t2IPEZGuuM40wpbQvn
puLqbNJxKGqC1sVz0VY7OZQx4dbTJtvXazHMkMgMPAeicfOwgAcT5HfGXh6zbxuMypB2bdWM27cl
X8F6cEdIQCO2dpCpUEXkrCi7/fHYA7ThQ5LSFIkQ1u3Uw4g9UR3ukjJWNxDdVzmv8DVvqCOXThuY
iSFdhHFfSqrFT+8CVdSzWaOjshJfPzUGT8eNbbe/P3h4DRxH515idC6qXqfB6niUEzLMvy6Q4ape
8eSq5HIkK5nGxDJoMhoV/fISCZuN56AXbD246uMQ/4F15c1BYab6i4VKrQ4+FpwSH3s0K5MF+0XN
fLeubhFIZSrFEjLqC7jzfNzlCGgPUANKcjJaPtc6Z1bCriPbDtkwNEmB3b7ngIl2eNbycgs6/DEx
5Ycax+EH7zgKIN9ijks6w/eVPK285DgCykSqMpQfQUo2IweYbchqdxaUn63lVEXx+8veU5eJ6GZK
Fkkv/4R6Skjbum6tFDT7y3r01R8tMA4AFbkQ9dNWqFKzPG2PN32KZozY812BSvmqvY1NYgDxQBuk
kgtGM+5hbg/c2pzp/VZMoM+PBEahTquMBVTZq+UgLpDy6GlbczTsBJlD3K2nibxi6y3x11qGAo1t
qA7QprK+vxpuUYUSYQ7P09EQMYd6xEFF2fVoNTA5Jhkm4USXZ/ABVYDi/wb+RX9DAtub9BRk/TDW
pZK0KP0NMPXhsoCHM5yksH8t/kbYf0c7n+PpsGs+GYjVb358QaCC+J4dBpoWlqHLjGpyVc/XZyF1
SwEDxW4munAlYGWhRiR54wsa97fJXcZsrgypCLgBsRLwhfQo8H0Rbo4H0qZW4NSR7D3XkCElk7sV
yMbZRZKERbMkzJyh3s1PjEjB4l3L1QMF53+NK6hRCFrCROnW0WlQXuE+MKinZYNLGRZDFljzTUbz
ygSHvgs/UApfFvnuk+FJ/lnENZVWrexmKp0DzQcaGjCyLKMzs29uK8nuDCuGI+8S3zH/4UQiQBNO
sbDWW9BFGEtrPlGSlPv1ejVfDtvV/gw/vrmVXy8M+OXT3e0iUaSgb5oo7lEbs6JPGgkmJpXtx8S+
khVLqJpA34reVGEE3hRR7UNUq5srFPmKSKOOGb03hLuGV+WMghfEdtI98MSv1WOPvs2vViodAwmX
AajSNnMJ68crKMyQNOBDIv1fEYMcgsxCv8sYU1BTvPsAZEMLrxBR3+s54C1fF0AB8vuraLWq/gja
sEWd6JoqCMwyjCr6OoXi4TnR1M/LGEnM6ft6X6q88f4gb7wSZFu0hYQGyhprbddzQkAtpBPG7N1W
im+EWC46xjAdqEo+rELjv618Z3DSPAyvZx0/6N2RvqxTwg+4+JPg+zrg9bkGG3Ulitf7isURI+lg
EOTF3LGMrQGQYrYpWepaDayGFUavvwVI/zssT3ox9W5ESaRMdNR+JEvvlu8mwC1gkpb9BN10yKFE
oDSBlwokBXcP76fREL0n+IYmz0i0U80XAoOx+uA5QAbBaiy81MMjOHu7nqYzNTR4AwIG/d7lCzor
nwhDFh8rPebLZDZpPi7UdW8rGGQoPPhoWVHxapW5pdp2IdM4tKos9rN1ZVVpboi3fKwxzKhM5Px8
uK4+q/PW3EcI94BMthYUjxO0Y/DSxLPy3B7I+mO2lCMxZhW+PNbf2hFdPTcC8RZ8RZ3/A8GkoVaj
OOba4Jsf2i3vU82V5Np9aaQXOvBlSEBZS1Z0YWZkDyywFhHuCM2keBG5hbxcLCAYw8HLjOFpPaKm
IUTTSABNSVX4440j4LN3n9Vs1YqOkKoTOyubERCEqnHDE/EKFU+p+Vw9idNkpuYQ0s0AJxRmjgjZ
RPg2NtFT+crHq7sXXgmJEKj/PItdVifjzwUu/xhS2K4qQO7tCDNCm2ZWgFqpwJkCAZnAUk8mTZES
hWsxSHYrHplr0fcZBOZOaWSkolrs225J73FyYCGoHtvu/aisU1g9GHSLdl9XaIScq261JA+8ItR5
XoAQTduBnVRP9dKfMWszW56EVXWodZ8gKdEiSZV/46OJjS+O9Agjy0F+pEWUDki9Gc71gCB+nDAf
6FfzRYrBPBWfD9FMtNUchpWsHeKITfw5TMzDdTcjxF/fOn2So7rFUzZfAiifLYL4P394bBJUIoPp
Z8QuehN7ApXEN/FTi7GJkqGPNTRJaogoQtlX0v51zqa0o8LQqpeE9djh5dCN+xqu9WwjEXPEOy5Q
30NEoPD/hozl09vuAvMC6gkwaN4hE5N7iuYOUscuWPU9gHMKxD13RGZLWDVzikR2iIB+Y7RdSv9g
Sxbkf4M1J+x2VLorwv3U6QaFkCy8Mzq3QtyISd6Vq5oQFrGKYGpRnLHcvQuIxpiG8CapsR3pRRjJ
J6YgSpznijv007d09tHRXa4EYsPkqD0NBRsP5KqXUKYG0xBrlPUn3PUQr40ZJD5NIO6+UXT8MOBf
Y9AkujN8p2bn23AuZYGptolpMiUphiXeOg+kABRMIMQ8DXbypd088sZ6LhYm17M/iRyZqJP0FqQ2
kzpJVYCcK9Qq2UwAsXbZI2F9Mw2eY8G4BLRdc9Vbsq0B3fSPxS7MShvel0uDCbRNWAjL+7f0BTxz
QsR4Oy8jWptnvxFSn7mzUIVmpK0gMawX0IkNjxK2Ldh/s3pdg//V8Kh8Y+syeBjFf2B68lD+qYzH
C+GWaNswcVJi4FxNI3o36P5t6wI7aXlHxku3bWMFzJu68d+oC0uA0eItJZ3S+aKAsuKnRJ/7dVYC
M9URWoXhNDw/S2Lz2xSw4r4OstLP1gMFXD3zMSks6obu+FyK8g3NJDP4j2s/LcByroeH8pPFz2Bc
OInzEVMOm1gPPv+PihM0pzSRJGeY8B5dlA6bDJ0j9DefonWUunrkjFp/reOOnMqHg7dZgFyZ+tzn
1lXkUq4DpnMelTsyNf9+WVu050ksyW7ErJPWT3sXRscR640W0HtumOyCFkNyJcDNOhYh5R6dPZoW
S9Ex8wJ/Ma0IKbWPwsBBACFUhTUKKvAwxocIcuqVeHTiG4D66OcSQ0+i9juur7YoB8fJ4QxI4SKd
hgNZSX0k4VPBs49/D3nv1HQnzOwecyVm5hFT+VqCszuBrHwErcLQlBAM+yd3LcaevXrxw3BeRd9g
VX/vioahYh3+b7b8uD3dfT14qEmKVr65UZLkW/HFifUUZa96rjjlDRsxPddWvR1cSQQG6Dbg94b4
z5Omx4qKkZX0IIMfxTcqaxLSelQM/ZhR+cA2PY4WzwqnyWTIbvgNJY8p1mRA+hkJNQteATMyLei8
Hfz+8/VPLdQyb0M6f/fTcOHQ1H1SMKrZh/VuLkirrB3v+XTRtMljyxHS/hUzRi0qHHX9dN/bHvkn
OolJ8ww/4kq7HCoysCsNvBX9NeutynE+DWW/ldqWlIJr51F4XZ4q8rYdlJbNjypR0AtCXSOa8WBT
2mTMmlP5nfOQUDV+RNWRFASb0vEpqNQgPImxA/KQzDwObc/mrtjIVFoOq/X8NfeokEb8u9wBASR9
NDkfx7aeKGlum+nAarQR+J6ril3vcyNP3KG0oARBHO4MQJPfonXHu+eIOavhfccxJZctLhQCaV73
Dh7SVQ+xOk0d6y2LQFUjxMbQOynVlg85mRgXAivrH4nof7MpjMT501HINHKbmBeZkNfTbCJsGSQU
inzs3Cd8uBYDGGpfMmGi3+cK3vP8yxBEvfzvTKEz/12X2a8YlrhJutFgHdJAr+/EYvO1UVBquyl8
1MupFf+VeMIiVR6ETwP3YBxPsnQ6c6s/DmVLuvRC1u8UjXxC2XPbsBLDTdZ5UfAnHNZRtPvXc4/2
YJdt7gkkhPXG9LokNMcyUJAx7FwpZEZ/lUANQKuRaSEyndl4DpHQOMpsKZP+qIXT2XMFjXqknc2h
GB9Tv0pSsWZCiBzYH2R9rmBlCD+IW1d2nuu9Zxixp2hKGONlBWnpG8ynQkZTknPwLxUBq1tMv+le
zixhytlBAMTXVeCqWAoA/EmDPqdstMTY4R4VfmkF2UdBJhmkky2GS/63ya13Hd+i34+2X6HGubTB
dVD7wGPfbp01e4ZlqhIA1GFaNk+osh8xiw7EPrA0NPqwbI51k9IT/IKtrbaMuuj2JlMBdZOOFrO3
be+tnj4IrAcO2vgmLRF/PVNoGbUjWGYJdNQD6OuTY8Bxv7jNzeqaWyQw7C3vYJtM+hYYwtMRyHPZ
tyw3bLSN/PyxUJk1JMBqJ/X0/sNnM48LZkTvgu6KjBrncA/YB5cKzJ5Ag3k5MEqy23ypWLfrjQ82
ENlG8O835mdFN9l69drT0lOHY2M/OVJEBdsUfeCs8ivCBNAkmKKy/RUxJOasRTl1T6rgWokGDqCh
+5agFe6vUQriqXYo2ztkZtAsP5+x3TDSustXVS9QV8pOvUZntyCggpNvmnZS4iVFhwsSr3T3VpOY
Rn6JXiS8xVtfPaVsBx+gBOVFDI4bpBxPU8cSPxz0TcuGD3lC55DPEcDIpcumEwWCqwu937biX0da
ipmaYW8V4dxtNaJCJ/x3GrXOBab7oIXMMtaKrc+5QfYUWDLjmydleuNx9UTtyFs3qJgvIg2BHfew
PCCteMYrrD4TWXEvHgusHo6zHBzYI9dNPGkV11YnKCf3hTjG6l7OdNXpmG1g5xKpRRosu2Xswx+E
krlMjbtVuDW5a2UqDohbQKYN6DNwzUYzBOSBCZK5BXlTWq6wLTHY1+77yNeSExiAKWzicIOPjaEx
YELsiiPtNUm390zjc97FO512BScprVXcYCLtUeE6USKvmsDDITBdZJg1gojw0vBLQ/eunXv0lH5t
SBSmsWdoFWVTw8cGgCz0bqaatas4xZd1RwsbNiSJrOlALxIsFI+fni7BHUlXsGgP6uW3c5/envsA
0vaw6e5Zm7W/2TeeGj0Vy6vryfnGjbgNLG8TwzbBIRjVUA/DIMEPO+XB5MGYax9XasS26fSW7zUz
Cr0rHtxYXWsykTKMlus/tKL0K6+0VPdp1x3KZ5QUynLe3XNRFClU9fCYyYZgKi5vch3aY+xdVeB8
fcZHdwpZZYGQC0mgZEktifJXY7QdO5/20k5uP1s2XdBIhk8fkS4j1sWI4ml+iEhn4FLm7vlr+V6b
8Yby3OMoCndcL0Q0nUjfsd/hx/dbZ4mKn7+Z7vPJGj5IwHN2TjVZk2s8kTYaVNiI020Qs3+cP0jg
T2zPfQIfQMikYKUdHdlc9i1Lqv8VxVdIhSnwbWuO7DRYmTWKGjHgM5keehQ6yPFNApnMPmd/fVoI
WOsOTUBW7PVc6EDofrJTZznzEOtlXu8MeR9NsS4j+aRwlg3SZwYU0+JAdO/h9WCNDbo/e/3zNAw+
bF/uyQKgVMk+BdYJUCP01WZ6ABMrYG/csP/Ql5V5BlaN/dCJdN9y/kgkXfi2VwTEWaHLvc/8Y7m8
WQnr4Mtei/25D8RKnJvzlmclilah+LPCjfkrfEZBVlU5qntithvSHSRaxYiJpKTFL4wxVIfV4Te0
mlReEGgLUbiJ7Jyq2NWpfQIj+AdqC0L4N1ViwQtITnk9xpaccFaAzTo1PeNQjnv4ZksJS4PHzdKW
oKs4UNUxPlBjvksWyFULvh0/8cxC9xHptT56bMP5I4qNKDjVj+2J0FUxGHQyQoYqCHaD0hv1YX0L
Pdl46EbVA+VYIycIGNUZJM4m5bQ/niOhDc+I7McFmU63OyYjc8Of7Xtj3UZap8Ak9N0H9hKPxDfO
QNXJPMo/X9MUkscIu422HMKT8AL6gFROUg4LeIizw/6qWYBo56+Gl47RRZ3ue7Yq+lxxwV+kVfA6
WFrvCBA8wIqz4eN1I5n7z9I1Hmh7MO1m10404yh7Bo/cmCp3cfqLqEGyCzymzQOPJ2OSdDPiHYGP
UbtRZiV1keO8OvutQTcmg8JUv03Fsoy6Wt+ZUfkQgTtk7CRLqYKBLQWsvdXaglkmQZkYE/Mdchqh
UXIvml1knOX3FBoOyeapERElxhQVgFPE/mKoR+q0TjgEiuqF6tjRNq+R1hga/NX8tCRu74yUEmAQ
7rXDLgh2kgvZLGDAL7L/najwlhSDHW24eAxKP9gAyowAz7nK7cUt0IuqbMPHFg6c6RQI/08d0hEs
H44/ZLJgODWEiw6b4NEOUionbszRjoGZOaWa2KzOh3aqPtKmTJZSKnqyqJSdw+aJGfCjpQ5yF+Hc
gT3805nwy9yszmCDpHqvgX1brkcc4d7mcRVYF3xoS07m/OYDHJB8xLuc7kIZ5VWd6YwjhJ4UzLzc
/35vgI8awl13Q+Bec88fWObfab8MI2RrK6oja/oD5mntDkCAS4fLkHWhsa3w+jMYaBZYmrS08vhW
+Vth0YPOH7jguUiD2Imsmj87HuvPWJin/eDokFQTESYZHcgE5AjX972omVvMd1p9hrmmAZKcg+u7
vOWMVrPJwoPrHBN0DW9OE7OoMR4/QsGPUdfBMX1BiH+gwG84bZCa7gKzcsYBjCPEj3F2VBNQRDWp
21KbwJE2mpI/jErCJbbzldntALVwDX28rPRPRC8Su1mcJgmqq+EojSLI7blVzJMmOX9r541bOCwB
/tNRnIttqWlTg6QmyavFMyuRsA5x1IFPdc9FqTT2dLK/fOJEcREMRFva8Y5wPmNZze8t2F8F584P
zajyDknqBBIx3quONwHsMGqFx7xvFac7CYzZ95JdLrJdwbcSiHPyEFkJuMhghLYQYDMSyiARzxxz
/cVLLLSDpZa2DEXHgz+KIMBd87hgkjfYtZ+o/PJhUqRyKrtAbKS0KtN/6HvyQ+W/uNtg4STmgw+T
GgA0h8rE9D+ns1VgcEE7XtgW9tTIRaJ25DUDVlVyoxzhIyWMKaMYouV7tuy28OGfNQFBxNVqY9nk
E0zWWIfYNal3r05eIWnVpltPvv29zqMX+kH0BQn+k+rRJlM2SOktzoKMuj1s6ogQhugYtNtv9sWG
8WPBqkuFdgURcqMKjMZOB2Jh7VaQHVNFRinVn3EJQqz16giS4DLpSng2DKP3JvAMOI7Rg/HvxpV6
CyjmyKiJSi739FVWhOHtUBQqN/xnaSyNFScoXThh2P3V/yibv5TL03J50pAoWC7jqmTcr54Aid+K
asgdfacFFtZeiXu9AyqEgV/4/2bVkSCvmgB2d2MLjB4lCnidceQJdYOt26r4z5p1dAXCNBh+GU+I
KUJ3EvJsh3C6f8aKtF0w56nhNGmEzIICKlzcZlRPUGX0rBx2yP9TdPZCmlmk6DR4LGKEFFnDrZyT
zymfhsd7NcuZ5KNIGTm2EDIhStH6cFjcYqxmspJ1VjoMz8iB4UzMB/ivPYtpFpQKdAlQbntgrwf8
Vf+itcSUn0PzMkk6sDaC2l236c15ReFtTI+7Uf5DATYTlcnawVtEgFvsx4ZA8BTTftRLE1t4XkKl
43sJA/TZPw+qOO7SfOqYSwFKzBHW8Q2ibeuKU5txnobThq4y2v7VNz9XkIHES14h+NlnM1cChl68
vCKH2ArS4WOiwZWSul3f5UjGbPEQ0q9gf2pPnBhzbtSZgGnl2GTAGcGFetVl70+x7pF9NDVHAfVf
IxpFvDaKYUDNyYgg7ZK9XXQpx34an94dMltC+36I0RcTt23WKUBNEzrjRhJKiQUIIx5D68W76rA/
T2wEW7LUrkZQSuatIKythowOm8bwasTQ7EBGxtrrq4hEP0TfdDUE6RVPdkRGm8Ea/7AF8LVwbNXf
FHdlDQENDQegrmYR8V0J3Nv6NJUzIyhYhZIVXQCd/Wlpk5k535E2iXMhPArU90zVWmy/t/pw+IUq
AIwnERCeOU4wMVM806okl5Dnvg39MeBA0Iys0K6Fu1mKIzPk60JoZ6IxmCoy8Mm3dwuaUjT9U7GF
1Zr4jcp+jMqJag1jjlG57OrLcAX9tPgsDBen6VCF65jGx9gLSe3fLLHHBZ1TEsukX1CaM09AE426
sva5rPgWIqIR+9Un8mQNMAs437DZvDismanIlA8LmR0OPbBkZT0ABP5zL8Y8pb/7jQiwJ4RLOv99
HMmsG9zhHwI5FnbW9Y/QErdu7LD7vD80Y8QwAVchqwqiflpUfahcpbksL/VMP6fGN2eMMB+OD/U0
+/YtqYDe2ElbWZT6n5JSoYvlNVGqvUCcRmkqRXzCWCLZcaZdEaAudwMH+I8u59oVzl1VltOXAE7G
OlW/5Td8rO2u9eg++nwT1HDh3pkS+39dAp0gZKkDdwzp+ZZ6iXrjJsRejq6cUt68b9bcMMJhlnbq
2frUsipGSJPuPMn4+3IPPCMpGy6gdLi10AlDcBpI2Zok0h4VMBkZqAKwKuvSU2bJLwOHY+UNk3XP
78C4B0OzbiiRo2euOUfAMG+XvZjByNUsijaxR8zAjetN2cGDb1Ttkp2QLJhzLhr6ZUNUcxot97+P
AxSHsNsyRINsZqvN585/JIgzfz39AqSl9hCZsy6XmmEh7Va8LAHWlMfZ+1O3AoDNid2YiRCZgQTY
mteNUURkJDor7UqhpZZuzN2AqQPCQxOQR1Zr4J91pZHIxG+vVv0NLXDQWCqcNtRP6Ij0H2ghl8m0
xaf4j5PTylHIeffn9eVjltgmOSTGy4Wm120VPrxxcxkneaV3Hznq3jxGFh0pqIlrguc11b3++we/
9cZVwtiEleNK1EUuTLnR3DvOYAMaqbSqvwFiG+8ZYgmBSoDlqhcMaFAEQogPVvugPDKwxK4pcV4S
i7foC40ObUEr0in4ObZI0+3YVxjmWe7nClEjHWJEmvW23daShjEVa1lnkKIPjaL1aGe3DS5a5abx
Gc4HgJCDveJX1zKALXKrvegFwLpVKbrJ6qg4G8TWimRQtCFu435bddlUB238i4wb296R2PgFk/BS
thi2Ck+9/no3iLx7e4gdN5n80zIr6WrcQwfsLSB4EU293YD2ugh846DUma1OjFDkau79wbMl3lr4
tTUTj2G7B2GCNoCnpaoFa87vJIFBZWEnG0i5GceyXWNTsNnOx5VioANCqvmGJsVEVWxj3yIVji+B
p6N2iKids+WQR6uDTVJDMv/5PD+uZS0luw9/Jz3Mj5A0iypaGFiys9G4NoihKfXH806+OpZaQYrh
cgBlCvKc6Xt+PPzTAjpl3iMjCuaRLr59LWb130TwiwlbnAZ+aTHilkhpogFan7pKgPs+JzEYNsp/
J0GBOWS7wLAPZRtHFS/QsrSuoIRdAFMiAnPBcffee/x99wC3c4CvtzjEaRXRqGBXS6ySmGP0pVxK
nwJA1BbduJ8y7k5Ybf7+Xjsy0ae0TMhYy/nIpRswuVtt74IvF29DSIMTwvkFv6i4xBYInfTDpvEX
hekJKlujXbn9jVgZhdVUGCMtQj8BFFGhE+yC7qjOBm6I/1Kfll9/x2HS96ydjgigc5+mGFcJpbr3
1dJXnI+McvN0vReZfhU4whf+Pb7ru6d7sRGzkXfReabokmNrp4DdLck92qNwTwA04QpI9p3sn4er
JjCOcEO13j1MZCIayiUfVzHlkYf9njeUqmJIm7S49pwb6yH6VxUVw5K2wgoeitHl9NEx3WbNxNYG
3raUh9MD19GVDrTnF/sgqZhPOt9jKB+/yRS6hvDlVTQdOWcSZ/K+g8Lb37czT5K/LU/WJESKA0IW
ldFlesD5ycSMM4o2rFJMz+4oIgextbzseCr3pkmU4+YcOSy9164VmjTDQzwD16/dWI3hcNwUMr6W
uDe1SXoOKUwXPglM25/PBtB/ivZq3nIkfQz1dRsR/J7q7a6em9y8TCYIcd/nH9ne9NFpsKDmdBbu
cLDiEJw0xioU5rB3Z+XHmw6CRFLth1FeRjXY4s6/pm2zm0Njo+PWbSkP7X1aOkl9b2gkuVdZH6Fb
RrbJWJ1zX8YGxaw40Kp5IU1sILKORFW3wH1nLT0F/1NYqjpVmcwAiYul+V+d711D18koHz6346eF
HoC/4aDQZcYFGN6VveoQP3UPOi5q1VOpEPQDFn7yWtx51SWusX6dcbDYT2V8onbLEetu7onbbWel
MCe+794S43wmlJGJm+SVn2wD1D+5kmLea1+fki2H8Whd6Ct0XRckJmU+XvPbeas0HiCnqf6ktWxc
RrYeHNQFEXAcDBhmg1qjd7RinMq9Lgj2tQENh6GyjmlJ/vd7acX41s4obRTMWbgYBSRZoD1ImcnD
o95YXvR7W94XgD4K4QTMmI5cgEyhXIaSqpiRzk1kENuje5V5mJQ7r91HtPlXnTNtLwTJV4ag5KNj
6QBkvrM1KwpvtNpzk39hgnCVh67TgKfQ6KFMRpi00Ny9W+Nxr5lzbbf07+nmqEehRdJzMTIAQ8rG
NogL7TxXuC+lt3yCo29gaXR94pwKcaz1d80Tby9Pa2/1LaX50ulinMs9Bjw6WekSgBx8964/g99e
jCjvLDgGn98W0/DU81MEpGyIDidB+DSxQztUQX+W36pJvGVs+StuXIwarP0HxLf1R3gMq39kgJOe
5+Hc92YfDPGsOv72eqiBhM7EJ6E8eTpL/yxAb/cxAcBB7wpybwe5ulaLoLrbDR8h2n5YbhRbNkKx
rEkvX9Gua15S3R5zAzN0k/zqFQZuTxkLpI4Q1p6f1VuDfTNEzaTuRMCHR0F9ww0eRY2qI8h00Dwy
UdBzQ9FUPRiLJFFLqcfAzezpc9fu8q6tPZTqGRWT28NPKv5umdvh1zC5k3OtUpxo46vTyakxs34B
7oZZdVtytSEn+cUawT/3rq1uN3wsprylzNY1EZD+w5AmniSOLwqmFvcIfIKDsk9UYDjk4gzxn0ZZ
LATGGElw4Cvj3h0V9M03sdFaeiArnz+ZswX/311Oex0drJ51KcZ5wKHapkimZlr+vzB8UBlWUmqh
7tTeGIplJata4kN13pzSC5DkVKshK3ZLY1YfSn9Uih3LQUaOYliOraVeMtBir09EFUb3H0Bc1dU0
uFnmGQ0c/ptcC1WYnorsAUFoCOdrQFCg+ZCih2Gwb+8/JBWEfV+aiFkWPdMZ6iPqfVc8oanHkVgu
0ZNbr+/wQB2AGKwwyV+x0IOZ65MC75ltVYAIyYZDKaFZcdyVWS+2nAzJ5hdOt6bdafjqOU46KhK9
kxX/01sCbwCSR72jm4lwToEX2Ds0lzJNaCd5XfpiemVUjK08GzCDLYqFf/qB9qZtlTp2x4NixdtN
ldd9Nf9IO4F6xwklQcVV49dUr2pePJUdhvFM4x5/tSOTkkOeHfbf5/D6dWHkr18jfeDG26u/3tCS
uqUGRZqzPqXtv+r2C+7IcglCUdspENZs/s73MP6QQy+XMA6NHfs9v5wsJT4Xuj0GryETggWwX+Z/
28XQd/9CXXnKY6rgMawbbOhIr3RtimyaZXkwOAVvdGOpb4GpBtluAPff0k5yvpjRyG4HPrLLcBLP
WAdbvV57ETAZgLverfDqhba9XSfDVZ69zEXXYJGIEn1TSwQztSHgKCSqNs5k2KJQVO/tEyNPgEmO
tqZjzrSRXyAr0enr3BpLWTnRTT6zcvEd/xPJpCDpC/1aLm8NrofdiCsrapcpHDQxb2AgB3PVQqaN
3yizhSKC8znZlcDVF6f8SCJI236EnSQASwC5ZVccRnD8unnI1AkCYgjlycI8NULiRnvn2aIcmSUP
Gumjd7j9D1+iUtPIg3wnNBZpDx8kHGy8VEVs8Q8hT0wo4GBCpqqbqil6rI/L0FVS72VBcNHQpNrK
Ca6SM3pbZL1X+wS0bNGl7UOw/DocDY2TiplOBZFpV5AsDbtiDRb6TN7INYVy9WrlA38GHeMHY5K9
SI9nri9Hcb4j4rOf1tpnfYFMeD1OxNbc3C9Ej6JHNQ0hD1WuuLVwmLRYEiHJNW0RmfkeLOf5q89X
+Ae3NZz4DlMmKru71a8VIBUqF+SGs7eJHn2g/Jgvuzwe4reZKzCFAknNT5CPVk8mCmgQ8Dr3KOji
1z5PYk7TFs81o72cxGs7TpZf1eEmmyu2l9++drmsjM/IYFAZvdqRAE2NRDnjLz2OLJTplloMGnZi
WO3nfZhn8mkchmBmTBGnaWofY/Ayg6Rsxs4ZGG0ILlLw5a/DJ6cxO87lwI8h4ryl9tbHixf+O1qw
AV+kSEVkqyDdZJRqJxmtZcBvIe5UeowHycYU1+Kneao4GGJZMG1oQW4s1NZYFYMthR8ixa3Rwcfn
JBiDCF4SNIA76W5LCJfpD1R3HKfhBSdWp+Dkz2N7KE8pJ9eV2uGaux911BRQiPJFgu7zr9Z0sMfY
inoyrrzzvJyhULj37/dSF32NiZWaiv7kgIrOqWTRgZbJQicIY3GccRXxhgngj3Pcfgt67aCROaem
AqJ1cA5rWe6/JD7V8DPJtiMtbBYK8EtltpATO7XNhy5+yif/5F4fLF2rRKhxmtYcohhDMKMOkuiu
RSAuQUt6KIiYkRSgbVNm18DKaZlWMCRwPuSOVWk1Ho1iPZ34IWB9HY/sFO40wzmD5nhNLJ8fecNn
4phOIwDW0h6h/9XqUhEqtJ2UYJhKWyDdJJmO/za9IkoZ14BaO14TD85kvk7umUQHb1DNs24cIa+e
Pe8RCldehWzzRjQ3GMAiYKVAq44GwA1m+qPX8D/yKDCCq6bsINxKeSMF++klK5mFgTHvPU7/SWKE
CXVT9wYggH4qqYOYwW7jbg2cd34BZAos9lyiN2fnD/fLu3E/4PxquYm+yFlZaoocqRcyGncE/30Q
DbHkg37sn5LpC3crhPGjMYrAEJbcX8xX51B7N42ZHk+kKBIL62rRJtGZJxbm5fNjL6LZH+gIbftb
B6fRfs4bOcX/6TniXR+lN0Lwx4lQids7ZrJwSXqwlL7HYV02RF8zSHJNpBfHC0rL8ILl6fEMJE6r
IHaUM7jSchbORxC2E2CLwSST4HZpPwRIrT1e8nOXbGifobqx02bR0mJP35jo0zSTyLuicnhtVBo/
M1KU+RUgKFrh4SSgmOq0eJ7VewLUFNxJCZNsSLgIecW58cpkDXCLCOaMdNESdZqSyLBQqjDekeZn
f6AXOThOQ0cgnS6AwOeGHbIGMB9hEH+cxYzrnL/m8wPmGG9+UHq8Uep/xfAA5Bp7y8AmHD+YTm6g
/9/D+T42JVpFbCpz3r+fTHqoQro8sKgD/yztlDutiaMdkMwozfCOnqIt9ngKbs5OypNQ00M81t+A
3uUsgDjtPJZg9NiMHoUFQsuELHn3WTkXHPZAFQJd54BsEeVtH0hS8iADq0Axu7N4s49ZRCWDYrD/
P1Yh75ogFrQ8BbLqj0i6gBfEyqWM0/4SQUk+c7Ac7tk0YPqR4edPwNW5/O8GIiEbiXfcBhiVZbDx
Q5m8xH6WABV+TaeL/6jHUhXYwf6QQ4WY8oEY16+TmFZwQpRACHgIRZCJvxjjdv8iu8ieab/OjmRw
1Y+RQyj6IHUsr64Ab8+/avwADOBOj7hjYmND2Lbu2m6nGromVT36wZgpKO69bjyhIYf9RuvEBvuy
rIs2ADqu6z4MaQvyCCbuCbetsxn56i7wGRTAnf/lEKHFZgmr6M5jPK9Bxqp+7wSSbVr86eMwC0Sk
kR7ugAxXNbO3P2owwoM4Fsud7kaJ3ZaPrQ+b6S+dua9iR41SXA1HTTAcMl6BRBC6phKXr6XPXDMl
r13Z+7/33EKC242SI5U9YRVedvmRuAMtvw3zG+olwZqk0Ehysk5WopLayOzaKOIigRcqjOutiuUv
56fpiNKatxrNMj1hpyMNiyI3NCKVqXsk58kfGUzGU1YsEnIEzlh90n+lsiFVlWdjcb8J01RnT4qU
RMB7nc0/yLQmxpWaI0+fjXJx/3cUmL+dmPlY9UTZBKV0gr+K9jOCUW5WpI1/493MEHNI5xP5b3/B
tqWPwbN+2A+akytGTXjMY8bMFI3uuGTmRj/ugonWfgc4rbSxNaWLikajbrh+FIwr9CQkRhfNQpzD
LR4ycPBEpvCWI0o7AGMeKBC6r/Gpp6Bi+FO5nhZ9ADmR8+XLeaAFXMMeOIpVhtjcYI1Kequc2GkF
YdGYB51bxzJehpbK/MtyBjFnCSJBPmOJUz/vHeUaaIT9hHg9BXvdGokJySywuanOMnHgUtmMJ1tr
q9k4ldAGtBrCsKPcVkLHLBgepJq5F11ucgrl4C1HE1t/2PExkOkWT73SDPt7EaNPZ0KpDJiigBth
GqZpqX/x1g8q2WgIxdc0Gx6sF/NUVOF/eMMnd4g0yZzqioN/xQ+MXt3wsPPJxqITeCQuibgBHVGI
6NnqLm9D9bFZmDkP1BkkCrZCLc0ZJnPVwJpTSpYekksMKQXvU0omX2kU7ECbh0DQmi6X9v0O2vMI
pkX6Ij635HwifYvvk6KzA+T4F4XKoWMAz6/wK7IEoFSOv8lRyE5c+9SVtPiCww3JvOty3S+NHRr2
WiFYkBp7TZgvLBvIQecjEr0GuHh4Zq53Z9JgQfUD+jR5RPXOr08vn/G9twK3Qyq4mr5GkFIbrJrF
jVumhBlMUgfEj1LCn0OT8+0MNty8v2sDhE/Kmn3b7UtID876WTYgTXECb4PJ/7Xk5uMqFPgPKhzl
jmzQRuW0cCyZF00mylsUH3RzTh777uwCjbBQWntUnpjxldG3/SZQCE4GhwNLTlCJXvupIDtzKrS6
rSuhzEnl4+ZWrGOsEPrfSqn9j76XxbZGdmU/EXLslbSYm9Xmf18LhKAxauBarRkidh7ZsKywIOJ5
EGmn+IPxjiHiAeC1/j0zhqoS6TQcioo8cxlnMKzCcqFBXbQMUm/WK2VGTS2VrL6oUyRlfUxwBaB3
w9zH0gk1w3qs9WFWlsiy+5QytH7myXM2N+pTMyLzvuduQdJhkLS9yJL9Dy5bMasg3ITf9r4nb6QK
97IZFg5m279XTCmPSZx4HKSezXRf1he5KAjZxO/BeiDfCZVBAdjVmCeNkB/3AWgDudDN68a5q53H
RVeNgDlkI8OdLuAX/+cpl/l6MTPF+iJWb2YzuyAqTv9brT2Vmb80307/z0SMZLt+rtzJ/yDUvtWa
zJLL6fYhlv3zYDkGsrBTQQDwvLitof8prKO6zYmXdfGhb+qQm75mgoaFK18WRDkYE6TTCgtHJEf2
beyRs2CqwbGDmk6McqAa+7tc+pW5ArRRIpcHntdgw1Sjj2UO/TJhEx+xomElCHw7Bbf9mD3eNJbJ
GCe06a0NsbzWdxDKmSH0oEM+tYvhs+5hbM285mokLpiSMdYeOAii2znBsS//eoC7jipSHBm3nmD/
fdblpOIvGsaAa80Gmt3aUQtmxEnSjcMpLnyDl1ihep+nQnTZ7pMw9AL1gooOL9yYxvK5jtjh42hw
tIgEBZOLSrrkv7XXOHEJ5Nk9N57x28mlvoGHyQ6D7pLzJsE4lramIHNfnF8AUaUbL8bvxpIDNlAc
RyUrkpLDeKSsjbzTfdd7W5wF2ErXHFZIQosnq7MEaj9Vf/75NEK2XJDChrfk6QPePnXoLeNLvaso
kuQM5SgqJABqSc4NDHgNztEsylP8LydoyqDKlKVmksl4avfD1SJ/BfZC52nbrI8Llv2Ojyc7gDSt
XpAymtG/PvC21oajmsmYbcGIadNsub/o693yRCYrd3vj5/8fc16MLQuR2mmOfCo04c62ZubPglDn
lU5pQ02uZ13ljY34bZroiKicgtlUu07LVHNSdhDKCMIx/Wqm0Kw6nwA+FHSUNdmtS4WnCpjrs14M
GDoQNs8CMPSTHCPelJkIMsf0B0IyHU4ozhOE7fe2cWRA3rZDb0/ixq8kgP0tU9lpTZBlmOcjSrxm
T6OcUdaExVy912wrnzRKguBzEsoM621V47saeyae7cNH/jhfR6EFUFwYUl749eR8DIGoWIS0qX+s
QpKWZ8kOAv5+LmrJA91xzzshxLDrIoETn5RQ/rKDW5cqdywtKiEMr1jk1z076x08ieeZAMkvtruR
hzcLg6IkIq+Gi7xSqHpZJO4Kg0nFP9Ct6wCzr5Pbs9Mm4TYTrHP0+I3t3N8uohWWqfDJWgy6Pfb7
s5jrm/gExm0SbeuOcC0p3PLT5jSKilM7j1QX53WeHDyTK6aBazOiVGyE16v2y23mN5coInHnfmsH
LU7x+n4dcVyzbRY2fOm6W6oKs9fxav339i4is8FsCCKDROAhYaJzuiYw+79QEsKdb56O/8bk7dbH
13lBdmrRp4OyEuILIPEt7cKK97tx0JzbxRn6tMrvKN6dpsVSJM8xBgIM8AwxLGUfXTFv1eabDyXO
ECW25MZXxhufSsD/obncqtoUCX/KtueNX7ztu/HvPoMR9bSrTv0aIXck/wng+PrvTeYNWrvNVGeH
zR8La/kp1WFWl22i8h28KDS3MyvmO1B8xSNrfqzBlghOtjXdiK70JCiXI2pQ4x6YBfjAjvJ936+n
PZgaW36KSUdS9TKZmrThO7GMbJOVWz60gYE0zMl8BtHoOIW5gAAhskPq5P3jd+rBUeO+tmctwZx3
8cGhM7SR+nVwlFhlVvLgmhrqw2rTaEyMrl16SLZI7t66I2H6srah94dQSbtmjM+yh4SbSBkRPk1W
vjPzgnAzJxjE+aUsQcEeNgijO4+6WOC6ucoxLUGxOYeMb2OjoJd+2exgWGaBkch9lQHCce4xotmc
BUzFm9dSn9p6xj+k5PVaqpSxVP4n836TBPUYChYfQAF9mvGQblhajuXBkaRm7WCQjTVz9FW4Dqw9
gSaf76PO28RpnVoXsfXzJEmnWXM23ymREk92FbHNqlLTJ29RAu5MxfwYMnsRxcdsvApgBIGioQY3
MEklGN+LvvyA4FIhfh3JcIASZo4GH07Vak5irdCiusYZBEJxMxD+9JCUn+DNdNJk/Lsd2EQWtY+L
uydXK+m24igMYI8rPaonPyvCyVDNL/qMMkDNsr+Eu2BTgMNu3cIomYpJ3Gtpha/NAmxU29vRiyHL
OQiW0dDcVgDt7jBJZaf6ZjuwoAUpb03+UVwHoZguCGJ0XTR7eR503Tds6FTyNh9CZP2EMmbnONc1
T5duxYNrSCW6Dck/g1D2y1wmkVonZtwV2y6wb4HvhIq8gt4gTrW3mX5H+m/pAyHesSdFNw79YZUJ
HH21Vcml7Q9ZmJ6pPS/8Bpw207Ody1xfZCF7nMYT9QmzRdGBnVrFEuq1EYwCDwgh6ZAoWsaPRQfZ
OQu+XD2BEpjjkYeP+kIPAScD9IK78Tm3EL2XIIm3WSkZD8zdMNw41+AsIc+zCrXexWmOzaHuuLrO
NDkcwTFun/ZgZfvi1RNMqqtikuEWYVYgqZgptyi0KwA3BJr/y4MRl1aZbgk7rA4KyhbyxfBtlNs1
gXb9MG+22JqjqexD8SDK6cCPXVfveD4qyJoM2YKRGeDa8S3IAOCyatYcOhRlSEp1aXnjDmfhddy1
irAFvJf+CfdH/8hG9+5kUM1e9sawnMR6uNF0eTm+73NB+pW+IyBXaXOcl0oO8S60WtHCUmL24iZi
t1p10HUrktnO9X49h1N1JEE2p7OKPwfNGrLkCYXB/HRiPCYCRS7i+cIbkENuAXSXnqHZ3jquDpcv
XSg/jI+8pNrFLeglpmO/U1iG8QUwjpq4QmsrRcYtlVKZhXWo3l1OpiDhlQ9HSMAwtqocm12D7jsU
lLtpTFCpW+ICGndt+I4RNJMct/263c8RbQiAfNvz8wPrcBluiA6H5A8Yh8JfhIgm11BGv0Ta0U1s
T023zQa1/iMSNrepsdffg/OkpHdj5667AZXdD8p0iA9vHnmmy79/BHEkMr4BFSGu4gq8hjqyFlMG
aNomnO5DgJ7tSblSeyrwrela/F2Z2RwcBt7nkK7+1NrtUi8pa04ExnJ1IKLzDr+MM+ZiI9dvR7Ql
fQ7E2hSNL2Xlny96erKcF4I8D1xQ5DX5korwJK75lrayaZbKYFmvWpM7ZgvNJEaqUz3h6vd8GHaf
JbuyaFcSMwMR6tsU2X7ze0Mj6EY0JwbaHWZjaS+Dn6nHMgUc1sgo1CVxPdprtA6J0MErFUITRdEK
7qyt+YrvbfY45Rs8UKNApJ1TXf7DXPBfF8Wmec+7RjIUXdil2gBQxtfU3WC9WRy1SBfOrkuCH7jr
nOSWKK6L5CRXTQPvcJ1aTW+obFGF91RsIpFV4TmGiFf0WMvSXtGEOgWUWpYTOHn9Qd/g9tGDQ7fI
mjRJPbdswXEAKNvml0ojkvEjaQ4qxNVOvUAtzgmR0Fur5rO2mpwWF3h1o6CeXJBRT33yJzQlp8E9
4M4CRRpKloH54JtA2pmL2e9C7Df7GGP465LR4xJJBVoKbpWIIKuz/bDpzidJIQsHHRfAnLcqo6vH
oync6lBKN1Inp/A/ZyD8U9nt4OQtA7H5buuKdF2WC+C3E6zyTNcrSbVkkHMCImSkNWnUn4sQfDAe
PZwz6biPEOMUw+YcIRiK5/8jvvICzxXK2I8kULc4fCZcs/YPG2bghHnYOeB7VgZIOm0ENg/i3ZuP
y30S6HBrvuQjzi+JivzYblB0VGh1seYxIqs6sOpT2RfMf/VP8Sum3EEEeCy4pNbpQwmNJTkvEFL7
NqM3WxJ0Qfh2JpK70T1eUDKSBHURD/027ndOolmRbWFB2xIkZApHlnl8ECRWtxcycF1mq9KCddl2
Z9JN3tnvybLq8QFs+3dAbfWDI+zY43LPhYSTpoddZL2i4M13YW31NFalPhcKsgTPLZwtW+b/+/SU
m4lqKmuf7OXN3KGesBN4XP4qF8pDW7pXh7G+tXFR3wJ/GWFGgfbkswTTfa6Iclkiamuw6YO+cItt
bczfRiyb8TKkemOj0zMixViFF9WjmqOf7B2kinFKaIsaGFYOQd1BPKkuec3ULykxQtM54YdMIKOr
qkA4y1B8dhZPw1iLL26pHDRGsTm9tJTzPiI63IBWVrziHbqs/HlzwEmaYsXL4YUgPGlPHUGOtJQu
KVsVV2Y+hfeeS5fc/vmHCYaO7lXl7NQG9wLYCHm2NdXAzeQtv3/IYyRJT7xZMUKx6gotupbWHkEM
ZdBMkNVM12Kqh3JBJa2eb8hmxy1MbMgqeQbULaGgzEju37p/ppiBdt/7MtmAPUU4nqGmwwAqkSTA
1NmhUGaat0+FsEJRknmUzdFmJPK8dUA5l6pKcBaiiqQiiztkNCTOUf7sNNr+agkdJj0ApOGu6w1Z
eADflpHhR4wvxRGY0ZMPUvdbMk7p4N4/5nb/9NBAybTvPpOFvRSTe3rmDpaNwbECgd46CW1x+dAe
wFIsWcEUmtFeQG7Vf+pO72ROmUYiW+cTURO8ejMRl/R2PBqfvojks/iTAwJK3SlCRUK0GJumGhKq
4hrKmmKaZUDt78OVnZaTT8tPZWnjAhBizcrTT5oQCqWyFdJlC3jvY3ZGYDEoIG7XNzOinCqpvd9J
CEnfWx070/5SJYsp0UrWptna+3CfHxeFnjOIPUXiIYMsBlWh7TDkrbm5qeKqrsUWFDUGno1wFMNY
Hf1RUi7l/GsO7PGeIM6Pou6bL/SrXx1n4vzghLhI+XsSiQhcLSPBprWPIxVHBmRUAhE1c9vSF+zO
4TtGpVe4kHJVn+SMhIAS0GWBCJTaO9BAODrdpDdozSPF/J28AiKlW+w0twCf1pDPzLtU+G8LPnGR
IarYEo5Z7fESSFS8xfkqI+NRE5GOR7j0Jct1BPwTNs96HYratAeK5fEIAzsd1ls8TPtDBPyOLqwp
DKjOAKZIhnFcZRV4Ip71IPruDnLYdPczQqZCvQ8qVYvzEnDxx4s//1quPAv0IGzacQHc/lvrvFBp
TkuQaxyBfdtN1ZVRAIWHXayDKAw8wqOnnLhf9zvdO/SF5rI1OllGB95Llei/1CmJweImxszs6NE+
+DI5DvvhAajLuL3WWWQkdOSa4QkzP6omWi1QuFqzMFPwKz1J4eFlrAaLO5EccqP9HJDdgyUdMJTV
kp/XhRiT0TWRol7HT0dnYOGWQbbYWY6ITKwvICpNs7xtGJQnRv3skGUm9Rf+Pw4z5RZ98nonyWHV
zCaQH3FvezdmyGk/2EzvZpgbYR77ahOtwAtikWTAUmOet6VcLg8ZrrYBjWZYEzmTFu+464Tyj50p
JY4018wZ1SaXYLCZEB6wO45gSlQVX0Ry2/kQgPqfkxL3Ga8AubVdikhXRfa0D+C/F8gm+EvSHTis
h9rpuS3RdFSwdu6OeAOdfm5j7LEM4NbxbaViPv0NqQtUwUu99XadqKXh1RVaAuCPrfjZ2TReC1z4
ingSwq3ofQ9tqA2n5qf5+nJu0fjsteBX6J7kQXw4a3Ar4DUfJ0UytqjwfxjDg3jqeU0a7fMzQthV
OdLuqFRBMxnLdLEekyUHAkAnOedqmRd0mB4nCytiH5ZvK8cWK4zwPbqpUPP3zmvOYgy9Wf15ohQi
KGSQq81D6ClibXDnKuHbqDUH7IQtC6f4KQAJvbhru/SKhta5QoH8XrFqAOEFHInIN5A/Kqr6fr3l
84Q5aiYzQhD1fdLsQvEzU0HWk5kcxgBNDll3wXPaHrDEtTv1/iPu7SZNPsppxP0SNFaIUwi8bfWq
gl9Zrg+UeRRpv93CyM1M+j07qS20vPbMzl4g8HDzxS7lMNEzD0dsq45SYYNX+AQYM3VoilVtOxF4
/TGrG8fxgW5oe4I+5Fe10qbFifMrQOH2Ao89VgB9HUtyP35llWK7iiyZhYvf2ywUIIYGHqIx+7H1
LJYI5JSH0FAomTWJzXToVN/HeHRwoiaYyMCF783VEYHvZcIQwinvZY3V77bWIJ4bsXorcWIh90b3
qgiTZ3PpXke5c23IS7qRGePhsJnVf0RmzKko+HflyRmCUNGMNMAskMQh6xM0pe2Vm4oe0g18MxUa
BXSKfo/NtgUzqo+XlmSXVLJFUGv+tugY81SsYgRlx9bKM+HJAhyE5xubsAlNsV+sD45cnxiKj63J
NUPTMl7DDDdt1lL+VQaI2xYOlApGWHua9uF8zUhcpfN7ASJDTC/h6+EMqR1al9ZbhYVflcCU88bC
McFejLb+YpxSfQtfw6qq7KmN7go7Sn1IrPXoIGtgrQCTvc5U8TmzXHwBKBPX7oNdG58VvXJh019+
SjRdV+3mYGsY6EgGG5+iqGpBp4Q+V/9M1DqqSrANnDIv9GXUsbBT40TPGboQp/7nlF4speoygU0L
Y16OEkHIo0wjBzOoToS65WmgHQV3vHGDxottRyDd+EWD4WQ1+aBZ18iOsD1mGgNvHaMv6BN1rbKu
oOrKqomfaz7TPvjAZxnQ4NfVnVPQIMcajQ6WFq8qSE0ysLD4M5bvo6DoesRGF+9XZVu+Ay2XwpBi
R4H5iRkXMy25Oh4MOtAwl6vKJ5XGcap7V/u2gTq7XWXXW5Qt2UgkISqc17pa7CFcM84YHdYWBAYJ
y1GvFpZltlHwIbvw/PQziC9JDdWhPCfrQIdDfDIMtsqENa34AX9UFL40wi1RtglL30941GuMB6s2
8AbkpEGDLr0VDJ/6dSnCNyS0Qx4APePN/fCYkJbhkBwuzCZNrz8O1izJ4AqMQrJg3MoqDmvN2DMN
tu/fbAOYNItuQTOInWf52s7fSNoh8DE8SE505+J6htgo8q3RidGiJeSte0FXnJoZxCiOnpRdGeIf
Eb8C2w9xKyz24OMtVkl0HYGpRHK09hxNy7MlPZWfLBX+5DuloDSjYhVUMviw1hNBNHMulL00CRDa
WNTxG50scHKzJHcCCAd4nRrb+2WNwSgfeM+UxWEQsgCunSCTj4pUecpRzL/DM27hM7Rt6IhHuCg0
/8uNCMNkuuC9mfd3IqzpfAlQB4xgjKnTtJ7CphkiIEXRPRHoI4JOQQlUf3Ea1CkjPL59s1eqILSj
JSZr2PBi2mJ3375X2MgCRBuBKxSp5Jp7nD5vMnAHF09aYfh7Tj+RdIAEWT+PrS9CP8Nutw8f7Jqe
xgRt6bnVnndITu2b2FyzGsfkCAnNy1fcHIMAfISvnlCXsoXr1yC4RCnlp8N67UXIi5/YB+F/I/dl
E9pd/YgV9D2CSBxpCMScV+Q3RhjmaynbHJR0Wv9LhFI2qREIqsSSqtfdAAyPwY5LohbyI/EOmfWE
cQEFDiLy2VbzI5VmQzl+aWrJJunBp4gsrysnp9NtdMY27HeEhfYBVj6A3z3M6+EreOi5UruauRgq
1MpiHuU2tOgbp4m+mgTFpw/DKxeB9ZLnBsEQ72BcYXFrDbv1cKV8syuJwy7gcM9WkT3yOz52iAJB
8+G4zMcxoV1Nt012cf6JgsNSbBOoEpFs/oQ6IlgJpStOColW1r1jyXH+J/tEu7QsbUixCjz22oKe
DZrulAGRPcMkVwBCl7EMfo5B1m3DERRE9GPZ3JzrJkQJDN0KqMR8Ya68ru93gYIZrcSQsbAM1L1N
FFHuOkQuM3vtThMG6BJaKTI4so92YM0/nyyErhi2jgaYASuger1iF5YUkvgTb8/tqgwhTrXlAfjy
bwNk+yiknmNYGsQsxwpbseh5TbCwaZ37H02uk6Moh/cUVmq08cva3fXwiVdb4QTuT8V5R/ooXSI7
zl3Fr56WLLVR0URRtulvIbs42+tNMT1qLS39on4cnJBJim6llugTpc1NJf/rLE0W9ShsZ7Trd9Fr
rWptZtzzxsFJlJCGxWdNW5UAVg4m+JSIQDny5VaWkfOOPhiVg6LK+5AXdhT8afxB9QOzO/rVuKQv
D6p+02Xtp4cAXP543ci7C/OMu3zXae+Fzc+he+kJjJkpgYxyUbkk1SqrBm4HkP1uv8/tU2VkY+XP
OBqxYLX5B7KuJdqHPu4DcFzFfT2eKcey+tz2ssYFtGy+WMW/JllxGVxe04wflWy7uHvdl791Veau
GHkDwihSA/oVCVPplMUpjSBN/OfQ0ERsLSuLxRzipGfm+22SLSALyeib8AuKzzJPm8Ga1G/030sx
vy+E685XO5vDdGBreWVXDtXP9UAptSNsQW3HQZOCvedejcG2dFWoG/8KCzpLW9JPggwBhrHN2L6P
yQBRB5YPnuiNYhIcAyonXOpEn5mjyEx0ITyqvMDCTD/FmDkAj9YW3AZyB6qhE1Ck/Zwmvhku5Olx
ZVvrPU7hh9bnNdZoiXtjecnWNhqryrN+DiKgCCEUb773j/DkbVwitPm/GLDF4ru1eN0RmIMnFN87
/TzSuswJqzSOWTCEwmOixn6b7bYFGaTiz8qW5rvn8Ez0+hpy5hm2UBMs2wGhxdQByti4rabRdFLb
6r7waRPSr2alyOTXtKjb21ECwzk2hwYEsTqninfxBZz6101T4Y/h6ANctApTb8DLRHReN29pJLXb
JHf9WQBvzQwn+9V/3YAZe2YrE+STq4NCxzlYIFeRQHyFsHam4bDfzo29QUmhezSLNAXwDTmSOY2E
uH34cCZwndp5j0iqb9Ko6gfrAo6zTey/n5GErgNZ8cVcjBN/aWPmY4mcJ0na44zcVyQy39+0cBXG
P4suppPk59u0hSRU/pJYCkTwpWO3GTPlDUKsLXvwn000Ikm9J0z38HuND1TuqiRax1srXCH7IJ0Y
UFIBV477vH/2zeIYdSr+K+Hv0obQuZ/N+wzRXp6wvTCCQTfzejEiNu6S3B4M+ljD/Kopi3R46Wwz
9BJtHsX9FFyYmyJbcuJxs6A36FnuSqZYyjkVr3VpUuPyC37NinM5kAqonZzOva67ZPIq1si4uKrW
iej9ybpR+Ucub2nOOD5N2ZALWQCx4S1yps05VhmwpvRvxlOQKfzCEgOLXe5ld/mDN0Uqw1Q6JAuz
Fm9YT30CluzLbWCC30LmtFmcaPVadt6mA2uk9tfNk1AQFechcHvV8R6/Fut7l9g8a65XhEOOj4KC
cQptmWskPDUAJ4OuJV+lq05pdNjGAVaNf342y4YxFLmNhNfeztYAjAef5Y8WgKfvLBALyjHWKtgq
kC07bD7l4vHv+s4exZi6PWff2RKQvVKrVx936/nbjCR9iEEX3boquKly8W8cL2M3O4bd9pbB5sZq
LnyJQsCi7Eth6g7uC9yn2lc4/1fa/+tV4nkwlNeRAF45Cw4tv4XC5Ue0WH4GQByZc5q7zgMUZFC2
6lmkuNhbbZ3+z4skrUXiwoYtWquZVhNxefFPc9x8gsSLDljJqXjaLcmYFa+ZjSF90sl40p7Goy6J
nxq+sPgibdmdca3O4BghfAZga1l3HlfijhqBanDyuIxzn1l8x7qre9PaSdw3MVKyJJ8LqbwmpTyD
LjZXVpTrXVBWs5ZOtHnE4XcEeajrHatDBISZWp3k8HreVK8TeCcjWxryWrNSTyJ9LpUBlkO7OIAC
FSOZ9VXxYXZ8XFKzqXB1NG0tdOKpsJmmjEzQGk8i8F5VoUiZYqKQupT8rFy520/IRE1FKsmhM0gU
BSEMGT6NHFscp/cQUrRFtcFZGRsrs8EzpH0h6E7zW+Sm0y5wxWtUQOt88dNAU/NNYM2KrJulEI92
7PohGVAyMfNMwyaLmlYcGiUh1HddberV5UKwqQEjeZA0p/AOcFYj6HnKH6oleRW0If10+A3R36zS
ePffWz7HOkfuetnEfRPpFYADP4pTlKbpuycAljarAgEkbWLkmdsKFzMthW/Y3GhYhsahhp+gx4ll
or1PIZNDi3RHJN/BpHl+hv7rpNxSHiAgO7zRVn0jMb1EjKgk1sNOfLTna9U9pBHrHyfoKWQCNpEH
pbkFOnQi8IAdzyzQ3MO0zJHIxxlJIaeR+xhl2gp7iUVMn958EZRhpaP7+Xvb1Y5Lke+e8xb5fj+o
KcUqu8Z1rn+qx60cA3MXiJtnQ00X5Tl+UqJYoqObD4ZGvbFVB/8OtCiBf6EoHYNjtEgaHuwo+OAA
WlH8br5GhtUY5D7WXL+W8JZKJVl2Bbm2CCH/RdT6lIpY2AT5cJVMOLHorfCOL0F+9WA+axHYGBHG
zmEbESJayxutuR7oUpcRMllSoTIPwMBNZcEbnWrudpnHYf7Aj64bF5LeexTk2hjR7Xja0OV8b5Vf
NFIEb8W6O8ypUH0QbVseKNl0PrbfjafN9F/Aa1SEK+jgDJKOucLDYWap9kFTDY8UaP+oEXcMfSOa
AurzwA9Kv7McRQeN3VyK8zZYRaiqIDrOrY4iZtuCm/2wC+vdp+uGrnlbf9dW9VUPF+Kb9nEQ1GHF
aeRB+ff/j8bFm3V8yV0bZ4BmkTTTcd1scB5tuPF4ycavdRGUZ33ebVX+ByDtNORrqWgpLNEepTmw
mLlpB3FCQ2BJuxaGMCQXALnAUxzJdr21qB0lb5ffLRLNQR1rKu4UY/6kn4PGIvAi8eyEU58zknDk
wJUWKnPZL9t5DDjwSkE2xpWmuAqD2RmZ1P/RDX2AZGTgwOPx2epbODvSS+rpUmoMuEm1clJZWFog
aon3fUilsIwvlceAsrfFtaECozZKR7TEVV3/thylOlKH93TsI1biagWHsxeZssJ8/ck2lydy+DvD
hsi/UVdZoZE/uIYZjLsckZWT5UZ0MH1rnhSJSDxryBexwg9j8Cuqp9YQ2mMCmHiW9n5dZoG40z0B
GBFFmxgo2xDP6mCypLPIHEuesxvO8kCL6WlDt00AhqNNSmZLX7R6Iyx56zzDu0Tn1iIre1M7j/ZP
Nay2Ru7jTuAN+rmuda4QRDrSPwtXgih+XXMcdLr0agAnZ1zXyTXBBkBIWcNhc9/G8knCW42ImyI6
qn0QDobLjf7xgoKTzm4epI/kqSvpynZwIy0TNCeVP+rDHgoCHIc9/fNn4dWhIC2+7KdYts7QyM1A
foQkYEPR5/raBXWGBcQzeLX4O2jrc2gt0Ql4dEImMgnPKhP2rNjrnjpvr0lyb4XxjiLeHbrU9dKA
VxAxT9+bo+PKVXbfE1cakoP1lli1FV7U3ZhSCDg+W+N0pTkgA12Ml7Gd9JruO+K4dHJwDLBNXIlH
AR2wOkIUd8qXfRdmoKe+nh7uGx1xdzvk1QUc7GlfqhN+ckPX0D6qKa//4qraniM9pm7T0TMja1E8
540ADRtDO+63WkajkbDrm5VB2Z1Yx7weuEIlBXxuowBfR//hlkGfoubi5OTmSZP61U9TyJQHiZib
a4rBBr0Y92oolMV0GF7gM9hreY64a7iTtcqx52D1CYlMsqvqGBjTGtBThA7otV2RUHJI+S0w87Mt
Jt+qYUKDGFuAZhFKh4Eflws/4DuJhqlZrJik8w7zVOp8uBt8h3Zr3hjz+dyIDvtjP99B7lPm/Maw
gb3uyDGdSow/460ZsiZCeFg62TXsQk/DvRTjmrtUix0jEZ7KvB1EUz7YEvmtvAO8Q8DnjlPdxgW6
aWhuy55fgNNZ9dYIQ+siw6WZrGKykjwWAqvUi6Iwtdx5WKqrnyLGV+etrtKvFsL8tJRhIpIzsARQ
zz5anCr4xBA4KwTxCOIevZ4R/b+IhsUUdFIdzsZEiOQg6EY5LUARuvI3Q3NQst2u6eB8aoEl6AbA
Um2etyCoBr1r5H9ns6sKDFD9iQ0aKK0pSQW4it2KTdZBbzbMzWm3nv9CP+LNL+gdGy2iCFqsaDKi
AdFX+7jWjWw/N5pHHOdK19iZh+TV5c5fXd/pV/cjeVOujbtNJQlnaPL3YFgOtUMbHD/lXRGxbk/c
gm+QYT9nyRg4j9DZUz1UvVd+leJqpuaov+J8CBo4tm7ZegRni8Qq0EInYYAVUjmfSFc6m4wGmZ7X
KLH1nLDzKnyzAEbacybA1NiuG5yWWgvYQYtxQzIKj9Ee3gLo0/44jsxhToSWBFmQ3SIyMV55nHxc
9E/j138rObglzNMxjuQ+ppg3RgfQN/f98NzkMOthvD+xH8sQinp2/U7ZhVhWoB+lSUhe1Rv/TH6l
/CoGbuIgbKOPBm9nFcRcJ0UTCI2gsNagm8qiJbAD4mxZCFa9AJi6kgaSyZrKHGU5Bh0b29zVg8Yl
yn5PKesRpbXZlOtE0+Rx1sxiBdWwx+ZDPK+rKupySAjW3F4cDkdMhp6wMLtwdM0EPfhjG2vOaZQq
kGAQ+yXjGuyVQ16sgYrQYsqTfyEzzu4E7nr2fezTjss9hu8hm4nnNSksUq2RWMuLeZf7VbPFUMk3
W6jdnNltLvehiyqzNJm5WnfUBk6veuRSifdO6c13OpDUeayitPVIZgstd+BkncHV8dWOXS0yVI4t
gR2+ZtxlxJW2uYhvPSdL752cilAL/lwcR/DLlD+FHawylUQCmTMVPl9lZpd0OQe1YErSrkjIhegs
c16VDC5jwwntj6PhQQ0RipS+80JfIBmDeSf2KmYb2HD8qpQnTnb2IxZ9eX5BZztjX43GTnYUhRNc
8yy3oXR3ZpQW6itOihJl4sNtQ6LOtUG7cou4UWPb4YVhHwyRyBRS3ri66mxhLtOOre3rVjIqEYl+
UhDDscCQDHbSlpmfbP2FIBjsLbg1+oN/4y5+dvAjl4CbAzCpgyWzc7MWzrcCvo4iWG/naNhdANj+
I6v4QtZDy4EiUiiSugzibxSWo7P7LzlJdG82uLeyabkwvNkB8eK+mUO+oMTA3NcGHMXVn2dhdg3E
eC+YYAPisGA2naRhoFauHZHWOaeNk8MnSg0gzfvmnya8NKL0m/YIY/QrCvrlw4BeiRU5kuP0Qa+M
AU/5cBHpbSXGonWLidJOr5rDLG0cVO63eyz4mLb4GDtudIw48G/m3+hxu6072Pd8SVMIe8qGUmi2
pJ48pwpxnFlTPsGHlfPU/ANbA1hB6K2C8k7NRcGkMRfmwX0GmXv27gYu8d2ERR2d7evHTgO1f/4z
AfyYn29EmNMssLqxMBdFrohlymPnyBnrHMy++QNw9tZNXN8tEZKjB6AY3dXNN4KkfU4OJB9g7Byr
EFojkDZvW0z+3GC4g6Fy185nzX/cF6+Psi9VD9OvsWHFU12lJdqiqFLbTD2FlR7p7NnYc9qZjPCI
vXA/DRe0S8mzPBl3ZwC5XrtD4eZBWiIzV9StUJybEPWuBCH+GCbdVspGjqi6nCbt3uWbQAiTFnD3
6v+uIkNixaNygiSq0KL2cMdocipNiiNm/hJwYUmz+TIMHwguDifzbwzO9VDxiWIUkit/1LQsH9QU
uXdckkHjAw8s2o+64l81Yar5KpKatwNHEqyYJqFxsReMPjbyMeCC16nRL1/kwAFVpjaMN9p4lmCr
kyCo118pfSvvCDwS+3sRNo3FhapnDGZgVmgnhjHu0fxH9yDshO0UIPuzbSGYVGMpuab09R8OVw88
wozBYEiyEqT7RPewnzsfV4EzDRBcFXFLJboR/FffxHUfSCNTRACdRarZ3BmrPxsezYwXvuUze1Q7
tIP/FdL2Xbr6Ste4pni+wmyN545VFHgbVVEZ035NNjrXiVNf4rdw827k73MBHQ502DVYX0Mo5p/I
Il/6+GdAB9U3Lh05j7MxrJfAenNGBeI4/joSUhqIMWB4cfz5gweiX6gULu/9SCp8kIwSR50Lr3Me
uh3FzoAODfVwTaaqTcvWICetg9ll91qNsmJI3bLvWUP5u7Qr6AKmcKEb/FrEQbT5m5Ro+uWk6nDU
OiolFLECivr1tWoRQ5Ezu+fXUZha0wpACkRCG3hRgOwjZXaP9/76y3AgnClUi143Jh2TN1kLfc79
gD73ip9qz0LYpdoRHLlpe7mm0qzj6oBBtPUovRU+J0EP8gSnt9cT5uHbTKnhdaA9IGqGhqBiYtm0
jep6Pr2mPSRg2k0v2jGjS3vPYs2xK6lvioyaMFCM1gdLcrliRGlrtBpr8fylSgnuCFHwtN5rA7Fm
obLyCwDDBJVnjJIZBEAk3jkPzDX632GP6tADIUIvEDC4aaIx9oQHxXpbNYMzsGKlNv7Gelt+fLIC
MsnngA+AivpNheBry/OqFlyuezEm7BWsy7Nwdbw3m0tSTGn6UzBMlH0daYrqNF5xxrnABl2LC4Cy
vO3yPH0EsTBr0xDZq67thLOKrZz1mSCHTy+eabh5fIXtXBZ3ftB+S64gjDZDfAKrHq2sns8rVGTc
Q1m0imkEmzXi6dXEO+3VoKiraYnYsGBxVu3R7GXai3Gd6c2+KzBPYwtCdHGOWWTFRpk2cJknAz5R
dnBQK8Gxz4xUTt71ATnnNAd2obGCnmcajTTgSnWyVqRT8BM2HEL/j9t4SFVLaPt6vEEAZX1J1QXf
gpszkS7ySdbFXy4RHNyuWOfnhMh1fo2MVejLnQ6fwlBSqE7h7xthwhfBBbFIEX1lp7IHSCpxQ1jk
ydbD4NkZIl0GSUiDt30zwPfnEUrvcdE70Dmai1vN3706OKl1by7IuZgLqnxwBhFS2Ug05wei/8BV
m3Z/6NBPxZT7DxOPlLxmIiQuqGX45tptgR2yp3ZsUCfaWtzLIzwq65DTF/EjbPk7RUPLmpV47jjY
EI0XMlVAC2WfIgjCN+qBG7mug03o15TMxM2VNrOSP1JB8hc9kfmujmU+NImdSKaoepbFcXqERWtX
eLpGtcQhNszaD7gJgT2hImzGLuAZwCl5z2Li8vAMUsMuIxz8i4EcDHFveS2atRKgFeDnkBQ9uAEO
8T0rt8b6grOuBOFvsG5anQFvixLvi4sDRexRUrLPhy39fRX8OH/EjpllklbWKrSq3W/yIoLI5e3C
JasWZKSpN2GugQynL1eJJt9rkNORs/SRdixRJ8/9einIkY+QyFd0VxISwXEHxXcm72EarpE5GHM9
jzrny889tiPzvWszOW1WomsJnpn+gj0Sbcbvy3ot3MljW1dPalCOrg+csFMB5EjWsTQuwPa/InMd
YztRF3xwXX5hCOUUGHLzubz+QYzpuKy9yItlvN8VM/usJm67xAKvAI3YyuhVh5XBw80YrVZ8HASR
D2imnojCdCLHJ4coCqIcdejkc/8sSd/hQqXXCFi9HuQYgC3IfhEYvMvc88GNaPBEskjM/sdiKI1N
rLZO6NgVhDr7/6aVgVCHB/JeufO6mI8AkkqjLCP8VZEZi3E7IH2j4PDqcMSby2Drz19/bP7LPf7T
2vt3yWQcmYIoY+j8SrIDN/mfItYwbyY3yS/bpBhoUXdyIEy4oZVc1OblZU9WxkS1+R5TO92j6Oye
FILPAt8mtp4Qnu5ElHjPvMecIFg8HA2Z1p827urK/YOjmh9+/N7j5X8XzRMxVK0hjv8DWl8Tp+Kj
V6U5x70LimKzr5oKN4Bw1Flf4QzpMeKSfcFCU3080Vb5nbrp+CuZA4OTttRrWw1ohu7PUxl3N39x
/TLVPtoQLQQy7YK+SukmWNM3wB4Rgo23T51JOOWlB5+/eqXDu87IjEdMXFcTb83C3xcVNy7V4mh7
2ihCwa3SAmFX09j/L0h4wYOCTRURqXqb6zSq1EGUhjh8iwQX8VRdf9UqvmwNppZKSSpJ+q/6yYuT
Y86TtqvclrO22kJIYPCEPkSzSc8L9rVcrZuXhsN+vfny3pC2k64uaX39wvRCnxKSJyKKpOyBPh1G
VuDycxr5vrOTxmPJpcASMumho+3LpwhayZlkBo5wA9YxJeVB9VZYFE62nmh/m+vke0d7R5AsXGvG
1htQPwd3CKtzp6YgBfWzMl+d7TAR3ZaHiKvicdNmg2di/GrBUlBbgZs8x0ZSoYYPOKEMojWh5+bl
DOi99VX7/t7D9H9L5s2d0PtNno0OBgD4ge4bBGejCxUUaTHt4gyxD7/M86/noV2iIms61n+armSt
dYKv+kFDHwMjYVUZyfE7PaDMPpClv9ht/Y3KW6EofZj2k57jGaDx8s/sBA4zu5k1WkhQfUef59va
wPqo1u0k41dmYSEsylbIx5A3X0iKZVtY8RFtfmZT/xVzDqWeiTLqPQDDreZH8sWoFV9SVvWtzkXf
MNgn8+mQJnvykYX1NUGLTeVFyrNnbSkMHauNxbaQHUL9/cW5DsZERZ9hPyEk29mOPnhEF3zTyScw
sCOlgyf5Ovr7d3Rr6Q0SbrSyuDD5AkoUdaoJ9CzEm2wAPQIwX9+wYToIMrxct2CheH05eqJv26px
zX8nGmqBq8+WSERDdbnNKLLuQz/WCvx7PBb8LDpzyFQnFwNFmuICrGauQHc+yKVGxpWirLJkYyI+
cjKOoeYKkiqPgiIeDEa1Zuz1xxIvOZLs3Mv1nHNw1bEgZ8oZA0Xu/E9dIdKzrhyrkC4KroKrm1d1
9kYFJzCraalSmowSuVJDvCT/DAdfdGkuB4BlzxuYlDM4w5Pos8awC8CGIlQcU44o4oJr2pyVpRml
0z/0+qioueL7sfoYOreKBLqzDemJXRq1G2cmYHhdyp30GyuOneFlUiGYvMUxuYY7Wnb8JnZg5LuP
drcBr/1b3wgLyB6vRLilLEekbi1/RVnblvDRSeZmKvS1ZJTQ93eF6rBCGthZxc9z9XcwhnFEPQ4b
zaY9i7cXVhSSAlWaGhSuX3ENM8kvbvVqG5LXXz2guewwoJoExXMp1VyFIDMhF5Kr4kHjUR88Y5++
1ffKhy7I6CcTZApNzW6sQ2KQXBx5nEQlD9ChuTTThH2oIbVAiSfMll9FY568+rZG2OZ794GUdLMB
W1DO8tZESfEThjUhSo1kziQ6WSFuca2+AzuoVR9D9j00s2te2W9ZifIrGEtkGyStBYSqkfeKWqtM
O3ex3LKsTG0VFQYgKdPP6Us8PiN8rF/HNVHBRiNCq7/1qxl/O8o+w+Ivkc6qRNim9W9W0KYt41PB
Jn3e9NpsfFbuR4Sy/hwUIhdKTOLfOAIIAi4t+v0mecM60ITsW38iMEM5JRXYGVpWE/v6g+0L1lTR
Frq+NH6BugoYxyPG9xU/4LiVB+EvilkCNb6bRIsKvRt6QSUMcsiC2Dv3Lx7VKRWDDgWieOq7zV4G
NgeliOC4RPBzm1F5CikxGGzVNFOzqdKsGZ4iNc3OMozOmZKUB2nrqOqM4tCie6/ESA/+eFTNj4Mk
r3wOAtn0+w1FXKMkBdLb7HBHMq3hGPy2xyuZPAi+KPw6rJKWPDxcv72MPzllHBGTmmlcrzeIbKGR
Hwc3428jmg1PhfMtK9vxILzkYUPlenB+ElWmsbpNbHEVngqEdZXU0cf4Q+uiWoCzvwN/c2IQtwSy
cTP6ztKYXIpLt7s8K/JGADI2QcGlyU9RihScOsxfcSzVdCA0hCvRks7jtjnmjU96z0pDabGI7vEA
2rXU8iACkByf1RyNPJNf4ZfI/OTWwaMtbsxS/tv3QALz2k3RpEuluqRmcipdPoj1hpeFMBJyT1bS
9MIPZeKPLLnY3ITOmQhF54T1Fz478UHN0RsP3OtJnp2ix4aK2SArz3b5i4TG0AmH2aYpu/x8bcNR
WhwHmtFc7rsol0Dqg6dbLWkY/lsZsc99VEhP1+cWgZ6QHXy/D6IwQwMmVFVGw9OAsIGZ6CrgsBBP
9RJ5Elqmm/CTTUmX8Xp9Q1e/4OgxZ+Q70AmU6bWNC9izGILDVdt7Tz3QKNU79jUlsGldr0STvYcQ
Czecpvi7uFtk6o4moYJcDchs5u512iNjJY+CfMQF48Ad+FqYZy2h1n947iY7JRRHX5a9aqLAhji6
t8BzMBj3977Vpzc09FOsnzFDpGKaJ1BeuPfcjMPGcPg5CT1wlZuJlrjaAPJU0ERU2osJ4XesdrZr
dQv7o+cItZjzpUAF+rJ2I43ZRO4KIrC6el/g7ok+IJja2kN4s/Nk/iUMjezKjgT6z2I50VXYB5cx
HHd9ZGAyzmhWtfQG6RjBKh6pOp2esbLoGyVJ15sYQBOP9UqGKcyjs9aIaGDnS+ECDXm+QFOjvIgK
fEhvPkgLQEcJ9pkAdC48vV1atb6nmVaf2r1DdBJ4va2CGV2CKgJjrxbYG8vf6+K4URM1trghMHK7
Tz2VPel7+QRdYqThUrFRbbODN0Bs8piNgfpnf/yrY9+QV0UU0PfC43qzO0Fm/71F4V/eT4jFbxn6
cywCdPHFHAACCK9fCi8bN1fLguDa1JVJYmPRSHibi8uWcZu43IHxa//A8+K6TTHjEqVpGUSs8Gag
BQA4QiaXIULZSVcSCN8LVT9z19FVsNyFW1jBtlD5+vcGoloWsmeaEUkeg/hejeUVkCRJIP594H81
YNZlS3/gqB7U9Dk/2yh/wnIwqkSvQWmBO1WD0TmDP1cbU0KzNsNRWUW8k422ELYOEtLy6kBcq3ZF
CrnE0YbeFCqgrShc8F2D4dLGJWv4oN7NJ7bRx799mL+8GFbwkdjS2H47kDpg0N3ITNibpRFcPf/s
pmSpdfhiLlfAxkiMSi/gN+vY82zUGVPWhys0xMBJA05rx7rh3IMJZ3V73w1HMUQK+AqsbekMHniK
D4DO6OhJVcMyzENuiHwwMwZDc1uoBZntU2JVB10zmJD/neKhzZ895PWZ2SFJw7/44gVQK0ouLlSq
0YQu6cE2akmdReVcoQGhyrkyopvz+6xpGLjCvBoYiqSQ77bHKyomivesJ6vB7H5miaA9DepqCzjF
8olT1ZUtE0GJeVopjWYTFF8+UNqLy/U3ZnopsRPvXeihQpJyFsAPG4eqDvIMu4hmB1zUUklznrgC
bJW1BeLET6/wawmdNR98vip/WG4bxR2Z6QUtZeSAcQkO6M7O5etLh0JZx+yP2zJ8RVyibe7SXYFo
SmSqi0SfjmVLgsgZ2FLIyculora4l1F488hJprNHxqmuJAKo6PV2d4oGxnkcog1FLMS2mm2MxKeG
Am3Gbz4o2w9eyCEFndoxGXaYAIlbTo7IJJeeR8136YRpRaulpZKfzcgYGtxjoFon4ugnt6yY58sy
Is0QKhp5I5MiVUwNWwR0CW9AO7HIHYk/cfYeZ2fHmc9yvurBHi54p1uy411GkbWnWLrVz+vRe6Fd
L6z2Rj45CUAJAVchKq9t/gIeFNMNOH2uuq2Voz0ZNQb7tOq2AO1DAoJizKU4j+HZEYwjSU6qzm5D
UigNRR5/nPM5AD28qobLRCqdbz3FtZcPzr/mQQknMFPZim+P13VYpuAEqY1857oNQzYaJr4N6/ce
d+BfcGndRA48i3bG7+YrghNIgUgEciPVRT8dled8iir+bJLGynLhaYtvdCwycHXbxxsvZ4I902JA
Pua6OOvPoB3CjFBX4aoeopKreoOhfITM8T4mx5S3FoNlq1uxlPlIpPDNYnyvt7uk27h7PffUFTqk
IDGOP1dMqfYWau8IRG48kD4nPnbLWCoI/FJcHeM7/nHMOMwDuePE4xV/HrjI32YeKUT31omVD/Ra
N2lu2laswcWLhPFUV+p6jk7s6NkYHj5R2W7Pqc4M0Iq2RgZ2yOMLFGYd5+qhoSI1q/57MJMBuvuu
WtKWP/aCStRBqUzSwiGA/fBB1HMrzS3svp416UHhQYEFwF0u/Hz/vtSd7vQM+MYrOIOCpggqR65p
eWETT250MDfhclaq6RgPVPTeFfFo1MTI1S9/I+/21UHdLIgLOKiGk+UO8PYS9QvtKDwbSveMrnHg
di6x+QPbM1d81J9HxpStJWw0C4HupEZbQFBmK0r7JprQPiGGBZH24HSWV9gBGm2kOay14wkNCgcL
dbB+98b4utjsXOhO7j+Dx/krx0w/bohOvYXlOvin1NuivA8NyDlwONP17PqhWbZegAbJwALgTuOa
Gk5nybw7FGYfmKHZIPEX6p0gWjnjwnp4q8VXMbYjQom8sjOy3tgisRDHNyKlx7oX+IWSrLY3wRfl
1+FHkl7u8ZvA4VjFT2PHpLSWi1DPkXR6BCQ/IRdi70h9ryy/m24Th/3MeLi62w+FgiFmEoPsHIJD
+inBteo+R2ledDrqcdl6yq720LMixog4BYqnvIrUP0CGDfRLqTKiPwBmEel7UkpUqvX7apf7E0jm
oO3+s+1ycDy1/vuMW88Y74uRwaxCRawCSGJYl2jirRIe2lHMt7uRGRJX0jxupHgkTRIlS8B+KGLB
kUv/gD7WHkG8L6R7MYdb4tPvh8m2GELXTuoZK7ond6NGb1cUEXWbfNGONXMuX8XyY4/u9iLQcE18
RwrcfR3BMJne1sRacTl0DyJY6Zlac0LvGXaXuBprD4Rp9I9QF+Zb3kvf7NCYu5Df3FKyos5fFqLC
/GTHjzWpcx+ThEqQf8Zgc0iW44VMuoch9RBPsJ1cd+XUTlxyt9W78++ueULOnnpXqMCXn/nZAYuE
mwWwsc05LlX0XABrOUYEd3C8rmODrqqIa/yb2XfE1hyAjem2P1DjsTnv1Sar3icfkyOlAKrXm8Bt
kXTGR+KcAV8lMx7J8kkNeHMB5Rv/r5PponRbS/Y3TTyX3WxovpmIuLwqdfHEbiZD14IY5QJF0Ssa
BruKZFfHKL9VLHb0radiWmkoXdfEZWKCigHzSjbx3d98v9mcJZSVBD1AWrtv3LonmEexoB/SFM0E
X2z9b2KWg3AYhOH1zLEj0dIlFB00QlNurtA2W2fjOPQd2KIPcbP7QqNfUDwLNLqYkhahMmNs0FOn
CAkU/sm/UoF9CzvtT0qdqSzLGqYgNe7YOs2tHf6XZPAH3q+nTHTiZRBEXnU2m8gjyND5sTRqolZu
lQ+Ulva6DGzV+X9NtgOuksnnsJKuNf9QhoN/UCpr7oaDVrstQ5JLd4hw2CqbdzEW0IJOhQgpOt7Z
BPgODRCumLSyKJQthmPMLsKusuTrOwr+w54Sbj8lXjDBnM53fmn7c89RHXh2QFJteWyHyWlMJQPG
cEaworyPa1JDlkxf3SWOqXGc/vQyKZxtdzMqwvg5V45FNU8tYM1l46NPJgdXWeeNUv3yMyTZ9g2Q
Lh/4XmsEkpKMfOKxYJY73wtcfEZ7tRoZr/J1c6MticCrHAImt30WDi8ZrDusWxDuQ8XaP87LiNzm
8zuK75AydYv3hVMiAtXhwHv7kibBIdU6BbRyb0rwdlqB5so+rvsdBdMm99N5iLswvaF6scBTxIkB
TPW2VPtCSZ46GnLJE00lT2leCLJS2BKQvZds9MbKOD0yDMgyclBzChTdM7+k1eP6OINA2hkIIXkj
nueNvNDFBRnuKZaEgQua5qZuJ5ab4DUhog8vxY8p+Hjhi2II/TbambshSSpGhoY2JmnjZ1t7q6gI
uX1RhMxNKj3ixlSWincLFy1PwWo5FF2FeR0y8JWt3l+Ah+XDcTNpWOWdH3HXm5hw5HxDWArsfUdl
h1KOleoNyVMEE/DdbEdNBuybjHSnJCW3vJ7KjB/ekDt7JdoxYpH9W4OCIf0uEQdkQMPGn9c2Hlg+
4lyNZGyL4RIVVR8kSb5YRSnvwXpAYMt/1tBhAN+KpaaJIxHRdBjrZ8Y0kDAbM3Yy4ajUEtVWIY/c
7aoFmRwQ5NnC3EUCz8JlPRMgxIYySDvboNPdK2Gy5mtyg4Ze3BykA1cdl904kGML9eP/wrM7YqN3
g73rHjZM/9st6clcGnRqD3OZLel/fomdk74eHafRKJoV8pOOfAT/BUF0JhxnlN3dYLQl2IOSmRnb
9pPLVr9EQWAiJnQAkoxWTH9IZ2IKz36tOw14eCvFCVdKXx6zAAyvOtn2Uwp58CwxJnTGT+sEDvst
lAykXZVI5pukHG50zLYbbx4Uvz3jT31fgVBxu1wyxyYHaJDQAwobliZQIfpbIPFZSE6bgxT4m6Re
LBOIehH/9GfRG7G3hEWZx32AWtw5Yy+Ejx3oqo0PsSMnSd4mTlLMgkzgP5xUl9UEt/sCnNX76w5L
yVm1pR37MYJ2lQaJ1wQ/JxIgwMcfvgVSfO5f37Ux2UdWTL3F8pVS7ZLd+81FTvuIZ6VBuHIuGb4u
Xo0wMXxwT6q5DOmfQIJBRMTLd9Clik+ABEOHu8j30LwY+FDYw2HUYyEbgIBhmxnrByf11bLRZrIk
nTcEbzqwujr9PMpBHz4a/C/61AfHfrU6q96owhHYawWX54M7Djz1wuPtQ78BNZGDoba4DzBRK8JY
r+DLCr3G17CjMHlB4TNqq/6V1O3Gr6QHXydCeS/C1RNJVME5C0MT64b0l5RZKMsIYzwiZqKqhoTy
OWsJ/b4OiblnUaM/5e06sPYjdxbF9VullNjkxfyRt376xDbqKjypdPKII58ODO/SZdShlqYF0erI
CL5lu4n5tQxQKIw8dOsQfTg4E1hepJzQC7ZB+aG+cY6M2Pp8vOB9zMlhmVM4ko4VsU/LoZJNvsMk
PypiiX8Nkp5o5wXpCo1sYUsomOut3FEBu5CAbL0vNDEoB8iBtjh9ljjjs5vyYsgefsYwDnTV29jJ
rrAUZfPjrsgmOcWE1JCw7uPNZnv8ClAaJq6ZAKRA8Xi5Mhn/lmpI8lpiVQuqTuusIR4gkkoERGXC
1mtSqE/IQxCDIshsTVDXgWBI09ajb10sk7C7HsHtXglQUV5KixhjCR7EMQhrb02amdH8nUAagVLm
G2kMZPAapg43Rnyb779UQlg5QtIBcXiOpuGjiZjsb5gw1U5TBpnWFcoYbcQTOxqgyVaXwTTBOUCk
kS5lSOhamjJSjqX49P4s5Yl/hqNfr8AwAKLAwWY+OaDH707Sr1ufeyICwJ9EwolS96mrgwJpENEL
b9n2hhR+7yic5Z0X8GqS0VQgiaXtzaIXNs1TjA+9DjdszUrUDM52u3KqCi7UMAadewISrIKSt2zT
+ZiKwWPsP8JAmYcRZI+l35YkbjVEbwIngE2GN4nKvWd/pP7N46Bgeaw/+cXhCUn1HPlpMOcm51TS
+dwIp0J+MhvvUIDevkr+KSEk8nPNuBddlnqPHXykaEhOVrKgNPrPfLnn+91jWp44T500no6A37Ve
b6Bymi96D4VaELStNm6nnjbtsXvsXRZzYlaJDBvWDiqZ6j1OGDjLkSBq2QFz+WhYPL7Mc4JHDOWQ
plOuBBhF6dUfiG6+IohEeknW/G7EhFO7cdptpxVhfNLDuid7nyHb3rJ4+y9j27Vg+NQB94OvdOqG
2YE5/71dNVc/kX5ghWkyYHcO9RByP0Jpd0s2pYOSwouZf3Q5mx8rORE0XBkL9unTvxP6O/New9zF
j9QZ2llfRUG9hVtp3SLXVWmbHtaTct/CUMp9X+k1ZKrJlkO2wKzsw6pDEjqSuU5wa0wIPw4FMXzK
6VoYMmDL8gGSnguhRaPeYEARJoOckogebvWLQ390St/jHhSC0XdTPy06fTwwL915yvPrBSu5axGV
12hjtiBZYB+2IDlanIQg8OlFraR8yJkbOMSQ/d+UMKI1H3VUIyQ9MwG4j9NkDMnAp0gxlUt9eN53
ai513vavzfq79dxCE4RD7R4sF9saIgJnP1tmujtXTq1f0JBvtmeLAYBBvWP8xJBlW5p0wWtKygVh
Ecf992OYY8ws7L+x4awtxsptGNUECFUE86KfcfqT7rPdNSF5euOhUlLNvUFlLhQYVxldItKU61QJ
tUMj+dvkH1t+VuqzkyjIdw7aRn3nmDMarjQ0jUpYywpAtYHP/UnVneHjTpUQvyAipmtqHqCU1VpE
C61OcuN/5/ccTc49RjKPuMitGwB2yRXzbA36xgjja2gx2ZuCacZ3C6MZNkb+iNesPcLf4bbR7D5M
B4J/PiA4L1ZlgD65qIpn87K/Z81HXcB0D1idcH2/rtSl6AW4d73Rl+pDUlBhPYFbdN+bSGQx7Evu
TDtFDpHyKnTDC34Lm1pvs5xPFwZwKqGeXDV/RlxqJNoGBT6uoaTUa3RkyJJS7TVeHEQ9e3g5cqtU
jn9mNdMdnG1uibIggPgnm62LyJ3o30kYgxf64X9smoIJhOdBp7mvYA+IGq+RegLq75zhMbTZuXBm
zUElO5eDRc16xc0sx6gOoXZNKHDJ+F0yvS2czL2y0ZxvzMiGBuFRrg7PTRjmIecRfxQMQMNdOxSq
VfD2uGhC0/cc0Vz0kqkcZqVB6CweEOMN923Unrp8hmVWPV8kRBFxr6BNszxt1bcQbwxvMMaem9XP
2GxXs+0/zdmaIU0aguEXGohE4sk5yAaHhCCG0DuVwd3u1R+gT2LsjCySvOlBOdHNOoWZ7lH0aR0H
A5WPNflDajbQBNcB1yeN6IeuSLabLTu/7voU/YdyPuWfb0gUqRwxz3ok4P17TkZXVJOmzXfCKA79
AAI4JYiU6LwJ3wSq90xBAefE1TnC8S6QjQAROBFIQ7J0eQf21BDjE+5NAda0Zg76e2CrR+yrRE31
Lg1EBZtnC3YShZuCvKEGHU8s1CcRvV7fu4ZJMjqk1hLndfDbJjnbKANaC0WwpHB/BPzvNOyjhQb7
q9M8DuZOo/9e5ld3Qv9a0o9eO8y0mf8zd4KWVM95pCnxq+L8frrBcIN4B9irqV6+5/niy9iXoHNY
EijJDZ0ZLO96xsUjFEBnGCfhBdxmHZgqRoOdBPqRZTBjwRbf+T7dkKoGlEoExqeU62ERUTDXTxj6
K2gHqLeDdR8hJMy2gJVN1Txk5z8fTANrqaTBa8n9+pNXpk1qVMc4OaPYyfzIcNOHZbL8316gVell
K6T6OL77bEgosZ1tK5TP3W6QjNDfikKEKRLbFEPxYb2M/NejCv7OB1rHsZfo+JMMcCbNmbZc8Mug
appeZWARTWh+H6FfQaKlso+VHsxKNCACE5X3/sC+YE8gpgyZC8W1KPFgExYrtQMomKFnbER+5t5G
GB2j40IgZOWcOhQNn8goSLIfY+B/pB0l9X6R3SveUuzcfrP78bVWuKf/tPgeiXjOAAi8E0T0lJrP
EvV/dVQTrt+WlirMzZE1qDEqyHfohj0lEaas+xU9mVYFO+JofQTNglCE938se+t+sADVeMpjZ0Mf
1IhSCOeaGFHMzlD4wzGzE89Y67vnNV6pF+ghPeb7NI30BesuzJJaua4jvcz6WCS8GzRb1vCCNP2S
ToPusZS/9XN+M9R3aOM8zF8DXHzN2IM3HIaM/P+h13z6/h48J1zBRymbYS74sgYewJzz+n8C/pPI
XphpK+LobUR+hSoJ5vD/xWZVWRhrE8kUFvXlEtAFngBnV1tgmhK3omJnE5aKhb+AcCZGfFG+GJeu
4vctjTWU96zYt1mR1QYZCKspfNoDfNJTksaoYnUB3aatb81LdWpxtIhCCom+7dnReYGsmPpu9kkq
KePE9FwdctfAYIrfB/HE9bbJYKml6bh5s+psFLcfQlQDTaLm9O41LTn4pfDqKdVNJh5ut8esuI5h
gMvvM+xKUYDJYRBlDzmmAL2pkU4nKtuf86uDPwnGZPEyKIoHJYBiaoLVGVnTSHmRj5prg+g5muAr
luK8VeEK5hSPS9gH07nyJqJKqSGyS6uH05X9TLeRAQOneI4amVqEOrUdBDL66uG8O6RBBgxpeCYN
UzqQUEu+zyXz4yw19wN/VK2oFvTvEc+6afy4uZ5DCMyfdtvHYkus2M4Fhatom49UDAgPQFlX655y
VK+CZJmSM79n2yyUMKd4OA4CpWP8StKGE1XgkO56f8AO6ov5K5btytCLauTpVxvKbRjM7QCx98jf
YUhkUh0ip7F7ocxSP3MoKpUTvAvp8+x0Lt/+PZmxSEuXNx1yCjASaQAxjXb8lu06t+jFf+qPN1zy
Kg3wBnCJkc/aqocCwemoUaZ+1ChkFUgD71WpObOr+63j3kELMz/oe9EYAqwb2408JF4VCQDLOhDp
iTw3twiAu0569Tvub8Dq/2kSVpS89G+EdLA8tYC1NmJ0hXs0MbkB7R4RB4elrXBwyYjiaKrAGQBg
jWc+wuKP7p5RO/JkF0tLMFdZmgwteLt/nZXBaCgNa75q7C81IOAnJydqFZw76feZ5p7vwnxVyc3M
wzyXe7zrN8ogdJ7OJ5HDfUah4bPqABAUUqRnA+4mi93INKNGYeagnpa7Bc08nZbgNXCM4WtMwCup
EzLsG+6OxMQ1j6vu/Y328v8qP55g+6Zy1LlgOxcL6CqwEMPWS0miWukwJJdPsmInWF3AQPAubKI0
Gsrh/nVA5wKjB4F0COa8QyhglAL8RcfZ3jloy7kpcTlnBbkCfXjnG3McaaT2HTDczSwz2yEv9c9+
c/fp9cAaI/JHXFPL24KpkT/MWmzLpbUSNOwmb9cP2EOP6RNIFi1qhH7Oft4y2unwM/HgcSatABpg
07AHSNDKm/tddL9yPZMusq/vLoS19Y5w1jFKXJWu8ptV/VGhxfOfNeYZxuL4GnlUpP/aZd9EiiMF
qFWY1QQlQCcr9L+VZkMpMHwg0rooeigd7ZL3JDEOp2OYtEbN4aWdS47y0juNHunNeexAvOyup0ju
r5QUiOBjElZtsAcaup7EK459P3IVrLvtpw4fxV8eEtzskieigjes8Irf7nfwqaIVbBBYj1kY7HxO
08sf8pmeVh8OXyegsXtpBeQPcK8wX7q1CkPCPxAdLNV0Bl3yCClhRoFZVCAm2ezMp1ye/T+gHkyW
ik1NLgi+VzecR9gipGq3PXj/JXvW5ndKKSxIN/x7L4LKRF7mk18Im/oqD+AM4aGUCgv1qd7bI4hF
NTS5fW5Jph75GYRgLaLZiKnCwApbGqxMwQM5czvYnGLgBRB6p6rsWjvbAam72lbVQmhojJfFCrNO
xCZ6pYJNGSKOhopW2VOsA3UGsAGqifETdzzwZpoiqrqHjaZVxY+jQUOZeGJaZ0EZdHfk3AKX3UEC
jC/xqLRja6HnsQjkrm5ZrPYkuEOxxEeog6Phd1/C6TGL3zSaXGEtfKDS7q1I94Q8iuwigdJFR0ts
FxCczURgYyJxvXP8YTzqCDpSTInJS41E3pdlaYJmewv4l5NkQxzYkYpZPRjkig8jGFSvnBvStfTJ
gVIDOW2PyG8P/rXLEz/Q/Lm1qHzxTaf/CMwAkU3pYMLvyJi5qVs6TgWCsS4NSCQmPLXwqKzMlDda
wjyWRGohLH1N1JdUlbg8RLMPebjaJOl5aXKdzzDspkurQQOcacCTXZlbSgvpfUDblBCRK1xyB+r5
wvQFMY8yneX3GXSsI2pD9LfMvAy5d/8vn5m5ObQdyGQ2laut3EbMmqEHsMEB1ChPfpUaON+8KgOu
ZXRvPGau39HX6ocDI12NONcoYj6qiT3MprL9Qc8upfe/+S+j7UfNMijTx8qfkDCUYN5xeRzqMq8N
E9IgF5r0om0a/uSyp6sVIozOAMCOnYWmOWohw63zibl8tytpHgKacjjdUUAzlMMPoex8rG8D3OUz
0STxzOfziYrGIl0OuTVmNxWCQ70nccDbKyG7Rx6+n3hD0lYQsH+TzaPu09tdJGqJI2A+rqatpY9x
roLIvITXTcKr5kTkdMCD8EdF2I5cwEWDDpsiPcQfPmFiC8mRzSnslZVEjs5+mvtaUfpERDX/fseo
C36YBJd1dQo5PR0GOujLO9eljLPORVGYVFjHEDwnBIweT8alISUvdaN06q2Xa1EVfTwbN4icsFTe
EaXMaRlKnoivLmtICtdPRkESu7Zq/jHneKXiH28FuvLwAow95EDmEO3SoThVNuFSVpFLFq7yNqgu
k4q9F2UIgBvLCYTpJrm0FsiQbyP4dmlaOclhRkhqw/29nZOPO6G3Nu5hAIRUhQdk/KEhLYaiIOs+
GevBga9hx2v0ma2jrnS99R7qNToJguxBXgQEy5siLQ0G3dzsMxZbO7GOCikTqitM3MgQDqsuewtd
LPPQmZvEgj6Vr1L4Ph2PWVPuXJDzsP372eI4PcHO2gMXwtAAx4SPIIwPimBVOYiz+ghQm8uq2sLf
Y055ssXokXWmkLqA1sVoaUIpHsTxiTsZ5KpNtO2QK7u+WskME9nQMRldQUIU/hT1yNOjqDKx85W8
Ip5wUddI9XbXZV3vhFSjYvHzaN7vdvlAfSDr6wBWlVDgjhMucc/qFlzT7FfwjpAz9B4kezcVeXG3
pJykvSIMyGI3p/oZgZPodgIxKul7RbAAcpvbA1D96wbb2rFiW4AhbUNIX1wQZGCPdpoPQVgJ/qDD
jj8CAJt56dQbRiF8wlslJlLlyhtC47SQus2D8NipyVa/Ugfhi91UV7NTAB8yooOvgF3GI2dK2Xrl
De9AeYCzz76XTU5sRlzqEuGaP3XPrQ4+FBeV4Lq8eeBB3MLs6XXK1a2tKcDQOK35W5eRjP8vIhEv
S06teF9b0pQ4rTKGUEz75O/3jMJg435kZDlBbOWI8coD/CGTVW6DD4smMwjMnDeIDmhnqsDW4vp8
0Ptml86gVnrQ9QipsI4cSCG+vCMenNQ54qVUnJug+X/9zL50w05Fgmyn2K/XB3ZsKrFBdZTglNOR
fAvjzKiCZmDBw5iEE5LAE1VQ1CDn4o1SJumAPkbpZ2ITEzxfimyWNGcB80SA0agDo+eIrQ61tKqt
rMdKG03Hj+MWa03FKjnqWNm/bEhOaCdmHaZZFWrm9vndd6LAsqvG8G6Ltz9NV3l8j3Jf8hiNC+GK
TBh1OB9O32FFTm2X0Wppr580E4gpx/HlnzMZGA2Z1vCC0fLZLns4YYk1lCuFEjuCZpie+eHQS9mW
ln2Jmc4tsvpTkga5wtA0r8nfR/LyQBlChrwFxBY4dPnFttVNl7i2y+HaqHgoRiTO3KLAn+xP5HOZ
hfLDYfM4zgSzoZiaPg6djEQdGtmmejTeLXpHXxjGqtH6VeMOhuK3O6oZfJN8YwooaopK2jlIlFQt
3Bb2tMUCScgFnzl5N4MRdnoJPrLEKOT1Ife8g0uzF3G5GoIjwEXj3VavWpYGkHi+5FYD6IJLAXtw
Ykj2KuDsPPCsMM1/IUvtS5JYVcy5hIXHmxkHWof7AaEyt2EHB+nrqnva+li9SNZg5wJ5Xs5A/IkN
vARuIvvCuIx/aWmsP5lDVdCdxd5YC72He3iPL031GVvn7amYSfZgJCHxtqbWCp6WL2VJIIrg+aFh
DqUbjbxIZNm1Hs9yBULKyzn72d/2hyAiepEjuI4kcYw5/alklmwPJ95mojpvVV7w7uJgZvYS9/x1
VjWKzzJOjx2yUQjXRKRclw1oB145V3kuJ+28cGZImsnDUtwhGOd1pKFTgHcA4Fv7fa2WKQpQsk5x
JuK3ns+qU0pftgw2u/arz7QL/qRQetSM3LmecyHOJ4N1u1Q7KB/IACcaQ9QhksGWGtjP+w1vfzpm
NMBY3W/wYVERYaa4IOTpI4oNZvBfob9TDFSEvRRFnfqRzSacI1Ik9ZvhJIEYR2nYnX0j5EHY7n6i
xAtDNdMRt/CTGt+b/0XKuWivOz5A/VWx/UZryHsKSbOGIVHnUg1/ysjOsd6m2ykCkQep2PRwg0Pc
bwTuHv1vdmlcs4h2wWONU+GHy2VPj12Wxc+TR7iOzL/yTl9icCbbKBIukvB7DBJCJharXyGKjTj3
2TCxKCn0cEkNFTK+5lyLkDpD/vJB4Rz9fSTA6iwkmk1WJmr01U5VOVujO2zv91p/NifogDVWM/uc
2VKmkG3OpGBVRIYTuuO7kaStnqCh2FV6g10PcV0LOPkYxYHQnBJg78N0DiP/2kvJnZBAIYt0mTn2
GThro6LcOLgy3s7R59nqqTxrx7mO4eLZpol1EGZ+822CRO9bVUJANr5fOigQSogXypzmQ38xmb9X
Ib3Qwu0kdH6Z0VqWa7gv6PaR0FGjLcexSE82tmd8n+fAK6aaqqpM8NcLYTZd53l1YMSSHTNuYH9k
8rF5FkRKtk6fDsFiQ+Nti5t31MjchrnB9Gwjp4HP8I4UtRsAkCwmKVm5UhRTpIOWJv4cK40ivlnd
GxUc3lO3R3MVQJsA5cUAleqVFT/AAcyB2vrFyUsj5kEBnOrtga5hecR1n7wsobk/1TJksJ8ggEiq
Y/enyCB7pFn0IqJJ91PbFOLHYTRiWzmhqR99/VCoo2Qu4AerVbmrw0iHp/kHOetezOhtJaRn8w6d
aG2JQcObgDINTEj2vexg1UHsX1C97aEWuEfBVjpYZxPWYbl8Lbk+uemusSkfsrjGW1YVy4C83JPT
xMlSoEH8btjb9uDg8ezH/+RWlxa3RoYx61qTyrozMXDUV0REXibCn+fXtgf7f58q3S7wfQkTxusp
xKwbnEVVAwDOIEHwfntOOPC0AFtZLELHvf4m5jzBuumUh7EuIXjl5RWKbbfvogrrJh1DmrBBLi9P
ubxUbw5B5YweIEpThIC3J1Bt04SQHgTf9GuNAW8mZNpLrJqPPuFs6YaaG2p+L/4z0onMBN/mpIuL
A09EfGJGAwCBbasxcPfKZJSO8RFpT+3mK63FxuieKcWmb3aQStk6vs3nsYYKJS7gI2ySps0ZKFqC
4I8TxSGWWhWQQbb/T2VDp0Ceee53ClYwx2j66WIOaWuX/GXi8mLjcdpLzZnm1pzqafMrIb17J52t
xApADsMy09Ja8nBHjTL0ubn+w2f/h3FtJyngt/Sel3+7S7p5qRVJfByyRPsoFmlMEFUqMTRHEseO
+YCL1aCfIsBonbg+vsHxk4SfgGhbw+DlsnsF4brtmhtlxObSJOLxdyGAoP2kjsGP2VwaMJBfyOIJ
Knd68rmWZ1Y/xEadIgYm/KQT6LPIdGW0PeK/APBj0lQCXI4iok4iBqbjwQVcoXAxTpiNnf9gHKEa
rEEZBFZW+0ID15Sh6Qsj9pMda223hjPpJnrrPg49Ut1qL10kfAcmeEk2/50/OqXxfgon+TrMRb1V
x+TT0nP8gh1xV4Cde311Wyb0VbyIwIPUpa/qjbF/zXVRQstw+CLFiytXvKJZGai8CH+ppxmJ2G43
FsXxQ1JJY43ELCNCrSVD2L6b4AGrejc6ml0CqzwOidBPeudDnF9oSidlh/XPXL1Rq1yplfbm6cZj
yardgK48fKN0AX2zxLqGJJOCMABu2q2RP9baV+OK5SOZWOu5GWmw5AwO0jnNIb4P6VN3QcRaVSsJ
VPQOVLXS0xbsep3FybsXOKw1dThX8uJEOI9kNpAF1TFnOFxq1IJ4UUSuXUKJdGFs+a4EkOCSBSQc
YqtunSdiSlg4eGjEBCXlE+v4Gh4wM9E1Htv+8lQ3Xq36iOfiMKTdfgHmlkUGhcobv3aU3tnonrDc
7T0UhAUN615iZmokoiS4S4XnM34MgChFT0e9izcinlKgErP+A1vt5SWjCobeBmhI0H9M+JLYHfmU
ZgDabxUipp94ykVubwtSvIkGjYhn6eR+ZjdDbYau5OJn0psaOrxXGNevmh2Bk0krvI3WZCkA1JUU
AdcGaVnBxh89XRiu8gKe7KeTzBg9bUyp5cyUlavqcqs/XN81pa7g7lBCCR4Nhtj49HO/wPzmYJzL
2d/J28oqLPQ31mXenso7YwRETvU0jXKFYg9yNGoAc7sEJiFYpF+b75qR5z9qz5HytYFA10UXIDC5
TSjuba7wxwMUTNEOj0jk8V0HabJl1djkLpxb+Tl3qcao8DbfIOCEYfsZ2XZ97vyM7pTIYUBoxJAY
axmXcd+xzYEdS/rZix+aqF5oYg76NLntYjg2bAypxhonzCLgHEe2FM1RZoYdM6sFR2H71cz55PEq
+OIGhQGX94mW2dKg5sEXz3UdM0U00X7mpYOyOYCM0tVGfTQwSsdfVlUI2OeWxlsaq5vTZ5wfF5Vt
HkUm6ggYCeAie9VGRcu/L4x7R4X0IDk6yfat+GUJ5kuitkAnDn4H1Td4CC3i5faRmX4RU1uSyfgr
q8MTokmQ0qSyCa+4yV2C2MwsZYdBvdP8ngUGDRfz5AQtgnVEh+ZqLmKnR2XYc5aW/CrwU0fsGYMk
IrpS3lEBwOU+kJQRr1co1ascd3JRBzDlqUqg1dAGDpdGcAW5/oYcO33jNF8e4HL/QnR7TPv0+wLL
Y/nKl9FFyMWbB95aoS6sYvNdeHyVsJ4idLXdn3LhaZgEYRxsHBuXQNS1lUzIzrDfhxRI/0+k6UMx
OwUGkVdR10juEhw0EQ3FIORTQnt3WqD3VgQgQXnl2lEtORGHYI073DjM0q3MIbjFdWNVHYvT8O56
O5sgXrEl8QZd+F5oVbvNqic4Xp9DKOdXZvdUc8A2jQfcy17MIHi5FjH7WcSOw8SFCUvQi8aeFD6X
ytOFKmez25xZs2cn5BzP2HcpbqyDU6JFPC+6BKtwNm29IQ+BXc5sJ8jQ9En4NTb8O2gh04hUM3of
ajH+sCQFLqecFl11MOi1zHzo3cv725qoqrr0lWSNjiNnybjzRiaLhhaw5bstV/4eKmxYRMKuGY1U
ERsOK4Bmq1/H4AtL76IDpX7Au5PQ+sJ11lxg6l1km7Dmh1P7u0Wc80B4rhM8vT1yDkFrQHj0sDrt
BEnHGnHuCSyipvtFvf/SDxYVNtznclzwEK7SeqrMKxlTS6D3oASh2Tzw+n0oigx4DI42Tz4wb2A1
FeUWhO4mhmhaXSPoje3wb88NHeT7gjWWIjrk5J0MY6CkKrYFQDXKAgFdCThHuAqQTxdCliwTpNkM
Bw0+Q2LzbNV1UQlrTwGhmcLmhbEQoEzWfq3160GVJFsWFNvijxoeJb9xSDSz2zMDkXsTtuIIAllj
dc9EztH2vWFKuSrRq+s0w8T8Up+dL0UqDhIk2p4uQInAFbaQr1MyUMkeVjfS9Vin6FBcvqH61GtN
UxXFW/0LkuDrXa+51AQIOsxs3U2PeFpEHQLx3Le8Y7J58KkxBAJJPHP1/3BfWcSO7le4sBhRAn9O
+8yZbIGah6j3feHRlPE3FW6Xy2nJ+HQbRt4MtkIgK7zh5EoBDCwykGxkMweWYcCLZygBr+iBpktE
2bTXcT5c7iczRjFhncGX69zDESNA/1LgN5BwOIQsFA/QxHYsJppDoM71LzqogYbb/P8VZCU5/bW7
pUTbQa/4z8jjUyl/art+bA2RigHSiy4rnD3Xfuy5HfrW2Fn4XWeW/9zPtlNo83cGk042GXdBIdhX
45kk45HAzc/hsW0bLVpDXKCT3LwLjCO2HPVnEJYuGzoL0rOi81MEIvpRsXUbEZYXGMejy0lr5nHG
zZeHIrrm9Qh3PAbTpFVjw/D4kz634cmxYjNHLbSSMZmZXRrKn61JJNLbKmycmMh2kHP0QdPMOnTo
7k5Rg4Cbd0dX0/y74/KThDTW0+Ap1WUCteWtXY7BapfcJUe9RkE9R0ds6mGH8SUnPvD2YtLoQ8U5
+nIcAZBKySXbobx+MVStOeOFqUkkaOcpNO5XHZ7up1bzgBMIVjaZHHjS9d/CSnE76+M1d76CpzFP
8Wiwo/omxexVB4FsXRRY7DhbwBCz3s9GfUbd50i4dDcL6SVmOewwGqNTAnWanJLrLzhb6Lwu6nIe
GtJD4abt7qSp89i/PsAu5c5yVGvTtP6CCuUhqbQ3gYy/cZVAe4pjjRXDzfIR+k1EWejD2IrKq3+O
lhsHjhSfYj/mUcXb2vmuu0qA+Ue3pJJ1TBf4y2q2J1DaPrgyTcE/JcgnO9VxUtV8+tTqSdFP7T9D
P9uFoyfEvb4gswWj2JbeIs1UoRjeoKKZcT5XGoJXkstLqY2Pg/28yNI7mbmwZUoZDgLWh7y+EUXT
QbBMj0YmSMrf8uS3drbZ0t39PXd1JunOpP8sj5zT0MQPnssPpYdA4K5pi+rwXq60omJg0Hiwl1iC
jyI9IrtdmONlB1sNC1idlNW/EA5mUMkvmsZRPWABj/GKzbLnyuZGY+EWZ+txTpToVE1YyoAwhLN1
ivJdRTO3GVhXwlGzPw30jfsbEqHarmv+IRf2RbPz1BoBKPoHbmFwSg5ppYtb7jpnDB2DpC1Oigrg
olzkMzILzeel3kIJdBRdg4U9B+5S4ukfH3/Qp4Fm8qv1wOlDkM93ZgFaneLbah5z40fTTMh61+nm
lQ4NzAf8NT1rQnnESUWlFjb2603qdLqmUzzQj9bKAgfHQDmMInXXqHIECxf0HWBLVMKEJI3U1vEN
9CC6ZmX9rXPgkeVVV/MM/woSaks/sJhJQm6IJ3hqdj+bvrKwuQ3DApb7jJidnKxkMfrdS08oX0b9
mM54z3G755+135p3BN/wpFNkDNxBrX5dMkVXcEZx6Bvcs+AanaFc4lix4ZsU5FrAJZ7Gb6V4EFkI
XvZFHN9cermXjvLjAbsL/EnCMtLYMjrcqjd1fG2UB7N7mUb/NuRy4iOFCYPjqX3Pl+aX424eJluf
6kBFAWcQ6BvjOEc2Wr+5S2CNxeBd6aoyIMbwZRZ26YoouUhDMdO88/0byHacT7fiSKatU7OIeo36
/M46op5ViIhSugf3ptuzXFW0LOpyzuV5xp04uODc9EU5pKv+3kWSkMAeGRQRl4IqFK5lBHXZQt/G
8RLyTdCWSbnFtqd8kuTE/yTfnUH9NhQODYxVenFG61MwJf2XJeXitSGbsRspmVOOinARSll2OH6N
89fmK4UyGob5UmqTq+o1gT9mg6qnN8vP4tGjMTamXgfiSahiY0nw+qyW5uKV8u9RKgc8fhCot0nN
oSjL+ABShi1xRx8JgmpHmyukEFAa1xi0K1O6wUScFxEO7h3jJeSJ0v5AivteHbpTlmpWoMYNMClR
c7wrFh7F7OiGuHfcBPTTYeqE7Sa8idr1E7JtF1mlgp+oh7CqD6tYu1McozLCfTIpir7za3VoTO7g
valhr/LkkULBQN7FtO56nnrxaVNRADTOj+XQ2KroJhKrcMFEA2axg8KOODu6jPwrpr5iW97Lxpwp
FAHmeKVq8XZNmAuHgQ/VZPjXEK99+ueHcr9DVJzXl0btDWSbAiPHh3mizZdm+OXgkXFui35whTmj
EnIIc/c0eRB4vEpMTXsk15K9WNIgVJQZNSSlnqTEv0ei/WY/DD9t6r7VQ10m2hZwROPO9bS9R94t
0gXYydpYrvPE7gGrY06CS5uBhQ57svB0ErDV57D485kPcK/RRhYq806MPnUwCOaHaXRj3tJcG1Wq
RVIEsuC8VRNGpusFKS4IvDS5Uh0kXqb59H1gnt1iiaZrnsocrmxsr2BEVTKsLAAX3d3r6aHCVdSm
R9AZDmbHgoO33I3EvXa/1ezuQBo2oSw3IqNvz5rH81X+sqyGoK2761ulDSj0JWyJvfjP5Vxp6Aie
lpcA7G6/O67iDSgHT48wBe/Up2MaZZqUJyu3d0mWEZsyLX9OR31tSYyu5IvJxBk60h2aCFj17jov
7VXGPW/1tiiSUugsqQ9h/J4dRhTupSFHkMQXp1ZqPqA27vxuR+/RAN88W9YDPT0UOZttDkKBX3OJ
Q3YeTEC3Gq4BPl9vLbwEapQjWxjV9tQIz06biXXcXeyhmeLev0+ZRFD9xGT88OxDkycK7HU+pmmu
x7gHbNrlyw/J7mAokoB5lJN6A22rlRoc1oGVpjKW8cdLnS8dgJD22pvGbMEIgrqJiZGPslIoBxdf
dvWRs7cAq01fL0FMZB5kbvIPowxEUiQtt8slTwG++48pS0xXKgvs1WwE2Y39Z9uNAShW1gGfRwbq
7F3c3bD8cF1sZB8nu+mBuRa5dPsO0g2MeR/dc0FZcpKE2LMfnMY12VA+ojxaFUigkczT7dCXA78O
kwAnWdVbfv3thcCCLcT3pE5ooWc1wP/eaGwTm+c4fCPlqL1RSW2en5C5Jp8raSz6ryNGcet2Nuyt
WKwiOm/3L4irGhFv2ys25+93QIiIz7zC7jmt3LyrZMCME3yG2E5+zG21zBri+CJowdbqjdS/cliE
f59rOmWLe7x2hZ5epWhAycUv0QHXeu2iYQ9Ge4jYUJF9G1ckigh16C1nElJVLDIGTZNDxquFHtlJ
iQGaZL8Kjbrlee2TnZ7Fpq3EV99fJ8m0mXvwqr+a42pu+8wTeBX2PJ5tQOQOvC7b6cVfy9D/Ff5C
W5ewKBpl84WLMzp8qIE7/WwrHdWaEpKDRG2+EComfkT40X+Fiewmr5bfI+tpAocm1cDsGrIwXGI3
J7XaXq8V7JtVY5sgXEM/wsX0dKWz3tYSDqMD0t5dPwsxW4xltlo3yeBNg908jq9m6Xd0PHGzRH4D
2VZag20kknmZSkF6bLy4wQN0kHzYY1idRwblBF4BjP5fA/EdkOWkrgPJAynTM1yu+D+6wHGUrz7x
EVT5tuLjVjEfdXeDztx2vzs/djKzgLaNiJeQ+2ZZwIQWvwQOGBSFLxeg5Pq4OJpRPzxwazD1ZGto
ZwTYohUfRj0ZK/8Y/Y8X9eR+h2gVO0Z++Xtex88gdwjrihlQCzo49Wx8upoHN6e7ipm5WKjrXANG
FFUyYwvq0vOY6RnkVheXuRUvH7tlXHU6e55w8z/qcwfj7VWHLkeA4KkN1XRUU++eYpr0Zj3TxoXa
/BFFy3Yt6pKdHh1woIzOPJ1MUu0aGN3zK3UG1pdqNoIzZ9y7s7lzMOJs96OGJAWTDCDiBPcQ5ria
59lYv65G2kMCNHv/0OYcW2gLOuyydiE6QcMrzv6f6Ol+LkTaJzZpWqyR79cfN8b+Uk+BdngUq2XD
F49Ey3ZQFiGqLlPJ9mipxpkto4LwFMLmEyJzAgM493ZkiHGYNIkx4wrkz9PEfHY1iQjvwmjNlr5e
AwS5TB86bh/6Rv7OZr8N9WWK/4CTSXTt/v7X19/Kdk/Ati1YXKrjvaaWiLpJNwXPsdWXWsIQBMTj
wS8EFu4XUPiwk/SXTHWpi7ZR05L8uNdK69HTjtZYHt0ARrpiUOD5XiRs+/thiYnR9JsAPXMos5SV
z1KIxMiExWlIXovn50RfSeJoN6SHUzXBCiylMZqehM7TM1C3IiPPuAwTg4YBXmMPljMhXAbwfpla
iJyOQ0OtvDR6f6GRVlIjrs6Go3ehNRRvyIP5rwqyxzUqE/nsfwB1bGvEm0NKDza3aRPU6Rg4HVxQ
54/qDt9Muufb7CA3cfhrjCGCEokP0IQDWvp7Arraq89f44B1CwWdQri5BiItz8ScJJgcY8nMK6g1
7vhhcXwr4Tb6a50rGsNHBVYzXREDIYx/1V6RVDQ5WxNA1WL2oz0Xdc6kLdi6TBHm93Vim0ftHhON
L7NNIDhu05sZbtGhTjm7t1NuIP5PAgxojk//gUrkEVSwP2O1vwY+nQHfcwElDxaMDj4e4wJQJ+Uu
09h8YPxSv7DOX/Ij6eGfFZFv/BaCEXpG0Hib8QkKYfikPveF62BtpdgbCZz7By8JY9ntmRFHfWPr
Z8SYhEuh9qIfcHTEc5a2uyv+wL17tCW4pXieABas4mu/RBUsxBwWuGd4BqvRcCLoFhKJ8Sh1aScJ
MYTsu8JTVtqBKp5+CxiUTT4Z3l4uvM2CgCCoWmibfrhoqu8Uhqy6sUaorocLeTRLeC95Lq2IjamP
5ye3sAUCFTYz3NfZL1VzDqxdCJCTX0E6+AOQ5a5nvc+gyBoD7DSQzArrymX9IM301JlOtAYZStap
tr5VEdnFRkK1WxKH193dlX6UXx4RN0lOA8I9p43T4qxYSEHqGJTrdWvbjw4cakuwuc9/bCGE/++x
RJsoSeuDDCyIBNFmXyjglSy+KgUDTupjePetEAPCPL1durdkTUKKIhEPao/G9ADE8qTZZyIRE2ZL
H5ibu2B8qGLPWp2UWIx7LGFrkxd163m55UZX3jVG4fULM1meT2hU7ZmwXvrx0U9wGGBjtFUprrPs
V6aqNcefYxES4fgJ/OHR+g9kiAIUArdjXsR95JUTrialNjwC3NVfmcmfha1u4s692GHWnJ6VMCdC
u0hMggKoZ66pT5TxjzAkUMJ8SjCWjXLMHpJwynYwtmIMSNvTwP2oeMhQZHrQ7ywMcaPcHVtKEQmZ
HVO0K1WsJqsP9FgT6OZSPC9KWwBW4ElZk1gfitCnamO0CEd9uh+qYIf1qf49PsUImu9fGqZfUr5Q
owDofaAqftFzJiA6oGhGyUBgDBJafTHWkvulkZWdTcHUvlE6uclF5wTrRoUh+AvzDrHHJJhRELor
z2i8+1aU1Z1AudU3AQiekhFb8jX3ygm2LJ/9nILs6jql2p/zTDF9egx8sVIK+bPsS0AbcjzvUHND
DjbvByByo/QtgaQLJaQ+ZPwclTShTnaOXGv5/sQ+eRMdBtKjfNNMiPXvJ5XSe1ESV2yk80/Q11n1
pj+0NVnKQxYe+9B7UDMGi/dygIUmCDB4eKgPYj7c0ugkWFS3nQSdOM9XpD04qkq7n6VsA/rhoV1l
AjBUsO0ktUjqu74YuoGgeJQGXbiW3wlt/9mPilOdPzsjqbNCV+8oLNyL6Vq4yDjuuXSLGFTpnbDK
kQiTP47duqCI36b40TJBXcrF3YRAUOvzRkvB9b5hfupIA0OkDIz7pxLvT50CWN1zd2SVCECER7JH
b+8BlaNKX6eHvoHLPJCe7zBHXQAD7lJysJHxDbwuuu3pkxAIEWRkYZuuYEMAtjhsSRfFNEBN8kn7
s80MQEAifIZRPZ/UF6FTvQywgRmXOjtQpSCRxGfAjE0Cz7bnfjzMsxJpQ8qdjBX8E8SArN5j+Sun
p2qmJr81D8cmLXZvMIOXPeCxt3Bxc7RoZNLFXlhYCg9SJaWV3FfkchpeDjVtqjhgc1vfOZKT6EUZ
EbFHsIiLBeUprohzO6piFpMNxycytgAaNlQTabJynNxfIsKuH6QEAfCaSin+YgARovuRljF5hgfb
zn6H8Ignmrxm3lhAFxVQVkjV3qGfWvJOugbYPOakUIfoub/0Han5/iRAGgxEDS3zvEPocHwgq4ex
QFvYP72kdWRpl6CQZM9edZIpZM++7ZU1wLvpoUXTrLKrSFG5YXL2ujupSzO5kLYQymDbUf/jF4yS
q2L1lF7bWT9umS8vbqI8dXNfL3mXZvYZzZq8lP/qUjbNKck/GweSt6m877TLwhqel7ODlGqv+SAF
AqZNMIOfE8ksGox4AzaGL1Y4GGOKFpVqko0MyFY9CqsiX9iQD2GgtV/1B93dykKy2vh84QN3ruGg
e0WfLGyM7tB1ftbFmzNNXhDSLw0Z+L/TEHym8s71t3Nho06bRXihI4DFk46gCtwBAgv8oeZjtCeZ
meeEy2k86n38zQ0aGuhMA8LxqaQTlmBevHxOpV3BN3V1wFzx8vWsA2xJ7CYhAZn6+fLiu2SrfOkF
OpwXwaetAdKL5kxiIbnDX4JGBXK+ZTIPlgfEx18YTtjNLAEa6xxfr4FUy0d1x7RGG3fRY7asfhq+
4+rCA+29SLDg2U23OOqG1sqmawHAX7vhbUJFOLhKc9mnKVS1wSw/r3RnsQ1nHfl3ShXCVSvIdltA
7GPXhWsDbpPo/SHiWWuyDDjjN0jimnK5/1Tc/IHyoIsTo1y+F6Nwijpkl01S48Bns2OYYGhLEG5E
2ia3uJVBUIAq0X2QSxAEKS1w2GK+eM1/ADq+karMGybdxAM6R2zDHOGbcJyvFZRJgRhAQ3NOY1vM
LSFjdpMyUmChLD8rS8duTB+cO+Yn7rw56/Lt5Aw7/sijDGtr12W1r8EBAKmaAZJEtoH5/BEbsjg/
bLhP3jILrRk4T57s1qdA7CnaqWEDHdshMQ3/rIhSJlzaBmNlH+nyR0KZb0LH5NteAdYLhyUg5YhV
OJNJC5KHbyNQhfGmQyLFut6ld9M3I3+xAAPcb5zy7OSmiQCHyXNDug6GtccuXcGfyUpjXhdKf82Q
En29mHEDDe1UcLqFfhC5ouWcbq2oILu7+gIr2NSIDb5PEAp5vEolDGKSku6n5U2rPVdkvYxcchQ1
P4SILIMcCMOQEX3OPcdpB6bG2OjI7selPrlpv10OQ4u23UZTXZkwoQEHg355bLJqR1Q7UN/w/GYA
w1Tx49pAOBxUtmcNQXd6YRIk9PN/G/pyHBo5u2dVEcHONppc8MMJCkEQBiPpDv03cu4e+oKAWqJ8
vAjlLWjhRxLDYARzqi2LHaD0sQLHPA2dgQq5RZcY4LNF2zoJzidhNMbUmm8f4cKkycm91Sau27eb
kN5yMLQT2P3D7KP9oAv+R4c10pvatD+uYgJuqKU0XeWpJB83FhfyLlNMCCUqASIA1ALFtYdUgWQR
AW4R0ImPAl+cjCiPW62ltMDHbfjJeP9axkbehHm77V+sZhOj3ZJ0zjgBNZgVKws3lmxPq+juPz6+
enhKOhGDmm6m/pzOeauHQlTxqoeiKy5dGmzTQowRwxjFpwDChejq/RDu6rMxWy4qHvo2HN8Z0iE2
UDENgGDN5lOolPzI3WvIpe8OH/k87wsXVR/pawpUPuYFKXQSYSMgAD8FHIhmB3mJkDdXfbsrYmyn
k5IuJHKaTFHySHNb1p6y2QOvRd98EfiWKH/3M0z/zXtjdbdTVMPmZs+CFpYUJp1cn+I9VQ+v3zaa
4z8e1DuNHv3SkRmdV5ACjGoxa7TpIYp7cSe1YIQloP5azGj4B0Bwe1fajai3Q1pzwXQuQ5n2Mqcg
sc3pRd2nxLZ7sY6+VpbTo7c85FhjcqBAArnJcxWzt+WMN9sKfklgDj1OOsa+3FBaH1BN4KlS4+Nv
VTGXakbqQ0IE86Lj8YwQkQ9eQDl0WoHMGyallIo80f8JjK3W4SF32vIuT76K1QzDna8x1DOqSztD
GwZlOS1BX2vok96DId6DNZD6Ocr5yJ46q2dAQZ6jMEKPHJaHa86dSOQfWsZ/DNh2km8Xv4rlO5Mp
tC90PdTx6NPdfGrbAwS/YLNPH5+15QMAQBsut7ZTer/a8PHxIn39mzet4qyrj4DHwoNcphLVfLIi
AluokxXAY6Mzpq7TQVD0yDl7YHqdocXATf0zqz89B6nhg9I/zcAy4E4OvU3GJ1O4YZR9Y8WHMyrR
mxVsoP4OZC10ANddfCRXYSDtY6JJ1fhYTI3COcNhMrQSNGql/yhHKEeVh2LRoEcyndHHY55+31yL
nPXoqEG6UHAy8InQrrJlYKBjf7SxSGApWkD0UNY/Dj3S2Oo/4fV5ISSvW/HWz9E84gxdjkKme6Gx
2KHorcZOKoeW6whQA29PdNc9CaaGvlsLAFG59AAbrfzpRBbJjYNxXkC1RhxByyzqW6+Ok4rrveeJ
g4wT/lcUpNYkWUF9jwrW6Kn1vSs10Mxt4AKEnSWUzEwQ7BNbyKcK95RhWGi5SNQRDmi1D0sXHTU7
8cq/axuPL1c9ZJXWGJQ7nTkXkaVtnV7x5oL3EjX7o5oGRfDFmL774arn3NJn3AxS1z6zc5Duxmxy
64jTm66yxVzOhrbKZElpOgVDJ8NXNKqGaSC9QqNRdxCu+Yh824iZwl+rsyV4gRWfUt6qFna7ILFS
5BKT6LfSNznISC0tSIZrPQ2mIolgtdY6OuC9PM5a+MJB+eiFUnBJ/DVK+FKT9haJilwQapquW1Tq
K7fJ/fbQ6sQNFUPiOla5X5GS1foiA89sn0jngl6n7egT4IZUGf30M5jibbr0QTUx6m7U+tWeHhVf
OzFds3fSuz2v+mHgXMdfClQFh/HTD9GDuT4NIKh/rXCNjgbLY7Ff4s9fRAsQaXVNiGmWB94wdta7
NdZjVAnHX9bDSYfL0/xM2B4u4l+ZHPbzRcCgWBev06Cb0gVPw+qn7mD6eucv/2LQGiyYEuF+sqsI
ymbLnJyLfg1TXkwKKFIsa9Ybn9OA88/kNyXdmQA9MbFyJkEk1ZXhgfK/gQL/elmJIuC0iI0oEifl
+XZ1iI9qm96HjgiRxoSw+LN75YuYhKx1/w6TEjsAKMsiFw9AI3EGdZWgyCQMGm4zXYrPXw0oxhrq
Td9WkSLpqbJ06Uu9sjXYrNc2sjRROtzaAcyIvK+379QQ2RvnCU3azWI79FpaCLkuRsD3xDiesGlg
rTzMeTN+3yA5C1wNRx9NFPeldA/Ks15nSpf7kMsHRhFAu0bWsU7un2YEFiU1cPw3RjmlRq8Ln7dd
gX2yY1VO5r5RQoitm9wP9Vt08ai54c4VHu8Twv16T1rQys8RVOuKFWt1yc47YxLyaORcmbER6fKM
kcXLBjTGW+8HEEFEI4IIderFJaVB/6muJZ0xcfCBC5meXS3y8PjQAsWIx54N5JBW5oLub4CFyCzO
C/CkhqOMT/jhyti1uLfIH+BkCjc+85z1L/S/v68eZr3Kly84sSY/wyleT2OK8l3Z+m8YzHYmEYpp
FiJz/5N/ZtM9WrRxigt3yrpC59VnDKceWH+Tnj1IL119J0f7hPxMcz8fEIfQx6EZuFP5tt3FiT0u
+quQDqjQGkPReMJazGoGPeTYnRFTcoI/rWIuyJUmjO5auy6bOTEmDAB/cg9qp7u+inL2749FU0mu
8cWCEvb4z7LotV6Sco2rK8Fq882AG3oRDZgjkCZapYYiaC3Oe2oUMjCmMs7fkKJ1FEO9kvk5sLf2
kCQGK1GfcBe4KHl5U8TlN788vXeU7BDUEwkxbFMAjBZwiQHTAg6JvKb/bphnusJ9U5UMq38W/jpp
ZoIgsnabuUH9GjvaZe0PzsPj8WmKUI5k2tja/pp3NnhcznfmWjpdTZv+Ou/t2PPwwHj2FM4pFswj
M2UXdPMobI8+R46U+bTSfD8ayXFeoNREfdXviifajU2okRXe5Nlda143meCpESoX0nCeubMHE3iI
J1K7M1dKZCVU91lX1NnqZQPt0j4dQedbLG0IH+4nIlA0xDCBDpoqgGbII+fdN++8hBDBuhULsE1z
eMzzMet1bMqIvkN1Jr3nGycAIBZpED00uejVHTiWiGo0OP1qdi2gCsTlo7GXGPSV4cUR0BleGISx
InzZex8NtMtN+Pup5hpA4zr+mgivzJtI+Gbk0OiyB2tUN+X0JjJ1ZWtv1ooNGlcpbCaz/rxaFnQq
iPxqglkrZMYm+pk8uEKl+u5EvpXbVtW/Lcw1bKRpUJFA8FHgM/tn4FcWGGKtynQ//Ya8vJmmRJdq
Vlq2R4/goQHZHS5s/zKGWyexyPH6oIllAEmtVypX6FztZ4Ssz4jnB6x0CKHx9fZUa+O3wl+fidH1
Szd8b7axRmmW70xzoRtwQKSLeUS7koYf3THeZ7DNW6duXbKtdF/bY6uZPmz/Ic0L/w1yM8fFfnk+
S81u28ruzZoLtafdyt07qb1S8/Yi6v969Y0A3wMj8nzfTXtJCTuRVYcp9SfHWEgn4WjS0UAPY8ft
wUBUSwPbFswVlZ92j6nSmDF/Q7WUpmlA5lWr9c3t5mL9ZmqY8ANUQebjJMFpQ/3DJgIFPaQsjmnm
w1lBIXIQ7uFN9CPSZw1zI1Ykxp61Xokax5Z6bHnE8iFTq6UvbAmzikiFgrtBL5ot0wEsNVCRNqR8
JnqBn2scYVHecw1quUgCIJdVV67KH7HMf6T/VEMytQa7V0EqnDHZCKyfX+S0KhaYtJIq1SUUWRk3
YX1/gPsz/h+qbzFx07TJzc1HzQvpwLB3gpLVsoEThOet1K+Sp1vbL/pOXcw5N8TFpiabKGK1jYfd
Zj7q1pdHvksENSBY/CpbeC/BJADCgAz+MXFPie3eNBWbrhIn1+D06nvMuwkHXQ88BHk6pdZi8EqD
JtgGD5GrUpBw6LM/pkghglS+TG249x9MOVK71fYESUexr6Ts8MhbLoPQ2OWXYDSbtE2A2qPknGIP
X2lIhEhIgRilVXCVYZ293KWcc/Q3wQEIIILo4UFRqy0aFwq0hbLba4dHbD0ukrooPg9Ej0c697p3
Izbu9zRNSLNP1HQt0XGt3ipXEZpao1PYPJwhN2ScoHxaxgFjdIPCPcXqNO0hem3zp+j60G1YyfSJ
dtKLhlGGLR4hk2Qzrfjmot9LlmnFdEEIoGZ0z7mQ2XwYSQPv5yp3CDtuJ7Sy1OIQeGOClFYYF7KU
REDO4FNHkLvQZGf9cuPoTLAFWaNfRUfnE++q9aKIS1uiaoGqG7rlEju6HCWV2DiBCr76f4ipKhBI
Ga9sst6Y/34dey/I9MutD9hmR7Vz0Seu9WW1KBF0AN9pKtNTqGZH2O0JG1Zl3uEaa9Ta6N0JOSjs
fBbBjwIDb53NSzHBQ3tCGZalw607HwQZEnTVOjBdyuzBg8HH4BSZuAsxhcQtcJJ0MBTLcig1CJUQ
UpkQxRxwUPHgm5mvSCErepvuHSXqxXw68Ell6IXJb/l2h5GpiEl668ngzqsJ8l7k4Fz6ST1xVV/5
Ckqe+LVjfEJYTL3nlDamFwXxJst6XwLOPRLw/yya8eHEnpCbKVFvavhzVayxkCXjy5EN/KiqPY4t
Q7AF//8rDnYLSrk/s/o044rBXdj8889+3QNjxE68z1r+/k63/KZgRnPny69KKJLKACIGPsEAr9qw
CYbkv14aKOpLlnoeFzg7RnGyq/Bte3Qq2MOSqO8D3hBd5P87F32E9Z+iQqCFunknsY91jhmvSCcy
UWIDzigYoq+nquWVK1zcG+n/DmGjV59Oy0tzqE3OGm/Mz2F0M6oMLbvALRR+ZA/YnGEKDZcN1yIa
F1XV+PC8JyAqaXpujrGBETcSgTVLlg2eUIz0GK319qklLqqs9gb1RfwPnv9OQh7MLIJFqsI7mEyA
Y9I64bkHrxDzz3CEDyXrQaAYlYcdRQkcyDKpC6sBVAzly2jTal/vBBCsZOlgnm1WOujrIzkEQfqx
fV79tVrGYBgp6AZccUgdRDn8WZi9NAkuCrSGqLNecdtVn+wJgjdAeOWXHPcjYM0D0M1ZeAzoLfrf
2sY9Tu6uTBofYB5D5siviFoX6Tq28mYkoBHdWT5gQr+SvW84z2tMpVm1vrTo08yCkGjDEjc4RhBm
QoiPrh9ynUk8UYCln68QWxnh1furQJzG00vG4//LPN8BEUNRcX6IO2W3pemVIsUXmD1QRnKGv/yP
wHr2zB7uObWZMf2g8IxnKW2MEGWd+9pJhd+qhDYExe5aSdiDMHVD66CG0sl1DWC0EOK6rO2SKjN4
hJSyM2mKAtrDEJLbK4sCqet5no2UUKlb4/TXNzTf+/fuI8wELzuHMdnOmB7lhvbeawgskodIMQnZ
6Jutccj/uUckg5d1lV6uJwLitqaNtZbxhUVL8wDnJXj+v74vIKGUVK9CWSzDNgtXdTC04xrtMNLc
4aspGvTaSpO7Qu3PSjPEGj9CU3zYfb6qq2a1CSfFqv5VxXfC/BKjFM3rXSRdaot2dm7y2XubgTlv
bh2nkKsqhE2/CU8VPPHu1S8BESR2eZiFPQpGeYYYXf76hRvDr8P7UNVqqWhJmliVZBv9APzDJ37C
1Bp5PqNgTEIKlbRlFN9qmaw1DrVAdeVo2aONoj+8RHksm5DuOsixApEH9IdXaKAsPgenmBrWPwoI
Kzjzxzqmy14ch+5OANw4tTlWbhbb+xuFPs11nsx83hZ/oHqq7NcJkB3UA9DZlcevSTG8EJIPmdIn
viYfQMascSL7Q4AuTkbQpDo+dwD8yvdImZoiExEsKImQHReErqF3rbn7mrk0HKe2jweaCFrU8AwV
i6cvbe6Gsjj7ZAblco6I2sDtPSBoeyiih0yKN0qt7dSE2R6faKdveQHXARpygj70HP1icIADtp9O
AeeuaVqDYPmk3jxHqvIbCQNm4aSg7IDUvJUazskkORcGbePM+y+yX7N0mRMhHue7z8BdsI+Dw/1k
+EVMh7kCZwG3dImroQc1q4mab0spcjC8HmHnqVTIsnx10h0viNRL4x2d4toh1xGodiTucbs+6sC+
jH3H345QTs9GBQb5j1Bhtl9IaVwdoxr8fKHHNFC0sVLnkqtpNKGgS34sbac4Hrq+REzUAEAcdFbU
str1mLVjvOjoOG4zA7HBRij7iIIyKSXCNL2pW8brY4lqiuZCEclauBtwiSnIGaGlnSS1Sdy6dC8X
fAbDxLDN5V9hs98GzWvKXmsvlnMO0qYZfnfw7rLAzhafZA5oud69lzqaLHcZBDu+SVU713+GPKMf
4UxzN82Hjd08STSY5I0Kv2n3SkUiaycraR9UMRaPrqVO475kTgddqloKISf2eQTq7/59mnpwHRKS
CxX6OF8iaNDUfVANoIJk7ekODow8mMNYIWCSnnJjgJ6cxkcfhaapU+P9LB4XEQtlxEr+rmBo3Pdf
r/lL/EH7WZFmbm4jOcMseSUb2w+aR7NiSnx9D2jCFnzgUWraenZrrNhHTRm5SjAhRq37emutJ3fX
D60KbLHVl1FQeZ1IwNu0fR627XJDgHQ64jTJMylQ8YetWCXX0fsGO2jDVQgnNMUedVvwVOVBm6QH
XfuL9rPNGYO3zR2VCwZAgLnHEVGpkqQNZKG0bk1ZcOHJpnvJHtzNnM8HBO/zscJ3nRqgkG4YkFDS
0OnG62B6Wiygp30RxFG2hWjmqyf9897eekyLS0DuSBcTSzDoXylYM4XoKxwleBlGpMLIpdDK8s1/
6NxhYqoRAWKYGCxFeSnIl6VBNbH+n5gPdUNWfMqeVI5cYXIzS/RArfaGM/ivjU9wX+DwcsqR03V2
tU0V9AulFCe9uIX1hYjEl55d5/swCA1/y+tL4D1MxdGTaRk0u/OPNn23EeVzEI0fkhROtnagMmLC
7uhcybX789bAxlLDnuqc2Dc1T3IfElX7BU3UoVO+/5R1VrAi/Qnv5L0Udv6HhziCj/RmhnsQsdBx
Y+uFcAUCIT1b4vvYkpn2vzgTYn7S07J1pQOMyl13Hq7GVxR9uQNGhAxM7maPOpmw5+b54h10jmPj
rcSqB7n2p4iIT7ewWTd1LGi34oglG7QJeX4YXfnwiJ0/Wd5gC8VDIXQd65A1sXsDPcOLtSbVjdx2
W3Mac7mGsO0VOH+78za/yDDXgTzP9vbYaZfETc10rSkgGg+OFQnGR3nL8vM2P+C2JIvyKceylfEI
zkp5hXTOA26CZn/nL71lDRkh2Xm/J7eZGT9t1q6goL1Z89k1t1ZpZPfJBLvrmJcyT0aLITaeamM5
yhK35RYj/cjlP/r9rzfqk0+qHBV6Y9RaLCiHwz0kdwNPgwG4g61cZyJItR5vPq/VocDnQ6nt3ptL
nLn2f1F9AUAOjKUKOEXDK0TamkkyYjSRE8uXX67H/7HWymZSIU26VG6frl0WonzRDcBLWu7IyJUv
T4OYvnb+KOoGybhBP6/fChzMH0yJgTL+IuZcTnU8vE0Rpr1oDHlJuetxQqb9EB0vXsDsdbJYSyGR
zZ3a+Xpu4ZsVUf03b79pSvAxSZthLi8L2bheil+sYU7UmoCIA5VaFXTnVQgv/ZRe3gojkeXBB3KW
0s6P22B3CHPUmEn7XQICWAsGszMufubaxcnnk/bzRxGmpbg2025KKdGHyIteL8uwP15nOtg9e/+j
g7LWXpI/TMvWTYDbCxAA3diP2rd1kE9herJ6om9T0a/lbhH4k4WbotzEYBDTbRO4ZppB/tFGWEmo
2lixS/7naZ0ennUNejeOfxbSF8jAVsFdk0+ai4uzspvFklCY1IodpqlATE0+IHfmHd6BhMhivRj5
gxBJ66rQSM50MgUUk33Y7N9aHjhDW/Sw5+ctTkuc+JOz20mlyF5Zs5y43sj4vXqIe4kLKfhgB2dz
MBvl8Qvef/EvDfQ9eEUFHFnYHa5QBYygAYSv/pn/sP3Rye5BCNTjBHQZA2fWu8QN/mtRcpO4Xbd6
UJtq+VrKIBfyDK2ULXLeDA69Q1vrs5RI1P97UBsjMMsFksOFnubc4TR9yDTjWiz953+D2cMQkUXa
WuJEmRld/qvhFgJvQ02633IEIz0Ia2j3DZnkXpelmQzPCS9DOBajxqgLannGw3GyniTr9vfbxcGB
4hIeshvO5OFWMmMWwA3zn0x7oCM9WDui3gYGoY1KduKZJ8IIrLQY278AqJ9F7sefSyJK6hxDuv/2
0T71flLRXreIW8hHnskgOomNCTfN40fEkPYprLtLdSNuHBI69usfRAZ25x8Qs8WoU2hK4RvDVKVc
y4g9SUl9rOI38DE0hVwLEKsnJxpYksgzNkQ9te6MnL3MsGJDXIiWc45O3p6suBb0jiz/1+rUbbPw
EJLBXklF4YVqYl01KQaqg+c1JiPFUugT21t2ULmb7bIK4UGUKfnZ7U2bW2b5z6bb3rLLnmNYgkVR
kaqYAjjPVorlUuyPnJF1HDCARscB7/DZgV8TLEzKwObdkjgqORie1934gcLxLHHf07XnuczCNvng
EvRWQCUXt9OCl34hQd05OtRaIeCBVfsreZu/IQLaXP20zichjDKmhLmZhilo8LtIrPH9BN7FL8U/
p1oDRfJ66W13L/4xZfNL3K3hNk5O0+VQjRU5+9j+xmqubYkn3ep3GI2pZTN3dbqfraFWUYFEIdRw
fkp0ragsbrRqMLKaL407ksEaaMaLkgQQ329Jvf84kJvF6+EvcaLQqt7aax9lAeWVhPms46qRGQPd
CRHj2tHwexIHxjRJl4yoE3OXFwakYHLxfDRTuwlpYfGmW9d8ubQ1ZLZSHrEudxl1IFdCCZjn++M+
fLRh7KmTa625LbPVcaJBMpT9DY+lUXYKkFAFpoGQiJxugb6ClHt/SVOAzI2aeBopBR1y+86/ofEx
rhiYKfPKZjHMfmXn66fysO2g97OK6sRPtvqr04gpmNpTNt9rVgnAmnphb96K+uFbyxGPzKS17CzK
sfuoVUHXYeEcGGvv6ci74cQvUcRDPsCioy6n5pPr1nU/dfkmZoiqsqWlSZffqUXtvRBrSP36SUK+
5/JuIvjQwGw68r0p2ZOhrIQ9ujFE4LoC9/8z7nGgbzC7v0/gzYG4TVpgFYGgV4WA0YFKVrsNfoDk
c0iwrYJwA42WI4M+KU33Bk8SfkrzdCmEjDZilhtxhHpjZ4QHOyEb/bkKdMjjaZHazSm93d6rrRit
9YFEhm8MQGMKo4vT4B8gZNMRBKoGICjkodREIQ6B2loo2W1bKJDPVGdHlZ4j9p33W8oIQdJ23xrp
xD5XYDwbt9DqWdu9Xp1c8euZRzk/FWLn8cvMuKoDMUdLZzm6k0OkOXZ7ULvZfbkvaA49i501xOeO
nmSblleuBWFh47n+1MomfS5MvHL3+XnY9dqA52eVwN0SmgQ2/pIyQZ9eXafSl6hasC7hmE76W2x0
IzaEXA1z46SsQAJPRM2wNoYrgbMmTE6yo1v91NHG5xsKeYNUTdmnqLj643YkoJj0l/2wt8VU9gpS
RozLMtquevU6tatIsfpwqgEPhFNEqkG6/WNPLVbUjMYl0qY8D+EHF7E7VOb+9c6wGgkmXrrHvvQT
7S+/4OAa42hx/kh9bSTxoX6S2YAzKYTMzT+LWG8JORrfz0w68bQVkBVIP9GxrB7ZRTMR4i484cHO
XFJLWr8xlEl+EvtaD9yPTjWF60ILJKa8wlYPIoujwkXNowXp+t5+/FbZ1tOyCWIi1EJ6kWxYfArb
XOT213XPoW47zOgXWdgB2Vjms5Qmv1iEt4/B/Om9w1FNhRnT9W3R+qs6JxXaJZESxOGX7tvpmAja
XRxQJHPhtJNYPbk7BbJ1hpVxFo/RFPiFDa28UtmKMmbvNhBas9+zd+46XL+FW/u7EHH/1u4gfmpl
56jj7erhBVa4Fb4b5uxgWFj5vgrXI/srhi3y3t0X7wFlNy49qWCRCSfHUW3aVHRp8WA+zh2bYKQF
K7JhexjhSZHgHICN+Viw/Boz7dnL5stecMHNxeUfCayYQR95fIrHK+RHvpoADdnS2Qb/x2ncpB8h
IXeOUoIQgRgPbOOH6/U3QRSlXa1MtVimE5cssegRWfuUCOo5IRPxNjIESVkl6IGVSU/JgF7FQRm6
6fjhF9redM2StGMNpVidGd3oVBldW1gMszALBDxaKJWp0k8o9QBKfdkoqWZnMl3+AA9NEq3tWivw
THa5qajE0pyd+XMgOnsFejP+LAJI4wQiUmeeV2tzFE6CTe59fik9KrAh0ub+v120OMI7w9XfcDW4
TEn79qvcmAXnrLwH9TyHuEQ9ky/qpdwl+ThLMLlxzSNsptiA5IZydB0qD11gn/DBa3XGyAnDJVyE
185tYpTwqYrbDoi+btufoP+38YyYe+y/goooKjrwaGhLQxFoRGMr8W0ikvdXdwOfWJYQO/JeOCKB
oMJUJpXTh5faDAHjU0aDImo9+MfIVH5yghWQtDHteNTdhZPMkk+f4DL5MkxAslqiNDoN1mqffD8A
OibNdsoC/0HjBFhhUcVtt8IWt/t+rv1PYOtcRGXrcCD06LgAFp8L8M5nWE1AFWpvsxNe4pN9jBXz
VHjnpKkG7QeRK3sx82WRmego203lyCeu24Q+r/hGBo/kWtxzAb7anuqu6WcRk3x1zXEewCvQJTU/
XGF/5jvy/sjpFTP4LPciONJwUZaL8xvbcfKJDcmdBekFlTAm+2D1SfCz/yToj6rGldN8+vk+89QQ
ZQDOzukeKmT0OWbtmzT7hZdlQ8z/r9VZg8qxJf1QkDM3gORNfY3iF5sthzLoEzytlkapPm2QAfGI
/Zw7UYPIOcQxWWnv2Okso4fuDcF1OU3ZLxuPNToshV2MiX4rKSehLt8KhasCbSE6mnFIB87l4DWh
ewUXpvXqzlbZE24/SfpbWUNqKOMKd+fjE7D28IRWlytIq58mL8F3/6IIm4+dlXPhm/Vr4mAC7eWT
GpCVAmCTCdCyI0L0CQ7gffkqQew9PyDpOAN0DbBsJLVY4OOqWOCsikP9q8sgpMsPMB0+IM4t2+ww
Ke0xuCOgmxxZfjY8UHkWsOlWN4pvUedyR5TxqM6GR0OZ5VA5Uv4Lky2DgqpX6VaOKdwmF3lcW0Sg
2nblPEMcgKJ7/+bDBMYDF4FtgSVr9sjKlNJiGLGl69gBb1LJr71r+BOOqrwA44iuNQB2xgV3oYZP
i0UkjK3FsGSOInb8Zm3t8kEPk4PqGk4jF9d6RnxuA/OH4P6ZMSr5R7Vy8HMF6LOLMzktH6Df6nyq
vtEAi7dSdArqi+gFCxf5qUu1UZ+Z2FjNoO2oVRRIonP7Hr7YzeVYwJm3qEIK8gdc8/ZTO6PrCLty
VsMqYzdi/a7jNY4dZ8LrrIk3OVhzZax4UDBiMhGdDICvZTuIN+emsjsP2KnrKhhyTrmpbY87AnXR
pIS8lDdm5ht4OPzjeSFVZ815dPgP8+xx0n4QaIvZSxCe9AQvP2YQRTr6kzNpa2BtiJIMOFeLbXc+
46qDzmMgqbyTpibXW7E3d7/GpWomoE6hIhP2gSZMaAO5nxOBE3s0BnVRBWkDCcDm4M9ceFktvXsr
/9Ko8BBO/CDAu7FPves2k6rFiGndj7/fQn/7nDg10mPQsTXFW/t2V3TvHxqU8rwE8JmqYJ9DywI5
oJqVqG5udZGiZUvnI0VCgEO33J2i/2/JARnRgTQzSoq5cyIh3VLkkjdnn2k5/aNcXDdDLxjLNPpk
AMZjZPpwt9VU+dKdXrd0wKgUXIL7OikJbBS+voR5SZ/12od6bOsSUA1LxIzMp2wuFvBFAM8zT+IV
UOzZexkTvAggZScE0o+0GIJ6vVyggS2XFYx5XLBy3Fpm1tP33uQrE8tAKormaRq0vCDUM2f08UIN
hdWkIgYIKECO9/OAUl5LZg+CJHaEKIy8QmeC3Hc7kbKLhuFOHgvn3jjMmh4MQWeptADlpXYdPFoU
csw0NBzxr2GRAi6htY3pm6xH3N08v49flJUBt7bcxq+74OO+HC6af5XQM6q8bbfA1MKzI9pgTvAk
L2nXj6IaWKNPiprA4aWMGtpnvsPH6s6HKtLo8W5xUutbdyXlieF61b56Hr/o5ge1oaPBIWk/0QKt
LL9s2lyxwKSIVsMOe5FPNmZNZlmAJXRDcH5U4IwudVBzQ7EAENA/WCQOdxYLCS9FGdiM2DMb2OPy
oW5QwpNczfYv2B5aPCJopLYibmBRQkxxsKHPSlhOrU4z8qDVAqhTZztPwNqfuZNB9F170SGlXfKs
YZI3gT10ftK+223WymPg3DUyto/n5oyV0hO9FrUGcLVy4eMZBlhKxqnvP7OE2RVKFDh7rXs0/khJ
ogztTxOvhX4eBwH2r/CR7esyZ1dnRrPnzLoWWUqAGk/Zg5JludtMHUiZVkixrowj8QSNv5eqkA1K
NVHiXL8rxw+LG/NSKuqYhWxZMe5GxpVj3zIE4IPdixJV3lu8kY6CGVYBATy6T6YXR02mjNy5FXG1
2Fl4nNPuD2E/EIJM21+478QCvRpiRJDwPQTWdnSY4zlz0aVFj9T3cRVS+X8R1DmXGummBMqQ/th1
0xQvVV1UXtnlU9LWRjGiahL7Ey/eVQBCdURhEK1SBn2tgkbS6dGBCvAp4Uz/EvW4+/uPnLeXbeUK
Z3gkgFTPAA476lEUJEC0VFqxy5GMymQqfeOd6hYgjr7wx3UR5Rh3HbBLMs8612Buhim1xgTls4d5
yidGG2l7m2ZQ9wTCAQFeOKW61s/F0SPXZ/2rxJbtrhr0QK5t4lBHYNMap8uVV3I94nSomrxO+FTO
NaVf0U0F6f4srvzAGaHbvyVWgY2eDPZj+CknHPqJdr5BogH8KccNRiooHK15Eh99OVyos3sW9SbM
M7dF6akFpp0e3hrzszIP5T13qJdHnEJvb911oYjqK91rstOp+mVFAyoiiBxTkg2LuQUkWf7xs7sv
e4vvA5vLDwvZMikvUY303LbyAdF6DvTQj1CNJ1b5LuMjgett4q2YqFV63Fp+vrLo94KCqL1h6RTK
H7HciRJrC9FO+JvIveYTjUj5O18mR8dDif0kK2/48lsdJXSc7CqonWM+bRZ7xwk9RCNHkuWm8aED
ckUybMbK/+u6BS8Rde3wDidP2zBZczotW0l/HDigpvGoJ6EXhB2sQQmZY1n9RHAQtVnPlIKkHSwW
ejyR789IbfISGhhuHxHrCrtUTywJmwDfM5cJBPmEmwsVv9aJET6Ns9jzfLOddLDpKwuCcGGhiL69
GwfHdmiBM53tuqssRJaAZMJ6eMTsIQcelym9UEcPH5RvDzxSe79jrHEPhy0xk+UbaBhCGE+j1XuH
nPvmWtTRv5M8NHeeeNXkp4T/QSU7WjWK1zh8MZ6GqwmV0GJKrn457+fdm0WQaUzi+Bd9IiE5Aq3e
VYoy2jDHppxV5W1BPf8aA0NcoGUBym7DUaa2Ma5Tpy5gbWn+q2V3EcYudyD1ncvjZFfRPSc4loZI
Fu9+38glapbdw1RyDqYg2OjYp0Z+VBcG5qdmDZ0amEbZLIcTGVsVRYMrKhqKlIGCIbaz82xf5NBA
sVEnnn2gXg7sL/TY0hQadc86Jdt/2B9ffJ2LIMUVPld7cYKNLG7ZjMIHwTMMN1i4WiMETSKNFoDz
newpaqyMSg9Xs6yceyrRCo9h+Zihaf4hiG9wVJpRxFoK18Y3lACLUvBp8uTWl4gG51vcYX8R6saT
9nJytGmrsxwdA/YeFmqUwKRNr2Lwso5EqUzdm4vJeIECQoKadGzDZw4w5ru6LLFUQbSPMSWOm1hX
9aV6sy+vc6FSrnVhf28PReMkoUBWysvRpEaRW5/DuraaKrPmfuS2WnVhS2wGqtL5sJ4ZpI7mGBAt
io6RIU4+B7VPghDz6M/O3766sSx2F77PUWOqAJMuikiz7dIbQpR9NcLdmOkWrOFQ4XOF8r+6Yk40
rrs6edWeKb881njbhFApuqUQWt0bKePG93OzG4UhVX6Z+fcQq6jvzKAq6/HwkmIqGqroTZikiC8P
aitjDqwDU/Hz4T3obqQV8wU5YZlC2FOEa+nYoH5F2V/atX+1ZyGggEgrLMIzOFJmSqqXs+5hvMaD
sNiArzi8yrTb/TZqL2+sfPXxdiHkxqTMIg+PSjslerIY3QyluGuQGKepIaluqtj78ver9ajozBCu
CS15AoOQR1/FkwWhX1d4r2OAoXQ//y6T9PbFU6bp5BdNcM+tNe9XjyCDu/S1tlWOQ1BA8X7vvoSB
e9t4epv/cloQjoH7seYDCAPmbooDO+Of+iQALlNsVzj/chcylnixRh4OIZGhKUbvX0phRU/E8m56
KkcHwC2Ub1T9Ix/phWCgl4wl5yyTRZdUOvHZv1klSNL9SIUEfpzr6ft9TzaAxJsHjnntfUQ77R4C
OHAaEl96bXHhlTznZjiVtwRoryjc6XChyU2eV66Mi21sqrYcPXDREsndrUVG8IHpHnWcdSM4n3GY
NobB96bQ1/8MypikVA78gj8y/YhV4oXEfLj5ujhCMtolIxMhZIyWO/fvjEm/UrH+6o+ZJtVZC0Y4
p2BJs4USr+sAXdWXGJv62lum36FT3OC5l8DNjKrizrT1IBcCPXstcpM2xWM//rNToWDQJsuJfFBr
a5F1oajlaG1BPuOHnDnyBuZVTQ7SKeOP/iv6AnnhgId0WWrN/VcTSAPCH7lUUxA8Agb5Q06ByA30
SolB1XUqX7RK/1SpeSGFrOaU8t0IdVte0GRaHkK6ltaKMR6hnu7QFHEpDsSQQZPEI0L6DObHb7p4
gOXoRq+7B1v1hMtBPXdVs1xaz0NVbVBeMKTVbcD+cwpxzv6u5Csi3y3TFUoS9mesFvnPLBMKeb9l
S4L3oumrVHHLfPHxMuZ/vXP4w3BpnA/faDPTtsS+J1wh/5stiBTYst1FBnuVwMSA765/j7Ejdc80
rBZ6pdDdsDc+DfPf93XY1kfZyGcd/cQrOar4FsNyMclMa3FGCoLTKTX/RXtr6dPsw7kP+fe1XTGh
bR8sR6ONNo1Cul49GheLDIyPqlifRxuqVAxKQ9kkD75PVvsybjD+yocobG+BJbuLg1yNV0QBWEP1
WML9v6CkQoh4DIiqK4HZurMFjNGhGY1cfN6NszlIMKDaPl+yC52Rm/pMEUfe/QgUr6KsaDT1YB3p
BmHiexw35tlhsFNWM2VrmQeBM6LARGU9ZK2H+kawpSLQJ6xXjYyYSOenvL4Dzh8WX2tDJTA6K02a
5ynrNYvWNXuHJcfh+cddbYClZewKzr7YB9l1faXHtCKfwPJ13XocfTSaH8gd2Nmpq3asDGtYfch9
zdxdUuyfwzGmSdtJIFWsmsFj1YoudN/shl3ApwhMsD4Q07kE4GNhAHpBXWGPvc4+m4TxiwycTZAe
3Y4cRIIQ9TkJa1HAfOLtaG0w8S/NrpiQkPFp3fbDm/Aw717L40YyOGKzdeywr4t+jHvZUN9V+ZUK
5VsapWJlDHJifif1K00/iRw0006OfFQJJzCTubX/WW/sY1QsY2QTG+pZ7jLOiiA2Q+7MRVjgMZDa
sRdRbwhaNpO2KyrqCucHASnOBrxmzrET4MTQ0uJ9k/V5Cdj5LwGYq9fwqhP2qQTlwjW2ZqOvyLNC
Ua360B6YJW0qNlZwA4Vj4Squ3QxKW6V1FnJIcd58btZ6I9mj6JLYTXjfijwPE9G5iYlUGorNsvfN
qiSenx7s+o9Ofo9KuYbCexaXwk5fBeAVZWaYQ0dvfKFGwnlFEkJee4fXujyHOyc500YZVDMOiZIi
zrsNUfMxqpszKE0RzTp3Yw+qIwUSPkRqPCxZ/X7KqtHcplq3pnUtmmcwAPljOrbfeJt3NoPGBOyY
iSm+zDRY215aPUsJtEgSY2Q5r8i4voH+4Qo7tdREu+Nz7qc+zY8iK+a7uXvvLzQ/cwswZTV4uY+E
EFZDTh3RWK1FNDrcaxeyBmAUTr3u9Tam5Q6C9u9mE0X0ycZo3rV827yLZ8yjN29biK/Ezv7OWngN
6fc14MTy9Ti4kWERWiKqZJJbTRI+MZ5Z/d3b8dQkEEW5zNbhHckOtCTq1+F0jR4MPtg9ETPIhxam
EhBqkav5Vo5yg7LsqGEr6aBaWNsaOevU02mJYumEylok21KZ9S0GCKLhcUlZXBwDZC6XR64joG31
IGfeXEF5Oz5W/iapteDH/toE/FY8rc7q1r98P442CjufVrcm0NadXt/XF2MPhI15yBJ/hBqzvIr/
jRGsiwgKFLvvZ6ym3tUqlA/feuGnjJunwN5zOkjI7VRhCqOHHle3ed/AjqVHBfwPuiGRRAnAaz0Z
LnlmYMFRK9Nh9C+gouf+tVZ8Okng1fYyw5NeAblroC9hTpaKi14h5YdOmg3LJ7nATBEPZJFxuFRd
JmnFIZoOVOQbNOoWjaMka06cdrt547h6ncoGnzqPNkun9vdJjeVCCCmt1B/zI43N93CsE58nFb5U
/3IN5kEirWBGlHsQMmh3QxbT5Rljp5sMxqhZKiYCNhbWUOvQd7QzAnvHcZ8EaTyASt6fhq4bIbd+
un+mp5NeqkftNM6wGHhw3K9yCgddhiB5DnxJ1DXfMB9YgcZUN48oC3lFfXKsGxKdhFVnFFdahC7X
KSe97LJJ/p6gZ72BkRO8ajT9TBfgwcmpStjrqyXjZRhdbszObtRlWY9+BMlimVDNQB5akGl0DbAZ
1dVPXBylW/AxbnL91azF0AlAZG6nxBorlGncIpBUtY+YGKTGhXfnG60p/aKIdYWluXpLSuUDywH7
IqLKV+l/NnewIDe+nZDqtYFdmJCgMZYNXAnp7/OAseWB8bOb1XTb9m4TDWuhKUcvFg6ezLxmP0Oz
B9D8ZQjWidCUw2oLoRp11sWiLHXPFqHQWDUMnjc3SB0PmrFKc1tiDIKqcB1P9oT6Nmoidv57yreU
fnlVC39uF17Psvlq4ichp95TSIyAgdmqV5HkFbFM0pPlPD9ASBxOlFnas5dIFD99dBmDVFJXvWuM
gTHF4/7ZKVRVRCVsxNaQRkRulWrdu1WSO14VVzT0YRg5HsM10ix4pI9Hqhv0ES12sQF+fCMEtF+8
nO2PsHQ3eY71u4/eKDptnZb0MRe9uZr33H669xmVF05a0WCGxl9VsI9FwTmZp9PRqVYqlW6sNaik
KPoAy3f9PBWP+0g8Jk4AQHfekR6WXz3Kt3GMUGW2AMHqu/5Vbid6zj+OifTfsVuVH2BRGWTpx4wn
WieG5+ddMtDdS17xvwf+Xd6a1x8eS/aLfPseCfOVuZ+ASKkMk+m7UKUnGXqPck6WIkBMcyt2CQAJ
ldjFgtg47poHiq0Kttf6d7pB+Esf8YyGhez2peWqrnVTVG4QOCdBDVHY+5MNyyEmr9Far3NEptQY
zxdhB30LWI6dS0Yrkc6Jft6DL19iO3NHa6W8wFelgp9C1509E4xsqyyB5ekjBpJV3/wKLZEyKXwh
7/+cPpnFDOJQ8bc0x3QBO/1ELqiX0+eNQZl7jstOexuRT2EyjlyJYD6T2L6lrmhkEcerc7T3Z8Sh
HyS4sh1ESgNc+vUXea6N9kN5rV2HHnzmc4uph6+eaNK6xOIi4hdVufdUs9Xf9LUh8Mg2zqzVWa7+
eDWH9ht1NkhRj2IX1w04Gm0ux6+V43oCZkYVleyxZS2T6PL6HYbm/p4El3ifiVlzIslomNqgjxDo
/LCiatAxfpdeieHutQ8kkj8GDh6zSZOQBBYwjDmnnwbNGJnyLJnkCxyqfYlMEmPtU9JVWVCHlmY4
SUPpsF33PZUC1GLb750gGKfYVG1xfdm8XDGf5r/3MYHav+SFBp2p26tetIxmLHu7yBxBei94Vgjm
tv9WFqPUJKFgGJmuFVBk0SgSDbkr/J1N9A4qwis7knyj/pNUFb8OjeA1zbSVY/Kd8AgFdDGXesJX
DxIUXuDzJzUOx9s0Z+/xtghfHsKM2AhJXS44NBLQZteELDOjgFzg0nFHispn6NckUmztL0WkzF8f
kiHyD5Ln00KtLjchtblFlmZ4ZOQImVSYKdQAXmLb7r2UnXbg2nzdfXdExo5qEhiew7x+qh1DcCkN
MkWRu14ku9l2BOMFoZSNW9rE7D7f3yIdJdxb+objtFN6hyMYCGrf8pJZBmlXKDKEOzXWpRCQr1Lr
6FlfV5DKboi1+T+AUfYgP+XTGCQqaYG1mnA6tzN2s6KFgB2naPTZOEVPL+xyqVospJOGDpE/YImM
F0dcIxqrLa1dWcfM8N1n13pqNT7oL4I8uVqZO+WCh5oRGqLPHCghV5L6+HSzdmgUyNmK/pUccBaJ
fIfHkuvcNIhr6DLs2P4ebktrVkwXXbi08Zg2BxWlUf+ve2fNpqLVkV4hJFYseqFSudKGthv0QjZg
MTUqoI6xKe4qU5BWQVzPF3PHcslsc2uNejh2lA8fze1A67MFEHVSP2GTMF687JM+Szy4eTSJTFYd
oXb7fwDF/4cYk4Y+7kIsgeD3kOmpJ/5eRXQGEE3DNN3yaJRN7v1Wh5KwHn9Gj6ch9lfYiuSKADmk
yXExRfrLDHMDMA3GoCGJfaTgGpwmGMZC5ImkKtfqLR17D5ijoi4V5yB6V0E5mqeS/7MeM0FBDVXe
K4nYtv+NTYjfWqNLTBFZocnZqsgJ5bS/B+hhbPbsTH9gct1a3KQLKRtrDZMWSQLYwAquhLZ6rAVx
l46N2CaqyLnvlXacCeSAodmEBmyG9qIbDUt53aH3JvAWzP9UOE4D3SFVigO0QCMMlgpD4mXF2ycj
3+SktcPobdPevL00q/UDPCRPSL59xUAGz06fPoRerTUVE6gUMYc7MSknP6s5d3386jXxtqmF1OVE
j+pFHpPcFma/X9NTadyYqF7M49ogJWufU5Ne6EOXDiq8DTs+ojMyuv55qVJN5UKquZgeh0VcuHgi
2YDBFjrQuaoSFOrIwfLOsTLn5KSJCvEQNzs6BaTCJQqFi9gp7tmMTt+QVx4qH9HeMMhVd/lTqNuy
jFILd9b/FQVG3PiJlLdxdJatWBR1N16TTb99q9736t90ZWGHBsNCRlsXk+/4ZGj/uGg8BQdp736c
Hup7t9N68iuSCL26mvOhwXNrWFjybTGccBjXb6Jc2EK8dkG0DpPtB0oCKhMKx55CBcWFwBVd7AbI
GL6+ovZxCeErYWGtQTajCeT1HkVfBmeRG3xvHr3ZIYZmW5AvOJXSEJThhmU+E+ZANqmVhooGfku+
UUBWzy3B9llCLDHBMZd1iURA9o6h2c9RHE1XbeoU62zeUcEBjosxAVd7NJqj2BNsSoBbvaB5XH9O
OpNC1x9ka5HwJu4oUUXcs8jwKRwE5uCO0Sr3XHR1IHmdkTWmraOUs0bcQ5k7GQs44CzjeUk9ONlX
Kw7EGd0jVEXiwAj3aVgQb3tQT/9n9mNvsdELoWm/0XCxxycWcUncjn83IfXvS6G5uzxVeZOlP8HM
aOpF9sNc4w4SYEJebdoto43KeqO4WSz+qx19DPsBSW8ho23ZQ6akpyLu8lULnuGjTUNaxIlrVG+s
5gd6EO6afIxrYAa4NPtirDQC6MKmtTSnnjVGIxNvuWqZ6WA336WYEpqtXmw9oe/eXxmPVT55ZPKX
v9GzTaBNFj1ZJ3SwRStdm7k2pClkAB9UsS9hPkzwvrd/PIavE2PuCZTI103SpFO6k8v1vzYKAGsn
IMxkySOQd066wxON7DL815Y8JukouF0M3e+yIScJa4KxTAJpaIp6JjLmAlOmQYAN62R/n9YUeXhf
DZTsfRKYs4F3M9KTzuBaSuX3gsFaRwtqKDqxiL0GHWfWjNZfBw94atutKSIavwGyMGjQn1w18PDb
UAPzR/sRBpmIbhVK1X4JghqTS9zSg4pBmXp+R9JdGC3sUw4uitLSBXRBDMNHGjrC1M8xzn5kuDTS
+ibNzwhbdtyIomtkSPCX7uo0SDsP/IPhP71Rz6UDmONsnrlK7HOMVh+qR8vPbp8+PyV7W/YwfLbJ
1HNu3oGz9KpomIfDBLHjiHAhLe1L0xdw+S5/KCYBvOlmqXLxlLjzCFYVlFig49ZsJXgiEU+EiUcd
ySIE0tKNaWHD4jPcxlnwi6CY6+dkHmX1VHmklkd9BHHaibGO/Q1kN59OiMdCeU5ocGozoG2TY6vB
vN+DjmMD/YqD1Q0bx2ab8XtUAPjwC015OTnMJqGp1+Lxl+oxh2DjPu4BWcqhN8ZszmwFaU3M55ef
LYFEvTXVr+fV/kF8QeXonCXknOxIK4HK8MYXbFQ1Su2aCiJu6DKgDRG6/30oHgflcc5akmOEXQHS
7J7lx3rgbwv4MdXX7q8HzWEi7kHhYq+hGsCUdOvorm1Hla3rpz+yKkcFzx2WVuEi+xtnMO0v0GH9
87S+nV8h8xXzZLFp4xJSnOzvievlvEag2s8KnJCstxCHSU6pwk20yB8GQ3nJXbD8zd2fOU7Rw0Ee
W4CM+BgFNHpZbtgmd0GhhLuRFbH5dWlfNeTEumOgEoLADFHP6/oQduB6ZzT2QHWjU+akCyymmJJI
utwUpE089UjnU4HzKmnGdSnp1n7jGQ24+bMIF+MknGFivarwrVkDrw/8diuSRdgmn/YSRL94sUE5
iGR7VOFG1RMV+Sv8RIRNaKXXg7rcPnjRywz540pwFlhouTKRPHaSBa1fWffB21Zu7dbhIBsw4bOI
jh8eJO3smUpvtOOhnnb7p8pw9/Clnkll7Z2ZQtiggoyMDe/u+hB+T9QrSYYAU60BlUM0BPopr3/h
lXr18wfpDeC/BT2CNtuCowrsnMw39Z8ESeYIHu021TiZ87V+zd4NCwOSdndWfO1ISvSldWqOFu6M
aFN3hwVJW+37wyIBuzhWYjbCkd4rQlqkdLM44iecU90KJOyqpMTZ4ld+/d3E+Oh/qxSpF+8SPG3O
KGNR1BZGjtzwhLrPg065iRu8G17JhnlWSbqqrE9FBrM1iyREA5YoPNSF5Fmh3MYwifkMgKlSRCGG
1tIUqa8ePOZngDlJHx+8QdOWByYLcwo7fQLmlEJC1UZ5FtbY0wEJXRz635o83GpwTDuzvQ8GnBJg
R+0uTdeYs0ACXfZgwo8x5cCcUUXt/9flpO7S0fI9pkmUZkfDcYUGYJdDxSXvnQwwkdPRzhUxDE6o
YML7Kho+5yswG7wXhN30FEZqVPaTuLwkMmLMYZXdvazvoATTPX6f5D3deD5eDA1haibv0k8Et7Hp
1FHArWdVmL3sBspQDQDjBERfihrTWnry5LaMVIQYap+bGf0twFBA7aJcAqNLTeFEWLL9VKExOFIf
prO07T0eVLjWgn1pUIRDYlf/AoIp5Lu7VGqhECRA4OLVs11zgdliz3fU4nvO0xZUSpALBU+MoK8g
7dBj9/Hja3DN0I25bczoV8pMOFiXpiWEj8271OZ0NqM1QiaGGtgztiG4A9lVCkzCQNr+tMXzZWWP
fSqYC1bexVhrO956XgtEO17w+H5zjVWKMyBl9F+ZIDIkPxI+8C0R/loDErOZf/y6ExHV8ibwAEc0
W748uFT3z6L0OmasPYw9gSVoNTr5ExuuH7TunSBxoufTre+QEeNjE2oNJfAYpJD0yXIPRXgrEe8U
sOAvRubUhQTCv8WqFz/JFL6J6+imedYR9OGyr7ZhmqUqpp5CgZkKu6cEYIxRsI7dCCWHH5kzfLpg
r4D3lSlNUoWhPk17IpItdhnobCNgOnK4rPWTvX/nN18qgyUGRpq+j5EHHcLPoXzaISZROBeS34kb
bz96J8ULy93i0GBOnObUNYWRsBwT9MQ5XKexHXcliG6QBcRbjlVmmdgfwLH/v6Ikz01IQIuZoMLP
skTHsejvTH+X4Vd+yqFxIWyqExP/ZCcJxsTiFkhsgX/ykqKa6RdMmKvdDROQKBxbnZLp9NgcWHxk
gpd/Jnmp+5rhOcI9zLZP82qlXI0/uP2O+5md/RY9dZZp7X35v4GHpxrv2W7ZMVh7w79liMkwNpTD
4MBCLAktk2cV+siiciCy7r7H6GcZ6V5BSd68jDCTniFE86jhA6OSiWfoxu+ZNFuXmC2RRqCeQJ/J
2dowzDgne9DSuIEOWUd7Bl+Tz1ssINUS+5ivviuTMbzn3/kJMYfrPsioHXpHRv3ERI0ovqiXc5lQ
UjJVxkxKDfUkq9BqZpL31z+v4E1rKguKzmFXbVyHVTepe2HQrxIdL0UEPKmt535k+lDyFGkq/Klh
utO+3/lPoQRsUZOKNgkN0ye4/soBs7lgSj1HOe6whgM5lFIDk+QvDtAhz+zzCMhfmgqZU4AP1QgO
C2Ui10RSs+hUNE+K1E5dAC/a4xvuqYcoAeHFCCVQ5IqKJjt29irc2dkTVjl7+isHj9e/AdXd98c3
sczoR0Z8xOK0O+hMqnyeJKKMPoFkGSTvpTxaqH4dAEPk85dRNASfqQp77bHOCcPC5gW47BPZTbJ5
wxaBewEFzoY4d/oTJ+NLXCBAD5slnG4q/e9JkIbtcqI3iNM1Tux7Xw2x50ahWNQwhif7j4gfupse
Z1ISUKz513E1l0whCSxMY7rORHuRJhSSk5O6NcvlIlUtkMlEps1mPB96ByhQKtP+w0f8VlACtv2T
CSXDEsVXFXbjtpgJSBsTKmDndgmzru7COmwIghgwXdnTmY0luK1zw6+HYdp1hm5/SXiMwcRnN6MO
g0lajcGquRBiawMAAF6cKqYmtKrfAfe9xaVFafn6d2nfp2ev/vM6EVH79izS5f4nZ6nJICkU8nSI
q12qk4H5e+CRCgUMwKHA9sAEGvFXORVJ4HNp/jXo51ohVdfAa8BPtlm2qBERPkgfrZSOV1SiPz8E
pj8cZQPVImsPqHND640a3lBKxOGI8nIul99f+mjD2UrZaWweoai6hLJPF6DfNTLSp/90V4i+LyO8
w6t5AuceYRbw4FE4kuOdTC8Qk06y5BHecF3WzHnTN4Shvr1zSj1xHfeSwY0SEcrB2wke9NijqeyO
/EGl7HYr/IxoFqVuCXFhRyOx1hwFSChrBu8DWsFShkMDH0t/aHHUDIw8jOmginsnCquAmeVs55z1
cg6338JqyjMZp1YSmNxrMxKGH2PyR5vSQ1HXZWNMLN2UZWyVmLb5gEd/kKPQaVgtYlfPyvqrW83p
a9DHXOjWZ4cJZvfonQHGF4edWtOmkxZWgsaBmwoFqQgIPDt5YoGSZd1ukFy2+esDhSBmBh5HXIjx
4UAdT+kDBRu2y1HGGIdRugwODraFSQTAro5RGMWImb2j9hc3EvRYl8d2B0t4YPl2lE82GWSZ/ega
/81A57gr6A0giOe1Ak1zlVXyEudFdeM4RuiGxRkL7pPKS5KJaNk75KvUhCXpjN09c+dPLKpBTCrE
Vjn0MgFM5nmW4Lmi7/AE1HxjHrZfUu0MidUXyJ7uavJuIRqmL1vaGxVY3oTKn7b4zFU9JNqYld9e
LSLSiTI5VyL10EYbEtDNXcuAHDDvtJifKKbThgaGQzxpwVo0QYNPxbYbvDEo/Q6J6NH7yO5mI9J1
y1xeWxlilpxrl8M1O1JqP/2DBKIqqiYDBFPIHjk3JO45lqEL0fnlh3EQzCJxmYexdt4TR2uT1vzr
3NmlhH6FfWGWuy9wBANiDMlB3fk2kbOOnIUfTrQQcT1rZLlDDIHJ+LgmYh0/oei4O/qgINJVuHw3
Vy3SOY8p6YWlsEu+WYqNFekhS4t4Sw3gnuLKsla04HC6VvHc+vzDPb0UAiL0o0cGA1SXLXp+0BKd
NXihiDQjXQ9UsVETXCvT201R9s9MOOXs3lYWYFnOYLvi0/5LuaQb791FQDEBsP9sAGLjbSkKk1yA
6Jj/L6p3eAUb/2EIJrvXv44Fzh9c4/5hTvhHrg4NlgngHKjh16RyUq2KODWVJh6WImrU2NrLEwul
NFeLALQ8eepqBfvDwD/SzvkLNlL3oHmnDeL/tYsfIGiFfjSXSugHVgf2pl5/orGszQ2YSKO/55GB
+4EPNZp09kBHsVoBzgdf9E5rkpmWZMV+dYvH2L5qd9jakQO6x4sjkuVZ8ZEpAxhbER5Z2rTw7tYU
8pd3vjbQsv2c2AxXgZxaSODr+9+AcPnLuauAka9R8dyRGwi0Zq8HpgAXy5jkZtBbKyy2BvFdZsnH
+ZqUDY1H+JtWVtbAejFBgjDnXwdPeJiDipyD+rHxlMOIsf15XtBh8e1qRjSoRvLgAeegBfilU4Z3
+CJPaG1tMOGkn7MfYW3FzsssklmJFBtk4guAjVkwapV+IGPG+dchMQRfsR3zr5i3153Nnde/ZFzD
H9Vx3SBU6v08yGI2VAp0I3HfrkFCBj/cG2VlSh0VuRVMnNTZzCV5/uPu1KpxnlpfXEy07UxZGJNP
3HJQwgb+iEdhnGsSiL6jvNRyZyQx5grCk+j5WZI7bhuSJjKzEV20KIKQkzFbBokFZxyl8ccwxehl
oicfv9DuQzQZoW0OsZsa8G6FPktl6vMpu4LkDnwdLO/fpyn4xCaodq+XK2wJpUs9NgQfmL7II6nd
d5toh4TNB86KhkwGv3XATfWVW9u173Hfkj80JoAgx6xmkjBKfc9aP3/KJqU2Utpj4DT2LtWGYrW2
CzBEz4SSwT12W1tMl/aihZ6OQjO5MOu6WY81Jx/EwSjCGTGk9EDl+GpJ68tIp2mpplPGK2NHZSQu
xgwVRZ7llPI8QPY1+Iu53lhz1bdmzhA0kx0kgJWqjhXlkT7VNAwXAQsjYvFWF5xpYb5C0URnKJi0
OyHHFliNe4so5aguta5r3ct0fKyI//dW18QhcyTJUjprdEndRSMfgO3OZxsZXMdgiFJZK3aYL6nV
DgCFKYH/aVTbGNUvDE6Ze3DLEZ1x3DWCABCdhCNSeqwKZGHlQ7anK7/7Jlb1yuO/HnUtNK54qTro
WFrDN2aIwzqCdLSdOQLdHtOy/bu+VHmz1MxKA5JGpHSy/G6y7q5i5mqI8FIfVuHBLxgyQrSSc0tL
WMMddzcaMChfTtuLa/XQkW1Qskt0SWAM8R00pSTrC2i/lC0JzIFOe1S+VxLqcj9aHg3LZK5qKMNn
3SzQMZ7ryX6EdAM4ZcacerP2aRTIdp2mviNZhMDFC3dPhAMg/gGqykpmEVdO1LyX0Ry7OjHgZ0zw
AUQDvD8PctA8dxYfk0dC93JTsh3DdM0VPzweM0xcjkBsvBXPr08H464SFhn7WU8gUzNQ4F3Nw0W3
Jk3ImFmdOdmM/5TQVXuKL6I8sINVr9i5dBxsNtLdbWBdT+DZBRhWeChBS2kiifQq5ecEHpBbMCsU
Y68qBO+ApH2vpa3VSW7PPjLuuhf9hzEqGW4G9ct45L32fZVoyhDPIHI/0JqG1v5tlB4P11I6ooUV
REiOKGsb3fJU0xZDMdS3OcuurHHBNITjjOUi1NqD+RaV1MbNXPpHN/wUH7ECVkkhTWxQKLb0UHz9
0icqwlRak4zvB03WmUZzAO9tBTPvgw2sohwYUQoZEVidY/GOsHklkE+SbEMYO64b48x+akcFbzYt
ey1zJXpnVsemKH3M878k3GFwzVOtgNcjZQ1ljXKl7VElvGzbw2Od/Fy1EX3mGfiC615VSAAgvAoM
JQrO8RnahweQP1dgrRtfbM+O6ehA7QRO6Z4qcsOVQxm6lKSSH/7FpH0clUpkHB7US2iGU8F5SGr3
ZqMqvEaCgNdK1JWq4LQLfzOYXuHtCPYz86oPO6/xgRgPXmm58DkomntOtl1OBf3G9jg4XV9MpwL7
vldONgTbMrCorSPWUTq5iBA1Q3oVqf+tPQ69pnF7ezX8ju7XUSJOqpUYQFyGOzFHvLE4Vr+x6MpD
Y9MRB1FkGl/ejv8XlfbYARy2B+r4VfBC+ZsIVpxqljKI7vKaLSX9if03SZfPkItTfqHd7gnEfRfZ
ZUXEpIi/oxRi8QnXAT10L4Alu4J9Fve3X9VX/9lCCChumPtU8t+lGVYbvujZWuK2BZIOOjOblRBs
V0WBIYbGG9BYqiJiq7jWPrMNSv2oVl3vaOfBrnG/+GDyo0Ggnsi8v/VxZtFMSaL+8IDt+ZtaIqJb
D3QZzFHJYAMZmomWPRPa9/DUYiHILUwSYyZIOMlvy/iqqpbZljCEoFOobLA/zmYRsJ5xaONQ6/y6
HGl109mndrrBtaDBRVxvQLbC5jxzjXU6P40x9wYc1xtLyFJfLRZp0KWc4yGayr6zzudh+3EWJ7yl
xAgDLrE0uKTsbJIan+tO1vmhnzaj3U3C0+7Z+xI9ZAyH1XVFThLXpYYW89JVKekXju3RVuaCjBGV
yWaOk9KpdKAR1iSv9EKh1hhKvoKgQkDkwqoKHXXbqcei/0aNzhqpCPxV0PWGKHAyv/veICfYoRKH
PcTHLG1BaCamcf29zCkUbYQYi4oHRJ3mtGMOqjiZEo36uXrUTpRhWwl9YICrFQuOuotPt3Bywv7A
nqcSbBS2lE7LT8sbxsqF6yZciXvsnrDA/pIIyK8SEVS3+5EfqKcjCoNVo1QpIUxAp9XQcYMw2RMY
YFaMz7Ae2xfIDDFqGlRy8e+SgUVwcoJg0iVPdfw8nWvL8a2NvHOXXHVtn/6LSOxZLGeMQXGtiBUi
SgWFsLOZzw0Qh7lR9tDuc5Dn2xKW/TB/m3HT5v1iBk+PuTSEn3PzGH+aTVRr9HdL37+OOST5hi98
fC8mb0dyWujr9DlDC+3NvFAq2lvlr9XwYwCHhkGnnp2hnt4v2QKcMh4XxnTNc0KICANXdkaluWjm
H4E1vudFvXA/iSbEqBUuFkBY65KBOV4k62FMtBNy6IKqWSBgsRku5Svxn+zR2ZeViTI7tnkcJvqw
EOtXeowIuTxiQxuO2LCHrJI0qeURNq8XL0DhaZRMtplhgUtfnf2BGbjzGNGD7vgGgpGiPbTtSPWb
mqEKQZU8Myzf9pm0oaKV2GO5OXE9pHpudUCp6dgODYnIaZf95Kpms4LwoHD1hiZ85HbFnGwamdua
Lar0BrsKV0v4xpt+fSJtXG9KfQt6/0vHDCNyLVWMNGCH3xOWZlH94gJJVRFHFVaf/aeExLMxuUOz
eJEZowjcfAJ36zywjs+5058DNarXApgiJGfoNkwZoiA51ca3SggDWSR5/j9pQN6iV4hwkVhjqFbg
fxcK5YvjZb/MBc+N2UHbgCjJwc27mhOSrCskRCZnpshPxW1QX17SPdUjE9fM2uRAuM60xa8iIxut
JNCLx5xHtHYX65KEfdKoWL9FMl9cHy4WKs66YHAjEECooTNbYgrTvP0uKlSqqF04gN+JSjZVAH/P
gJUH1w8O0MsSsikB5T9R5v6GNNf/DdRsAtEPvAnsHqxrnvA6nMg/oWAOJr8pxccn3RnPSELGq155
+GV2rLeqCWqq0Q7SR9BkOZDMh1Md3hyXVLrlfebxWcemtN55WjQm3YtWRo4wsshXBxXrrmCqvXNV
iuJ3BZbHTssoKceQVYeH5+0TK/QZSc4uXGMPVllbkIPCxHSrea2XPVPlnVQiOxKWM7bv8wsM9mtt
q6DgeU2qV3bpj4odJvLCkNdaxWYQnEN5LCB4r0jb4aFeLGTDK3kl1gPR5sV7nKTVS2mpLLmoUGbA
ha4SaJnbRE3lm54DLgIT9uYMWx9GMYfOaw1QVcbm3a5uEcy+HP7RhxUzrsCNoldRpr+D63v9kt9g
uvDX9mDrKl/2RC6PR2RxC6rryRE9Cx6TKl7d2xZ/LzUMxC8UeR7/aVypTbH+/Lsxft59T8htkC0D
sPxFRr9wNw6d3XzxmQssmfCzhwVrARf+ncRZv594hCKoVI7Rwp5TVuIg430qmrbknfKGQ9hAXHFB
NgP0lPmc7mL9PmxGElhQSQMxCuSstfUA0tX6mbPvffS37dU0XrhbozXabGYVFI1+h3lWOZCgWVyS
LeOU26uFDRQWc5QdbCZvhHUbeo5rv2BwDeCrMgrY+8RG7D4TY5hbGI2uu3BEPUkHG6QTV5iKqIA0
vsT4fmdgleOnD8WMUcOCbOtNLZXjmQ4nEWKUClDkDCQ0RApTeJRdslQ/9Taj8MJX9ha30qYFdJeD
s3F3QNjdki3W10RmNefjNhyTMjsNug7F2hw8O1S88NDfB09dzZJK6rAAAunvHP7F8AV91UBukpRY
xT5OCO4JLH6RwCfRhsa500Ed41Xupirx3p4sRoyF5WlisyM5KmIpvzy6/to/UfNziF4JU3sqkNEP
5SISG6HBmW68PZN4gvRNiN2mi5ryYBadKH3d/Pu1iaSYVKP4m7YO3izpia5YNpfnECs8MAKJzSDs
p7fwcwuXsU5zFGtVZ8nGIP2KP5XwwcZKddref5bck3thn62AVy2F/0Ct47ASLwk2uObsqxXmb6ZP
ai+uFjfe2jdUicZLYC746J+g8G/gVuM6G0AgXzoX8Gdg0QcKDguAQ44aqt/GRn7T07nx6dL3YgTs
IiT5R18q5rSd6aaFR4zLkYLmk/Diu3+GrmPw51m8FX0yHxrgZGHUUghSRD+4CdreZapC+dUyM7t5
vhNOAoreziT1jW+8Ips3ZDNB7FGhqs0yhBRGJqp0YMdr1u3m4FCmmcAxp0dO9NiWD+2uZwak/AbD
Ag1QSpBXX+EuGKtXd7twRCDtWaQeyPl0EoJV/dw7VIWnZvfJOIBbkScoVMcLH/JtcCVc4UmOpCmR
5TZvIYJ3VjhHwzpeqh9VPbBs5GPk0ziQGur+lDyPzn5zQ5G4Wm4ZfM5mCBLJ87cEkX3/O9xD0rrK
6oopME5bZTiniPSBHa8zlKFK/lhIJAojCHf4cWUWZAFQ9IxI9WJXm7tYagWvJcjGzTOtodEhMhoa
2SBkAeevcuQBJ2SDI+DYTFGKYHiS0fvUjSSwP+KYBPCsSydhkqX5WIIlq85Ru2pbT56rIDUOC/iN
Fs7z+4v98Rcvf0NuuPy2tmy3fdtFbEdwP6sdrDPTF0PT/DdW7UMIKFkYv5Ounuegb9cZ3rAD08wH
u6MFB7HlX+N1qiECqQYa8rt2Pw0dtllDqN1+Pte6yj2GN2p2nfM2mOO/0Z1GnGbERs9gtFbDXrD+
0rI4Xv23WvRPJFrajpNZ+l3TJznpi2tSDAasKBkMGcJ+cVlV1ychMx/NkwlpDVy65QBACVgc/9LM
7E/PVzP7pkRFqZgcE/BQZ12yi68tslhSQwCtFhtsEdfshqLeq14DouuouPglQ8PRarFf0bNH4c8j
rBdcO/xl1QrPaSHEMjgYxU9NI6oCfDv2d1K9rkN4p0aQkEfPBVzgdYygWOKMfXQcLctc3Sp0kDKl
GCvG5ff/OAtMh5TlT5yXW6kdn6KWbFZHoZzS8TxLX2AiWojs+OSpymTuCcCglTsaFBfFhLZYGk1Z
O5O5MVLXs60rqtG8Ij6WSdw/lbwBWZxiAyCLAngSrjJJVoSwV0Wr65UW8wdozMCYY4kw6TK1Ry7h
2XKBSHlEUc+MfWkF4AL1MrX9jwJgWVFR/VxDMEXW0272R7+PCnhRuyj6fxkhd1jE7XpS+hB+SZuz
khGNScer/ROpjY4a74u1EGlwjmEt5bZCHTlGaKjXXg7bu3VrZ9QqlXvIWjNkaHPhlZll6Qy6kjFa
oVtn2LqT+6Cv3B97sHXmFKE+C4GU86aeI1nFSGyZgQJqmR0fiPlJRZRe1Gi3IfbkcLdYLd/a6EEu
pkelXJhQ6AobksBZBz3p+LqSUTe0LHIuN45wkYjSpZRyZ+Gh0OijGb10Fp2qQ+vs6cxRSUzQ1KwX
QOC2Vfr08HjRnOLNuiYakHxqOS+s7vJlK9sdeYSVUJlAYdsKDrQpyoAwSlQUyHqYi5Cj7Yek2avz
O18SVI6b+AZaoCoQ0C0vqQd615XzCTly9SfPC/Se8RLk1mZ/NU2xxzGWWgTZuYd+aoeB8aW+4gAs
SQwknuzw1M5hU1h2RhYcZoNBuV0KIFVZ76j+JefjtzRe846ZuFyvvxKrYBkLUPgbKHNzCqn+sYW1
2AbDeQ6F/uLLBsU/OvoZ70ie5s0O8TvN2Q70YI3NpMK421A69z7LoxRxnvbILAFTuovQo25J0Eff
WF9cn5V5ntzybtk581pVtsKD7nCClMIZcnhW7YQ7VuCvOCbziMOUMLB2c/inV211wFxf7/B12bFV
V2VzV74kJ00MrH0j+WOtoa6uC/AjiijiixKf+1Laxe+8YWZLIOcvllTEjJEFZ/vCI6RLxmVfzR/h
jtMNgewoira7DND35hnv946+UumPSxhvdjN1v/iQ2o2Ir6iaKUG4WHgOHIVVFcqmQThdYUEu2BXi
r3UmNpoflbn2Eb7yizKVf48pQXZePRxs/Lc5OfLt1EDNcJBsiAv3OA+gtpKx8ZRaqnzN3Jp5WfLh
H15b7u9duhwA9N86u1nTzAhHFk4XGi454BNdBUMzMiYWnBeQVZ+oDxj40I4uEx/pJZ2NnOBlNKyX
JTIwCt4g6Y4GhR+FtH79u81mAZZxrVFpxm+eu1cM5OVyU7qWXWpMUKAn86cdLgt9VjoYXMh4CBNX
c63N4QcN1PMolpXBpuez23lNVlPWbtptJ662W6ILrh3puUpTaaqF4Yi60H8GJjhBKeqsBMRIZ884
B9LLdbGfzWGCDtkOp0rI1sMgxZS7cDz3L99oHiymFinnDJQRQB+IIFwbSJX40ZK9b+hcju9O/bxa
QQmM2dsc7G8cwWgHL0OVd+WAI0DLBpIGdYPzEeEwkeuQ4XxQOldGHP8HBo0MhiScb696WFvsh0pO
5YTRLINQwiXHadpdldjWkcP0sI7A17bf5xC5+kW5POuwIyzxk2DNoSyyflun8pKklaWDliaU6tFw
uzQ9pLQl36ANVKUofXNghz4DRiUaqP5CkgIKsFOG/3DI/0RVN13HnbSwugnC0gT/3QaU1xMu1jrO
4h5eaQYW7NMccJx9+ahfjSRUazGKmlxrD4ZjtKJEIpTlhAkmazgt6cS2baExdy+Jlnd9RDbO8vuI
zA+F3qdMFYEDJDWnKMFcj2siks+McF/F+UsZaTYEzPPoJ4QomISU2VBFeYtYdWagMKDVtOifXN1E
pWxcYucg2Afs9lDq7n1p8bpgET4CBtKJRrqi9uavPg66xN9Eysaeq1V/mURD5bq7o2SjXMn4aGSG
WXkk8qTSN0DTUHka8TG0TyAko/fMSLSBdL/v9I1VnZJyPvGOLfbSc936kaAelw1Fv0JGh0ygbhqW
S5LEZwCMHBvWnqr0j+Lw2D7FIkY7uvyPdckDL+5XDndCl3+Dfo0IvCrC847Uxuk6Z7ICQUjdYg7U
x4Jd5/Xczn9ibezF2o+XfPQGc2zofs1dFuKnP+2jP6Cd5Cy/5gXKAtte47surLvjL+C8/p5pni94
oyeZjadxFpYWiTpcKoVmewmnmDlDnU/oQSYiGEWBp4gN+8YZKJ9Hp5r9j6vWmXA9BfnQ2x4fGbc3
neACR9RRFhJa65aFXLiQt3KTprn5DCdFAa+Fyo0kMcShm5ReZrNFuTwZIoKQhEsBu4gWssGshemL
SOjULNyT1UmPHhtwaHlYYYfiDH5uWor9T/x5oVnGYoC3VPT4UpRqUJrnGh7swZLCaLLE/dbx4uAI
xd0UZLUY8MjX/WI4hBKiR2qKmoy2liHnc3+s+MW4BYU6ED1o/nWjLzmzOk222MsbvQMSq8NgmU7e
RK9JYfFpby1sxoXlT0K9AtD4QArmWA4AcezATINo9LDDkmB/2SyM4gRqcRGIlLlsKd62B+n8HsaD
QsL5M60ZYYMKWBXveWuQx6ALlEIsJlO6LqlRdokU/KHfxSZwXe2qZEmzaDRtGPqzZ1ciE6PwLhee
Vez0BF/3iE/cTAsssAbxbNofdOAYgzyfGpuyJ32cPjlYjhQwjk6hxfelVLd4btx2DNbqar1M/GxK
CcWR3O8U/9/hLLcIJj+rDUQjUaNPSw51jnUnb850zDca/xefklhv6J4BAcWNn2fYP8ecC4I2OVvT
jxLtZjmCx4lnNV9MZWr3ro2k/Gq1JE1Cpw59Ubo7npCVgrE2B99BKUGd3DmYkMUJmnGhhgS8t/Ir
hQSxgUbHQVXyRayX1jfu6kwhzz8gtLcJY+Oi6U8ckuz1gvd7rR+c6WKGgEetrklIEC+eSHNvi1Rh
3CsNIwhLzZu32GdxQJx3YmynCtqkHmpy86c5GsVpUB1x/fmgKepYLPHSHP0dYkwK+yhaky3f3STj
nlzF6XHYhv3U+sqqD2ea0KllQrrXgZnRQejKkfooznohOcow1k9vuHxi2gEwXnYtOAqmEpQKXFLV
2MMMX4AZTDp8ZZvWqMMFhUPkW961WgVbOp0jFMqAihF4tceoxB5oCT064YJhLL0f39+RaxmTlmiW
XixKFb2Jp7MG4y5gVD+OKRP5Ea225ZcCa8K+5GoM7Dbv6EwETTfjDSQP9n3sMcl7s6yMbGVRYvCi
RAXkfqIsQYGBovQyd0oPXOlhiKUhJaScKGzsvMmwxLMYDvccb75IoOuaZYmuj8izrp6fNmgHkqGz
WSS08Cnhz6JLpEhZOxia/WrggnixTWg873q4akFohoCNHaGkisB3XLX9Ze4OWNwHUpRKp59VUZ9n
6pZnkE3kCP4GFnBdwDpCO956WBm5p1PeP6PDjBxN8rpkAMTFcqu+jg1m7D/+xe9Lx62t2PMC+mSj
vxZUkuwQoH2onSchGFoq62SsipBLXP1XtjHJpBL3TeVVwhsw5zvoBSz6DyItonQjh5wtAqx7Ms4u
sxhxt2orVB/RJufCuLokdQT/aJ507CiyX19t+jaWRR5JhyhqYL995bCaTSfaCSmVikKibtFuTbDs
YECXR0P+fuE7jMToedYQLuz1MQL8aZOKM8PH+nBicDd6u7y9fxMNNmkfEcuBsTc9gnJxJNNzuukC
NNgchrN2Dw3ktSgtZKYhAcnr7Blhr7vMGjiI88rHiAQ9v3YRuNbhseNHbgAXLMnipQxC7mbvfmWz
V/LvbRM3gyfMg7h3LRcy6tmQxLnYnXN5CCU1G7Mm6Tu8RRQhuci2nf+6MjX0R/NTApXH/JbvkWqe
pOU3Hy3mjkCsc/Mt+1DEzT4DRRKfKeBgeHQFmY51z4MtV4j+47MkF5nsbnWHSvL7u36JuG4EWSua
lfYDrYL31mkELIGU6aTQOOHlGAVemjluve5A9xx0Y5B1bfidTLrVGfN3N0lUtg/AJ2Ahv2xvoD3X
7WBIXwAlrZCqXCIaq1BGevMXt4CQXRGcWfvehI2zGEpHqMV1tT97af/38BeJrQSMDVklNjZg+Wja
n76rLzzprTTR4W+hUMCwOyJ2V6rqkFjNc96DrmWuTkB4IX3FdyYkQCEWjD2aS6lnYvE97egK6n/o
SckU+Tio/GxhwIwx2Sa8TmQ5IPnBPac4rRg6Il3QtxLm2A3lcrW0WvIjEK6a5F51xXz+MBtnVgc6
QbgyhwgC+C/TSlho0ZYjMhruDyDrAIftGtFH/eRAyHeW0v7dRFXctVKN6whhYAUvZM3QsKRQhVRR
8nfDJfxVDAMaEBfGW6SZ3evELPzQXm2a8pE1ySx5mMJf9DXYW2JHIGHIFtRjd5LbP4UAEeFTWkS3
GoqZcWkIAVafPyIjYkYD5U470lGQLDuCRn/iVBscaK/N4X2Dr9ALDrdoWsYryMiTIYOFTMls/wAX
htq4PlYwBWBTVj6wgZG3EEelItRuBdHkgJILcDm87c2ID5a8/S6SMuoIcYbNzhBfgKyl95Mog1il
EiBx/1MLjUBQm8mrdjb7GjDQHRyajCKuOBd9Q+P6nfG2lbezZxb1/h814TGGiQG+u34Sua+Zf3Bw
NNnGFdmU95nmyiXTSmVIf0ycMF8ah8GxWqpxXzaD0V40F/onlvmggLpIcMq9iFHZcunu/BXrZg9M
uUyIaWKxxEOlx4eI/xVJLvdl1ON+7jlIE2L0NIGmi74/yQTn86UX33Yzyk/TvLjytV7Zop/sB3EY
I0KIOk0jj2fgE45oZ0fveGd3MT1UXvalPET/kMA7JsrcjTulog0ug57WucB/0WQ+jIHqO9f2y2Lr
Q0A/qqoVeTZAzcBZ7Qwr7MaKSBlBfM22T5l9vVpxr+z1+84lnTTLg5BOZ6uzXoTKxZDjRSsAghDM
/yAbshCA37eUQSyrwjIlYnR+S8VSmZa77V9ViBHBLdQsTTK7mEURpvdFhpRmtGAhvXmcB4n/5aRM
k6ds8eY4Bszi/zhInzH76WAihZxKOhw7Hlh4dIIG5TNErPuXzUv58JT8CwlN5xi3l/dyT5IX+xDp
Dp63RbiJbkA3TsPx3TRuRNeQO7sS4nvj2LdbFvGfTn3UBB4hqWIEaaqYclDcbVhagp4is68f17Rk
g/S9Bg9bvDjT6HXdEGTbuIJhJ4sKwbssKJGIsVXQfkKdAW1Qv5VtEo1HRLRKlv1ZF+2nXIiqH4mc
qYUNS3fVpgp/p8K8HDdMgehRzi9FaJ0DMbl0wfEyp0EblPXc4POSi+PMySCQTL3Kt5q8qdl0NI/V
ijjqSLNkKlyttS8cprcshIwgnQjg9y54C5Zbvx+FlttrtS4NcXbrbyoCFmZx26p/X0XJM1d9nwl7
Bm2pyHqfWXLyEBicMUg2SCW0vwmyz34ZZm1CZqFvSzEfEZJtNoKgqDSdVeXDkcpgCAIUAq/70WNl
tJY+9c0nMLuQLUQLZd1o8deMcFG0vtQ981snRnXOD9MJ23ag8zCaAqUWn/LNoAq1T7v/WUsJ+gXv
/huJPSJ3AmhUJJEtnBht9yMEBfE/1Nrcy5Az3q6zW9xnG9f4YN6Ivig0iFe+aly79w/Ik/8j00Py
nqT4+VhZYJAl/tmRH3kiSXeaxpwtY9gVBOHBMbdz3JQOCA6G2r/e5MLBOWMdqSC7EqDyCAhoUtUF
T8ADAFuALCetuf23El6VHt3HCg4wVAuqBDFOKAt9FBYz18CBCjeN/+5jo1cHxEj0wsct4fRPsKPP
3WOF2U4QEtfJ88PnFhUAUs0G7AYqVo44/TjLLo5puvplVBd/608O9oEmkonI+190r+CPA867YREe
pKHN9WBVGDUHqft6+UNcAd+pCb6auKYXG2ziIFaCLNZsfsofenvBns08uzQvlj1ulcath3MFJg9C
d8jl9pwqoc5xBQ6f073D8Ad4ULZtry9oG6SIGkW2GFDY5nNb18/VSbFKIIfwXXsckMil2SOAokT2
XgHGq2VbPNb8Bl8iPvu+CrA39KGcxnUKDQHRUP/gd80IOvWM2eeSYPSb43REjBXVio3Jf2Shn4kw
2ycghw6fE480UYNk1wU0yWhCL/kjJXzd5mltRuehCKB5eMYbr4CyaSusvaAcC4jNeiRZYqUThErK
aAAURy70bsPFNGPjxDFUuQHEMVSe66scsxSZpXy5Dhpk98Ht0QOLnGOZ9JFmfftjBxJh/3+9YHB6
T10HFqN760QxwbL1x/8zxPQIx6TjX4+AFK2j07e1A7ufur1eyqAKWUdmspuIBtIrHtON6pbV6Keh
03fEtaSaAo1iEG2k20CWfO3rMijdDyz4CTi9z+o09tfCcLDYNbsUz6kUjzELcwURbfJ2P9vodcn8
quXaNNhPZtBtDDzrRFJyaLKn7E8vzxPesEN6Wuro6kRR2Kzq4T6OBD4AQHLhGWgwFoonVqieXg1/
tV/KPmC8VF6AdXNQs9SLLAwNGQvVjT6mkUdqkV2iflDrwvoDoTHbw82eIGpi07GtTT7ub/Amf34b
d0Dy/Pj9Nrq9jlQOPa3HtWH8L9qzDpCLsKK27zK0jkk3ZxKKnxPChQXneHCYP6E2o3G/61tRuRfR
Ik58TlUoiKtv2KqmugDGJWLvUODT8IkswR2/gG60roGm5pHdHiYa9TyYqUDPNOOrU88ycSdYKF9n
5NVpJmHTLlUhSHKP9snFe1larxHJ8KZQZRUh5XDmdhWm0CbPz07dOEQIxtMFuCgof1+ifWGLiThH
rTSQMyKgh77qWXBFZGo0fnJNwxWBESTqbTRQtDndqFTLou0X9M+0TdHzF/xy0MtXLUiWKpweXjPQ
CxmbSpKLKEQmx/S6srbEM62eqr/sEXHgNjW19hoB1cxRBVM9F7I+v43s9zydNoxTASPMJJ29fwdR
9z30qCMRxHzCFw1YIfMbSfjwKcidSUKw89ec/RQMXWF7KF2A0dKatYhRBXSgKEc648O8gcDVgaKU
DtluKBat3ctpA6/b8YE+Irs+1yrngjWk+xra4gDxKg8XncbqN3F70KFzDAYtUhUbev3l4qwulxrh
XydmJSdJaXOjptLkcjfx3vfTN0lmMOEeUBpUi7IKd9gKFzKNmtGppetkyxBZ4KDQ2xFtpBlaSFK+
TZ4U9Uh7S3w++cDL3K22NE4AKgLApj5R5zB5p6q8R2pGfk+91uMnA5F7aqK7w8Ce+uMgM6FC+13Q
8akjCFC/nSR/7eBuy91bUJlYTopk3+oMYyeqdJPuMyZUunX3bjNzP88cPtpGClXzSG35sknHaeYa
ms/WRg2haJgaw9UoV60ISMas3xLg4Y2r/TWfu98BLNmJ5/EsHfoF1Yb67dMN9WO18dCxgAXgu7wf
0XIZVK4XxInD92eMRA0kOS8gbLIQOzgZd5J0uLZnZCMr2eC/tuuFIpEJHlBRYgu5q2oPxA440PE1
s8coNcmmThYbGGtuc1uR04BVhEF9lhs7WATK16qNBqCN+Rmc3c/VzPSegQmna/jSRzu1zhiv8x6P
Hj5o5+QP1JEzzpaQJn+J9S8TcryVwuZeaEJe5Va06MKY5fJeXVoEmPCDJ1a8aDMzo6iFGU4elKga
OmxtXIjCRq76mGZrfgtwimYY5oXvWAqmYgf7tP2XcZwy/r+0C4pkNYUoXcGykFVnWEpFXlszlchf
it9lHGRO6FStLk1W3SJyHRy+PjzElBMOqFG3v4nHI8cByn+pGAj8m8IcNXJpEbAvwepx8DWlIX6Y
7dXTvDEk/pNBkS4b85Ox9wmkk1A8WFAI3Utv0UaoggISNFC3K5nT4F2i9IUu0/G9+YsImSlnPYbm
IUYvWutpasc9YWImF9rbW/5mwsx4tHokVjk2XufIRWGyFtq9K/tpyB5Ykl6uSf6+whD9A6PZ63W6
k/Kv1Ic9XZvILV2mSnylDZYcwXkccGoKrocI/FKJPrJ/YefGEHWYq7hJUb0ykK1tZNdOYQI5cjAZ
s5USlD+JeYQQwp462bNoaLVUUMwBK9156T1cgc+ujZkJjQ1QAdafNvZazQLrfDRnYcCypmolp8xA
OVfIGFRp+rE1xGDb7PcLLv71TkrDS2EDik1cHgptmkvUWBYmuGaBAtgnyObHNwuc1uL0El+sGL+O
CO5c2n/EhhXr09WAYuAHqNvPUGunxX7YAf9la1gGTnMaTZV195H1RMMV+UHz+qkNIjCrSzCHs5by
t6/e1mzOUTOmqsNYSelf+nPZGeOhTvPdN79vCNqh5PEGVVQNPJMy2fkN+h5cUHP87xkij3nF8h7U
Ui2ltkoSx+Pr8BYhJcQWz5s1XB7uIzssH+gGR+dm8+Ji4ln8LwEYIFu/qZ7L/pcrXhTwdg13HQkN
SjXsC1MJaTQOz3pIy52z9zizzNUDAJi7ClR1a9w4/PV1IfQVWkEnoE4AA0m7k1mEfb2L0ehwpylK
qF48Pzlekpz8Zk0UTSRyB3Ut4Q+c8GlTsvyYTXStCBvCyR3s9F5v2KiDWzaloyHOzNFmHHwtERdG
GgG8eHihHH3JXoG6HNN7dmYAMcsynBe3W13wqGP/k5ommaGzRDy+OOLAEJxdKZkORRcLvNAvhy2S
UYQMYGSZKrIQE3K/Bpj7zRqJOYoGnGohDcBPNQv6sJVTz4oCiFadwyTLqQmAzjCUoaI0tMHcEVQ7
wU6Y05qFEhvAbnJ9eL6obDU9iYikKB6QSSC6cYdPFyLIH60QpUMDQSQOoVagHMcovXgNIZB7aYEQ
2R7e4oZzMeWB3a+Wzub1IZmG+2Hkp4VbQ6FMRYolK8FtAG/n97b2dFDayeWwUbMSh9DdOhCEt89n
uc1ciVsRr3qt4pjEGrIe/ZxXU8M+2XxOLQv9xSoKF07UX6jVa60jyhLch5a80ehx4Ejo1/LygxRM
Cc8uIfmii0gXPJRuZTw+Csv/el4DE1r0Te/RMVwGftSEzgjqbmnwhqqxwD5Blc4BLgh77BV/I9TI
jtWKSk3JCltnJ9XE6W1Jj6lwsnV1nXEgWr5jvZtByLekBhQlGhl1Uwipie1i22E+gfA2tJMJuUii
bQW3IDoF1VXFscKmmjbnso7Dlt/erCW0OQx/fLp/9PPvhp+y4wZW+1Za7MSaAogOTeD6j/clydrV
FX7UAOwqDjXcbgODqi7Eab3ck6+zeRMKXSfHEkVFZ/7E4Bgms08RBDcPTiVwiGFEvmwadGHRcsa7
S2jFeHqq6r+pByDI8pMlyXGhQJZhGxsKFXx3Ei3LoD934wPPEU0nruJlUlCFVgZovtPCtqdhDovE
TKw+JqM0EpvJoZhJGrPpV06tvRt4hWgLHItGdIYThDof3skcS/m9DVdTcUgfX6ikp7teQwrCTSgg
n2LtR4/6hNjhidyqeW0OQeoYGRwVsZsoXc9L+AmeB0EHCXJb7U/cxbJF3c0kHDricto1sHIwDv5+
bxwyOF8MFUV1O15gqxBlmp0c7eofGv4l4rfnJv04l0tYl104omfBgQR1S4K2d24p1Rgisk++8RQa
/iCXw5YWOCd90m6bhwFpVs3tbg35Zh7FWWPo+pK30JYf38oBh3L9+ESGdWlj1rqbEsDfGTg+S/tY
pyWV0nPc5R5vcC8gPJUQY/OQTysDWsJW4gCN3zRlAcmoZERzGBP4HG/VyG5bejAWb+Tm22yxVWLl
qZUB9HSkMnoijUSkedUEfDfSVUZaY6FSeH5ICwl/LgzoZiSEa+nPLoCGq6fHEK0Tny3Qw/q491rw
/UghMvh3S5w53DmkNHZcRjzE2hf+K+/OOuPn4lfYJSMl2MqDvEqQZIMvhBZNRLovsQJkAUjbLO1A
DrgYQxlZDXWUejmJBUxeKzuWwA0KhUrqk9nl5yvNGVY/sPQ2YoqN6kS3kUN9sT0R8B/SGpiFurzW
/NcTIEaQ1IfrIYAoPzh1xqJFhUJjkapWI/SNpcZ2PH+i0frfH+yjWvBMCcqixfxc4bFb+exS/YI1
cxajQY2H7sksInwMfcR9ZIsdAbvYftG7Ko3zF5YjN/j+pBQVwL96veHkbRSaS4UDXDLSjtS/APBq
IrIznJnTlnm3LtPeOlKvlz5QSbLQKMswNTkgPvbVKMeiKAw7s3FItKvjuNj79eBxTiD8apuwc6aB
MFB9pmkDDvOjYIGNouWzMIKsMVSK3f0rqDgj4zDGm1vbBc52qt6Mcd35iH2HDsHp4j1wwwyIehlQ
TUOR2+5wHb7larIiIw+mT17hAaVldPEvZ3nlkdpg3s2Z5KUsAft/YjOexMBvDXbkdQAV8DP1s7hO
UlJZfyVIF0Hb4R2CaomHuglEmIDIRpY+S6M0ePTLS0LVnDmM10GuM1eebuCP2wC0aV6Bjng9UW0c
kZW+L/BcpSA3q0uQFXmzQ0wUBRdvMDrJPAn6zqLZ8p+KXLqlO9BMSPrD0iH3tCREksr+pLdEPbzt
2F5h5hKpBfurDtXWC1sabqeaZfgYk+tIm3UlSoQXD+U2xnpKYXLVeNzbhzamSFcrl7cTimQuVNna
1gclKbXxxmHqkspPs/FqNmKiH1dVYE+lBkVQNtg79jIEp0BnbRUKpVdZmGg4QrEsh+AG7FJEQ9TS
8KIQkI3LrDdnFhPI06eLkIMneAAxT4HGLASZSh8pGIWXxP9nY6zfj+hyZynVZSer+XY0DRVxPq9l
BTAn+9SX81ziO+zfJz5+BQMW3JJLDLJFo4bdecNFTk5tgQRsc3D7GWENFMBrFpX1liSliG6cfFw7
UMKAt16uj/rmftaSkop/PouE2g3wowEW1mwGMMSFXA0BfMBwpWo3iRcNfTZEvI17FwjQt6VksC5H
hTNpgCcq2B41u7kU4uZy1FcDtV3oCwJ3MXN82gvCtAw5ry9IDs3L7OTOJr75fSuKV46wo0tey4GK
Mr5h7ULyjaU6b8CDu4v9H94Z1o0NXvDk5XZk6uZ+MS+LnVE6DSc4AvWWBaKWuj8NfRi25u0r2Z61
KxK1wCb3ocmt1ZP/05P+fEO8UAmApR2Utkj6j5wIQjVDyKCsRpDYCS64IVuXafK/WMyzrPlBv1si
NRS7MvquusYEljS0h1S99jbZk2TmYLsHk7gee7yAYb/z7t1ct/5IgY/9Sqr5Szm7KIxWiqqHBkHW
inmEl+Fp3C6gGefvRRSDQe/SvPADdyO92OMReQ1kKrPNNJqZV224w0l8/hI3mnON777YvWgOwc01
YutG/DX9CX98oHdTDhhIrKHobMXKTyGsL/lXAwJDeX6L+nn9yWtrzcIyr6smoorrynmIJODdRtnX
8GSly9CadqEZiLYoDMJPWiInPM8NyDlcmizleOPQ28R0SacBO2Q1ZDolCYpFJgRMCE4+tZbBzriH
pO7+MQdsvfqjz818YZBLYj75d4tlGOl+tiajPisbX1l+eHqwcVD4cPmaXn0hr/S8v0p1SaBtacYs
dllNAzg9tDz9Os2a38ljQDvSjhTefwQ4reXX37LndDFKuGknbPvNGa1fjSGJlmNFCsZSxktFEGef
3EC+nrrD17xC2eO256L+TnMj7OHB+1Mk9X4jN9o4DZMr8oGIsHS3PRO690QHC1a6qOazqDQMNwyL
AJZDczWzSpggX9l9gENAUuI64LkhXDA5fRNE+CnfYwNzudcQX7YJpeny0/sloeKQTjlTB13E3doQ
Fdhe7LQOfocTlOd8gcnkKuiomOpnXLwJtalsmG8HPEJZrPnpih+bh9Tj+ayge2kN7uy7wZSSEWcd
ij0m3PWBU2inBOchtJt7cbIHI17io6YFSDz3Xommbr82gTcGGkUs5pBxPjAXtlLR5HDSo0PPya9z
ngM9AmUS1NQKSCFZLVKQrGq0hKPakIJr4RogjBm5fm6UnPVvHaiP3T/S2Hfmkd4ELOUIFvw6LjAE
VKvI5lb9zd/Kd29a/eZi5aWQPt/bM0URxZOQ40zmu+BC4bgehRewNy1pZXdD0nezCnWy5Xvr6QRJ
QbH7NOUcURBxhVF5+xEUi2gtPssMc8YgORMIKuZSuxjGMI275a4e0ysLul4fJ8mgtICCH6qvkqWO
O44zQNlRAc0Z2DW9SlFnPcERB3j33zxc/d9UAAVjDKyF0aOgYQwiuDm96vYI1Dgd19dbMxGL0bsh
3Ulu+6innrFmguG22/wCNEMwnZ6IDp46ermSZzZ6qYer8/WTPKJCseGiMgtfeDJWF4AG/N/QvaCs
D0ihzPFmPn5P3+9XDDEZfNt5N+R07J1YZhnGqMccPCYQUowMs2wK8fzliobzCRujwxCy1hio8ilX
GhdSHrnpTg8PZYiOUoQpReCiuxQXAhK1kMFGP/Ya1VpSaXccjXwDAB9vHGxgXVUmsllFwokAX4Qw
UZRUp0WaHfRLSs/prci9M+YiEogScPxXTAab/nx8jCKjBfKVaIB+1Yo3Buxko/cXWWt28Q41O7iu
0LtDn1Mxms8q8sHLyHbfphlhbcSW6H3bwopvBTQ0QAFIhP9izrvms3nDaIJqXAj8JG1WN9yQob5h
IuuE6W1RaRUNqdEhCItgGB+Mrt5E09MlTodSyEVs3s126GljJ5zxMAx2ZOtO+RoGm8uzJCSr5gI3
wz7vu2HJnHmfXd0igaxlGk4Hrgj0Hnm+/fhZu/vld8jSXzbcKxxSXOxUHcdZkL39zpVIWXo1aqbG
+yc/aJLUo6e0QeOmnKpZY3RB8vglPvqZIQiYD2FkIZHPvdaT6XKrI6GuRDrxT1qcgupt3VhilST7
Sm1KlTIDbaok8Yp9CFMaIe/RYAPlOFXV1ZNl+uN4GCghYi4MtCrDYXjXFn9z+Nt4KaDpKpq/2rpm
2PR2hil/RDnjx+BCVbEjV75v0Y3wd26r/NSh2MGesQXGVUfxOW4VlKkbq57c10ydAZpJC9sQ0/cW
8nvLfRQvg+9R3vUE5xDQFIVS9iyFeHqOSgQoRy84v/kw2x9ZVun9WPjk2wzrO38UOicBlFVDKMvA
Seh2eXM5Ix6Wk3TIFM+XAW9RRr9FWSpL6ZOWpyLOC1ngYDw1ZF51HcaSzRxpQgr6okhLbLGHvWwO
tYi63qywjpHYKKiAsxgydnm5bK7QZyT2AyH6mqcYZ76P8a6413Mk6JseyqJ96WmnO3XOHVD2pm8I
oXaziNRtZMZ8YOli1e1R+iRX/NVdvQfAQVgL65M4PsskTH8BctV+vSJ1ldlAcR4ZaVzvWjK+eomD
NaWJvpaAHH9ntix8Ivw3dTO/eCnhWyd8Jrma4uCh3R7xUPWikkVCm8kLPTJBGfbECQ8PrOgIcsLS
TTAJkUOIPBiILd5fMBL6XyIS2ti8FjRdJZRihdVTVMb7fzcpGLmZLd0BNVzGVTnN27SYBlbzmEOJ
1n8IPtncjep8ecc3SwRzmgSlnd+N9BPCEPWKnEcIbYKb/6t97qytD45T8eM/Bu8uq+ox2ee87Cw2
NjaCs3SSfoShD/KJO2XNiU30EmH4vUv1AYQujek6Z7jMmLL2mluvtgs3ZN+kB1SxrtgC2cF1tUoJ
C8RDtFA+wH8WEzF5gpNwBY2nqyS6FR0dVcOOOgiJOXsmHaoPFQpS47NM8WQZzXkgvSAC3H3EohJ6
cbJ3hzvkTONSHqwEIXOYxJoh0wN3U623xkwaMXr+tow3ON/Xi/gk/I61tZrOIsMcRyaR9Mux3XxW
7PToK37Yyoy/rlm8YG1cFPjOuWvJ+QO7kT9lMSB+oYcodokkHgv7q2NM9pSBXD1A7lCNZqX0Q/rv
wcT2vEXbS/BY/T9gPFUD4lY/tQtQbKB9M+RiOydNLzSdOoU7auHD6iGCHRFIiVTtxHw4gXnvEI3j
fRbG01BVvSgfBDJQpfc66467/aBj1hLMmoIu5HKpoh6KnjBd+dkIjh/LL1lgOxbInLLVYkphrBMZ
qfpbn1BFpTJk2jwPbaIYc4Hxngj6U6XPGVPzaT9XucTQuTf6WsLpK4YlRU8FB36uPiEmmoBQpKAH
VvnZm3JMONaFgVM/QYCgx4qCfvJEz2ZXXV5NjqRRgZNX6+dUwL2uqEcgjv2DtrHnkD+/7RhOaMH1
AYVySpqJLvYjcJFFV/wP8vOKgX1ueCKET0hmC1QJCbMlt8PPrNve7P8WUzjmdyFMcDAHgGB1aB3o
aIgHzmxX7kLbizN7N12NwR79WnctmeEilCr/r5ETzj598LPc/l4NKA965u3QzPVGElvh1ms/epZr
MLXkeVTJpv4JOysGyMnMGEvfdesnDnnZ1l7+B66R5ABuXpx5cC4+CslsVhU9+5WnJW97/i0kk857
ECsF2tLRQZm1fl+4PtEewrDk/q7Ks1lOWhBnTWtEc1/A6wCiplxxMJ18UJzhgCLk2ITm2bYGqGY/
8E3aO1bzD0rsVf0iZmc0WH6U3zL96SU+NWd5wCwMAEa11ZGfS6kzjFXlGCA0ZJnBot8FBa779oEh
ICQpJ/t/CpaYnp2Kf4ntPwPmuGpddU+sdddlC7pTvbz7qWW+k3qokL4mwAIV4M0dj+xNU0yfp+D4
ARS7mkJwp7ynFZ9sfKYL9fW+SZl2uF55fv8jksZQKwT6RkNDmfss4j2QqWNT4nyctcEWiDFXsEPG
5XG54u04cJGVDpZdcwwd3qy2eF+6mOAzhr4M52VNIebL/Izzd+o7DsIf/ozBBuRskny1eZSLI5EE
2JiAotLr66X0GwREPsWPSJm82MEkmspcNwKqXAVy6ZIBwH2hk87cJaZrTUVvjepBvaw5nvxOIRQT
Y5cyw0gVGHWlFvGZda4aX6PTz7SlUn6+IaAJo9qj5N8J8wz7uOOfNx4xfH0lt0UT0DaAtOD1AAlD
9EDaGFEj2F3NCGmcNxo4txuGuMPNTbgfLnUzDcugRFpDQmdZndfCko2Sd+Y47pLYBFtH3t3Zed/q
LbBOCDzXTkvi4X+DJyS4IqIEaslm7v/Db8bI8QTEW7xMzEJQ4rGaepU5IKpFaThldgBAwD6FdFeE
LM+ZEwnNl50+RsjW51iEHe68BNS/hOfHQh3cKKaMtstre+P8dV2ULbkJGWnSxaFzw1QFihr4g7Dr
BsAZyUjZax7DEw5ywVVGl8oVj0LpzTaRa75cy6+wpuxqK0aeSKBUgGbQ321d6J77NQDX8XgnUf7k
CG7Ju83mZF3S7DIu1wzhOw+9dD7JqONkctLSh65SW4VxFPm38d2FXVdIf52qjd1lD4CsvhUhScyR
b5Om7w/MeXUi0MUXicqXWlKFPSgj/uKdDl9zoazjaT7NHrpLLBXnGGI8ivT71ZzylRi/Wcsu0+tU
sqvFmOmm9FN9yDfPhtTedNy9+y/lw2hM0zwohyej+fsOCLla7J9SX66kZamzbpPsTcgaoh5IRKkH
lUeY2R2A5sejlHHRcueBDSZ//6//Rdq+m8g6sPio80Z7ZhYJLvUJZb3zr0Y3YWDc1h4wzWf1LKU4
Q9loL6YCUO0QTzH+fRfCBY6R5Ugr2so4ovHOaz4fTK7QEmjenwoDc28Mo5wF6cieSzbktg5hULxc
39eeL3CxKvO10XmQ38ZlabVDPui03BMpnUYDFxo1yWWOll9dUagFIp7HC1xVWD1O73SRKkUuMB4c
HNays6dFBlkS1YgBfrVLs2uP9/zl7xAl/et+nHji4W0xCJJ4+PToV+xm8ka+eRy/mlxE2IvEqb4M
zRcTB/uaxCYW58t2Y502WCbSnf47Aok/SYThv2GhQK84sGj3h+zMJ5/9P6mRMf1lfj0noQ/+UXkQ
M1mdQEbGVWxbmGUvhKss0Sjaym12ylnCNF++EnTzhdKHcUlmYpck+zE6AoHrEnjOq+4kcB5XljW+
Z48ZG8nBVSOUahv1IRIdGCNrHer+QDvFJ9aBMEdJMkeDBewCkJbXxJKRUT6e1Kruv0JoiUqTTbtg
Gj425deT8kn4SA9WugHvtln4gj/ObQErJd2U6nrQetWmXagWuK+JamVbQkaM8bZZuj0ZVliovPe3
yCu/sSj4f+LyNkOMEYhuwcqc5zhMgxSeq8ocO5yy3QaqtYsqXwaKXlW//MuN9ElcAuXqoPIrskK4
WhuwIdDG+Rz1tF3fvXCw5dkryGbdSTUjz710ik++J1Y0g2/+QcrjqFTYiCv485LQNnVb2ZUA3mbK
T2KtqdGiBDWmXcwCGtQVWNzkEXVg4QjNpEm4Sc1AcjWRrNU9wk7aAo+WGwLfeHMaT9UqYrXkwLNh
U7d0yGrDEDnVPXVZvUxRVLqSWV5CZpG1YeK+qMmiJ1QOAZJNbZ9gkOhNIU8LXTvSmzquWRk5iKVl
bXhvg1OEeJZx2G14RbqIsCbQsNtW3LrJKrJr/Xz/kBAQmhFo+p2aKXNv3JjGgONbYzEzF8Kz31nx
TR5du2/osEyEB9ZIY51KjDXhYo7p3peRHKkhqvrmtNTGXADnX7EFjb6oDiFUqrqlJ5vGuBCVe9ea
ifl33NqxCZCiqz+Q5avyd/hSfytVn9Hu//plbZ8HChq1BNbHWqWcCfKU2r61jeo9y5miE+3UMKeD
rPcwXJ+RsvQh8FA+yw4GmzOF9DFZjWdAFBI3dWYFl+g5OuVfp/xmhj3PEGoN4lH1uEloIx4/9067
WBH7uhxIJRSZYDBOCPBAZffNTuprorcl0+4oDzge4QiXAiSIeP3TwSamss2p/JyIWgzZsMmZkc9Y
fTGCoE3yFiof8J3oIvUoCS2GXbq0dp0f1Z5VB1L3udy56SAlsgP8EmRubLvonQVZpZwdhAKF4Bml
ordrcICzSYHO3wC41JFWYOqiOG7f3CJqclItN9knbqYxiazJ+jF5ZZb6JETKJrzY7YtuOGQto7BB
D0J/FDpXtrKWPMmQA8O9uOX62ihvjneEnnxYGm0vZrmTD1gxYhRwNv8aSU0wFfy5O8Kw2I97ZVYV
h0phyex4pfz0a/fF5d2sMcaTafHopRdWCFIBGaIBINusSupXbLPGFTSQtCGQ3iQMLUKpKarjFgZU
vlFzYUYf17wZoKx5TzzHI66jMMMEZoRXq2iKRLWGfZamsrIZgRvw4bMx1lmvwWY/1fq0K1XXYCbj
EuBGIUctlK7SzQhWg8xaNUvhe10hyJVbBsQYENknsoTXqef/ze8tud9sH1NdBWFDcjFxXV9hWhj2
nd7w8sOxdihfGr0QWtMiAIvxPFZxWw9c+2n8Y/ITftJd1ePtefD2rqWOEyM3J7ZKLouXN2ls615Z
xaYPDtLdi/Hf8Ar9KCBZby4TTSjbhxgodF3Xq2xqMbGYYx2hY2DneZCgS9jDLkrIELV1nSKNLTvc
KW5xaTLp6pwCs42ox9odklpEJ8b4kGq35rj69mxDeayMyQ2vkKWxP4UtLif/l2yfnVudoZky8Qag
bN55yJZxVu2XW15SOPBFrtVqgSgYifS870XPB4sB4bwIVKxARfb+oSch+afdKJaa8C9jFpIO8F9A
xtnifToAuLb8rpDSmHY0ztxu10yyAra7rsxFyjUy3HT1/q18d9/Q4pm9sTbm7qIFSbB63tPnBOY1
BVr2jnANjyMvtS/kis3qALIORWGfKxCMf0zcwuMgv+sOvEiKg76QCF5wT4GrljW+M4KgA3foPQ5z
9ORsjMMcWYsS6Z6F5kyJ7Vosd9I/bxXMBPvn1q110kj3dPaSXdWxp9DOV4y8uDXU5EofpK+ejetd
AH/09MLIKYqEUm7sSCAwf9kSUeQXzPKsJMh7kUObkRxcmZYwJsWgr0hLL8KCzH7IpCSvlK/HJi8/
6sa0ZwShvjKwjXDMuTKv06og+Diw/G/XxIu2UvgyGuQR056lQ44xyJlno9DGwXsq58SDjN7Wa+b8
z/6gwRWZTnicXBlXpec2bNFtt1YWHaVUlCFeyXoYzBw9rh9RYWPy02WveBHXZng9aOfLhLefDg/+
wQLdpYvposIIDEb73OVNRKn4AZ+ZmxE2YHveZDw8r5enMdU7eLGPjzyFP0wLjjRHKSeTHi/+N1Rf
ycyM7h9PrbbS8b+L0cwOmodXDklV2kBeWEVuSVACXNaJpdwkyXbPjoXbKPD3GvYMatG6KMtL8uaE
orkAn+mlfU/wDAWjeU5cYpHz+57039N9WHyrG+F+qv7Adxmo+MJVfKmiButNd1XD30ncoy60RSZ4
BK5PD4FtE797VJBtlnnwhNeilr6PbT4EoDKs4CpsryV+/Fq6082E78t2vC1eZ+xHEvjq76poMKK6
uSh4iYJJ1em/u3hdBcYWUTNkuBh6CpLhJDirDdNATRWni9G0eN5CnBKSzEXAtCulU7hVdcvyHW1J
JDczI9h09x65mQCj4WWqwX2sDGLfHSEuoj3ftz9NSqHF5fJQma7Ep67u3PB7WrJwfQq4t8xPE6gs
/W12rGUSekIPf/OdZNidNjQmC56aNii0W7/zFWAdIKZSr1xW0gayyJZDW1WQFEJ4xNdYCgTtbxiK
+0+6ZsTVe6FznP+tinGexLsmYK6M9jL9bCTooUuTKU1T5CZelpYnZxm8gEvrbvnEz2Qz2ad9EtrO
dRlXty84e8XIqwBVFmzKveLInxDD7cE3Bfu/UENTWZ7UnG4wyUyXiI4i1QMt9XRkd/VvyZgI1qIb
2UANOwgJvyrCagOsndzLvXK/Km4F/5jaJ8DuBX0ELz8SQP/wxCa2CU4tY27f2OzJmxYvLkUxJIQU
5+REWkNUxW7vLQWRLuTkbUySGbi8+PymyH5W748Za8+aOf1B6NuZ7peCBt8TyXWZQx28Qr3Tt6M0
rEqk7cNRi3XEj4sepONpDYf2RkcsG7yj4KjDe5txT+3x8/7AHZ+IunqYvh/+84eSMfombf8n4+sO
UvCRa2L8OLv8QQpJBGHxUhRqZS3nEG9KQPyhtg7eJ49x442zKlqdLbOBHpByvpQE3wKjoq/OJOBK
wXwSYns+YKyi2rz5wo8SCOz2ymR0Hpnd0JeCdQPflZ4IgLCnYGU5oLVk/57+uE9VYmsb2mR4exzQ
TF2d5FutPwLu+JTgubVu3R+ARFuYHMX2+PizYoErBLOSEc60+YkBKUvsjxWkfzpDo/VDmXtqPAgw
W72QUllgSSnPp953UvUk1p7Cg1CY+KiTfo0nDH49kp9W74He6g8XikG5xqR7ojKPRt57YZzXtqN+
RmQjBbHwqjeTQTSTYDZSG69SOB8aAewyoj4fepBXz4T889J2LOr0IIfONpEfH9Fa4D0xhGsq5YXz
av/Y8qRHl2XV21g+28ZN7TNRz/jZKgb813CX9TfE1OXO0R5gXZ+yP6vV1DRRKdzC0Ra2gFjnZzqX
4O+PtegWWLVGkZsYStDSJSjP4+TehHKJLdDmkNuMclh9zrJQXKQxT9cnyP0S+b5YyJfmBcyAG6fV
2C1VwtJmGo0CIyVAI7QOFtUGomij122DMm+LCSARQ1GSoakGrQk5KbCTd0SzabT/1DnxVeXAvRPM
M4y4eP2OHeLxVzNB0ziFAu6EicAhNjoBywADb3cvr5NnfI431rzxmaJZxGQE8GLbePhGAkvYJ23P
7kAGwdy+PJBQonhZNDkz6yhGpR59qAx1PdrwFlNluGvtvXbzVE4prd/61siqFRBF1enUBO6XPa4U
QTUvcXf6oqd9Ug0Je8rE1/dM9JicsCzzETUv6ONZq/LyJ1BBMCz1MskYLkXWJIuL+lTGyAKwUs7I
3opNyWo5kM9EGyK+NpBAdOcaSGv6eHEDHyo2We11rk+Wu21EqKeIcUZIJAgxThKRL7a2sekaVByq
VJyDC2yaAZ931IYinosH3sPz28uob17gmymteqL90Vc4UOs3VssCNDM2CM5lJf6gXm0mEjKDCNUR
CBZDAiy9qeFALR1FOHI9yL6csDeFN7xLxFwxv3+kRRvuv+QiNRPhP7U9Ef9nFDNhHSAFWAIG9RwB
LPL0MDOwiY+fWkBXT7U3l7zYvmph8miLcRQ+ORHV/6rquWiyPf4kb4kL47hntF7TRCX5780kDX2i
GfyT/6ztg5qh3Fr2yBdEgCkqAxOKKsnADl6+IwgqrVNpRanHjlOPQNJBAHRklr3VJ5qNvR1S8NlS
Um3wH0T2n6Byek2b99tXXPO4abgg43qbNKQm5DibaHg6lAXWvM7oosXtHjhouAvLp3ydXCIByKpF
wBWxG4U1zJNA+2yCrvBql3aI5BjWCfvItl0G8X3z/oBK2s/yeGTWao4OCRcozupV9o++WpM5Bjou
F7xuiqCWM7SoGvo88uvxjPdydnTg7aSZC2FX0r6N+iHQFJ9AeUFs1pfvJHPj9CimcwRwXLJ8I4ZE
006HDn89N0dmw2qRdmFLumTTYWMwK860a+ytinBP9UyeiA3JGdmUxhD5ZgYJ9jOmZkCy+s9J1tV/
udaXoEIa5IZDlORxy7FDDsTStk7y/xwZZVgB3tXVLllEp1JEoaB7U4VnduKcMEsGChkw7Z2wIYCx
u78IHI4MFWkkDlLscBWnQBB8jAvnq2Nsl+nMI9EBb7a23fiVJnkfkiWn92L8Jj1+8GKX2aDBVsK+
qWO0KH9E0k4UyflsB7u6PwwWhU5afL0JuK0I+NWNeAvDVgUy7A3mbb9lcITbUGl+7AAl0wX4OfLy
ldPXgZJvWYcoXwp+z2Bpqyxu+bLE0VRQt6dxEHU/+GfiwNYqxwp/jgiTdFuGf2i3WmYAlgmrIdE4
6Jq3dGnhaISuMNplfm2wIPc3hZdm6nQQm795kz1aGhaaoIWDuTWgOU8m+nkl6ELRJvVCNqhofexc
b0cYWNhr0dANp3Dcw093qloFf/GQgmErDxzVpV5K+S6XtTKhT4l9vEW44jML0NcAbXQiI34ynrX5
g70wKhhfOQotSza+Gng7lpSnh20jYhPhkne7ZbCJaUpeQx7Jim47JyqC/JWpizv1JLoS2E1iLo+t
YmRovEARR76mUa7CH+afcV21uOtMAzm03hM6NqkU/pMWL/B+ZX0JHsouZZY/5ntTaFktmxXnXwER
PomNXwAQpmDvHjlUbgJWp54RySKbw5ot/V6238KixclwEb5l+v1k4LwDgOF+h6QhkRDSHM6li8ny
C3v64vQUf2wAlWJD3UmEaYB0iHFj5qUIGScAB75fNeAIH2Ppw0QiArqEBUwx0wKbpPRIFJ1BIEGM
3Y4JLHYTU3BBi90wGQCFtZs8IrrksH+jZ/ECaJADWQkmocDYTYHe1zxNl5dDOp2W5wBaiieaatzl
zDXs0pw5Vmwk8LKAf1EZUjbtWokYSapI6/IPUsSCqF8Pm2VSbc3Clk5faZ/uLSAWjnDUtaRmnkCK
Cc9/ijPN+CkesAu1RYFSf9QlkomdSdoyS7gtmTBdYbghWAQqbkcRoM1FxwbJzl39iEMiTDavaeoC
Bdb/FAfj5Xen8HEIYSBT9DW5+OaPlCYZ9MkzsLukIPDKOmZik6WAVEeF+S8F2L/3ETu9qGsK9lf6
rHPvtDzQ7PNo2aOJAVKba8Arz466wrW0cbnXPvHC0hswG29SbumkLm588yzyDYtnZP8VYU96Jjqw
Bx2+3kJZ6IZG5ip6oJvVSN8V4RHXwWmGjoaF+N66z9VZ7gG3g7p289N6Mq6Bhl9adjc84HJesZKs
tyMD4mHZoqWbL3brUEWzV2+VsULy0CIM7BuPnss9oi4a06SAbhRqad2ja3KcX6ZUu9lx2DBZAmBX
NF6ChOAY9fA1PMBx2jxlIWZr0yAwx/swcnEVfE6nM4XEP+a+vk81bOcHE3piAv4rW94hYSjUnmW5
a5t6MmxoD2PZyyZkcY7XCi+3+kHv3eqXY7p/nK9l4fm9q+Bvqjxe8cQQa3gY0DSidR9H021eKEMh
+inX2OQ/ejtPFCyF3efHbFjLrIW9SDaYj3XSaOT+APgHjbmRGmhmE4JEfTjCymCb6KtGJiTCqof3
aQq9If2vRqwogoR3oPw9POcn1kqjMor21B5HYQrPTsMtfPkpmfFjEO/pEk7FV/ziGUWM3NEOcD10
t9xFREmXrNwrv7XVZAogN8tDtYRQ8PzgmFqFnRG6D0fi6jwOKGWJpK7n4vhfFcnA+IdVCKaUMGE8
Ox48zGq/H+4ae7HYK2RK5RXd1VwdQ5XZELDr2ATpi+ytA/1DXH6Rp6ukeDB5PUrMKKX3DNF+74fs
MLK9VsqocyNkr4m2slu706fpp9moP32vxY+9iuAyqvCXc27qnTVxE0o9029twNYoZCLXvzYRhBix
yqYsbfxmnIfzio434grpGD7g2O1eyt6o35GPoBQiQ5duBfRiWd+iJqPLJORjmWc2lf+tpT5NddHP
Gu0BVGKsCs9okxXawdz+mf5EKUWKgvcL2XUabyxvk1xq+YriMozeVaiaXMS/Hjy2ZEpB4CG3Wqci
KXAzUwBuaoAdvfLqSQF9sSrGAn61N9tDcr4xKZFztRbcbGDRJsLWpn1raFB4yXhtWvCoNuY4r59u
9R/TlYayHG2wUOMyg2XEaIa8VDWS2VwwWXfKBX1z/kHVcjcD7qednQiXAB7Vng46qhjuH+wTeQXs
VbgIAb4VI/oCm1/d6Vp8dUWDfXiFXuv5LNx7gXu8nsDEeBgwb2oLvj63aJiWSOTUO5xJ55DXR7MY
xZH+Y4CBmvm81YE7UdSsLQRwBH9ex3Jn08KyvE9BOiVtifE7ADmTJJDm7jIjoTlkEwvB7uXqwlAx
KZzdHOyI7cWnYu5DQq7Tovu6U2oVijdAM81f2FPB+W1UjSe7VFZ9+smmCJpByGFf5surVqL+9ITO
0eVyPy/g2u8ION6QLhdbYSQU6MTsSBYlzdrjkwAk+ufiEVUpVItcb4a3jcAbK2LyXshVQbNjFdgr
LwHCVNIQDIt0ohToQ+MnNrI0dYUxNtA5bq+2+KATcgSfeEENb062jdEKGJTnu5uuXKDl57tU6dH3
qJ6RAsRB8b0/slP6Sc1gM3ZeUM1qq92ZFyxMCsaPPpcrwuuFAPpQXTb1S+Va8RyupEalPgpw2ErC
eCQbm0f/iQSAxUdDrILhFX0dKgmAnmIV5gP4Hvrqg7CUxlSgrqXeg1xQAUF6oJKLMytLVKYq9Qkw
48UCiwiJMrPiRfszZHJDgJXnFJepehH12AM2KyvMKgroPE1jxVGli9HqZvCqpTZlZ12zgKgRYJ4F
7Wb4C8jyJRZkPnZBP1cj6fkbIyvoVdCotH/4giSWDXpivxRDqVx3eA4/gkQYnaw1bOjkTIIhVUYf
KLyQ9860cjEaVsdy//N4+O4zriEOTOB0OQ3phRzT/Zb2oJysEkg5j+5zd307juSiHDPXm9xRCwmP
xzDf4u9+reK2DNFE/pVZtwBVf1eq0zOwNDq+wAnqtq7Nw5fk2b7wRETSCD/AA2DwTyFfIoRGydV0
kwrmNjtr70+1NNFzpLMkJ6DAUAxW0kDxPCLWptvCp16JeSogp8XxA55fvnIOXcclJR7VgtStm6zy
oZ44rmFYvVVWBlGChFD8/qW9yxyB3nb5r2nlo94A56acTN0wQZaljTWzUGcuauxo91J30bi+V0dT
eKZ+D+eCKe4ayrOLcItnisuOKCmE/+tMKH6zC0dmTWyRJ2dFoW1l1khJBKyFidSI22XfHhUJv71Y
YGwTmj1i8rH13FHJ+c35nNu6wcbMMrKwbTO0/+EueWtLExE8pjvlI8Pf9RJiaPGIG/BVM5Xz5FcR
ArU/BFMst68IYV4sULbqcvvAL1+I7Aasalf2rMMCpF50xyKctPAJq2F1Z56YiWUYHtCMKOs9GCJQ
5kzebwjmgqvZ+Y4EPfTC4LPN9JlO8kJQiWb2itcbeqEwPUEhXSGeT9ANxUH80Dq9P2Ys1A5T6ybk
T8D3xCsV9yh2O6GhRQvBu69aI35LNlITxZTHEF2TFyKOmv3bcdYNqJllcJCGGbhKPe/vGTL23TB3
646qMc4xUYaLk0J5dfCRk7nRKeC4zvOLziuTAWVvJecyhdLzxRdqqA9OXAAteF7alLQcR3IA6g3I
QvIP1lD+NuVM4wvyQWzTSNtE2F/ZKhNyuUNjJyUksDLEFONNlvaQR4Lj5mjZaCJSgDyaYGlkOExU
1IZiGv2j3kZSrJ2gWUqPQX2XuAkjRPdXj4YKP29iPhEMk5AxDQ/bOxSfoo/JkrMcr1JZ7Z6bTpOQ
gBWa11iIAzPeGg+vSXigf6S5YoQj/AtipiLW/kDa75nd8AAU2GwrRPueleHNEuU/lQLipjFvnHmw
KryHC1rH46c1r2WtARrMMr8YNySgkqbfNj9nG5LZQdr90b1brIRcdfZni/JmaFfdsWZaP1qQ2/nl
Sispq9azPHaPGal8oVleoovPnCDs/YtMANSGnav7LHgJ2SKr7Jn2raNb9HC3K2xhS//QdJwFUozE
dkJNCjk+LSQahB3UbvNnGARxMEi10VnaPu5NXNk9UcgcqohhyzeFYAyewVwLHDEsoSu4F89iHu7q
yNOHfvoN2BLsQzschCLHxwl0RUsB5R3kxu8el58NDhXAcweBgQhXdi77pGFzqBzN+F3uPMlJMExM
2HTW01IOzptI3nyRwGd9NNJOYkLFI5pciMSO5RRtLJGOVh+OAkTMEW8luG7sfQ2+n8XgEEz8cOSw
azFDFLiMSh1LFCT6Btm7mm7JwKNsgUKyD9MbheFSeUPruh/wo6xuY2NxQBPGqxHt3jqKSA3D3D+q
LsTROTPeJxrwf5UbWKaPbf622UVV97uX0vOsb90DQD8Kd2Ic1V3AHjKiPGfQoAn1HyEX2CuDp7kw
0SmaIEYMI4U/p4+Wmv7cXUQkQCNVpMwpl3zpXvWpS+Kanqbai5yL1qT9pfGtnvlaoU87WDFkAcgG
uXNAusp0E88h3+vnrDE5lrNbYn3L6lOzbxxPrDalmuYwnVV0SwR1S+uxDNuZB3I+xBK63IYJt3TW
ywSxkQ3NEmZ4HiPHRFTS+kO65faTqh1zUwMfC2b7OBzTZZiPQwh3CHyJicnFvmUPtJgRP+gdlF0h
cpba/28X9OJUaXL+JQO8DlAcdlOdoe9cEcKzvBqISq4qtkXsJSfs2PU4Jad4iYTLnyuf9PC6U7rz
pIu2C/he+tWAjoKLpmmeXSDV8ZN8LZZUtqeuRdaxuAj3QwTaf/rLm8SMOc1hTS5Ni0ZQiyuJVSc8
8pU++Pu0vd6XNctdL/ia3x5Ih6NJMiHJTQTasD1kOnZV2PFL46MDgNvJXvEmaWNShu40cml3jIbo
WY40rI+J0fkR4/jA4CFo6KCiBd0qeKQf0NyfednwUTZsvdYQdM7vk7zpbRaL8SRWsvSGFhzMn8D4
eY3fbiIwbvNbdbpvwraE10AeTB5vno3AFf+XQmwVkK15X7bMeiqts8QFS+XYHSsIrsoad3oOreMA
8JY12YWnw69NJIy/YR7DU6vRA+zH72ahKUdqEIRa4fRyzJQOerJ+yepQTssyzX9SclEKjTOQg08y
BB0ohIdhBORL/YVRo4k5TsI97wPk8j18wUdtwN2R1LHBUxImJuL0K1GugpLuBV7WohzHd8C/nD68
MGJFtYiBiylUtzzGoWVB2gthRHTroMvD8XM7ek1a3s7qUb5fKoRisdziyXp8Qvmjk/cjxZgN/qb8
p6hCRuoEFhqDgaa9N2oPfpkCCLyYSZk+yqmeU8VSUuqrtODxphN/6T1yl3kIeOfDs5s0J5FK7Pql
YhrW4Nu6hZ3IVM8g5BGqlZtCxeUVETE86y/HUCI0GGVn3uGMM7316d8g4ou3P3qGqa2BKxeariJf
HMwgK8dsALar0mFG6SpMlWAsr5guhaiMf4nR+2dGRyIHgX66L50EKKgRJevFZBqkznrZDawUCpAF
SHvZ0z131g9NKJB6nTpSYHA7D+ZEG88GGFYFxDR6V5UX5ZROIKq/DH/ZUmppekiaXEm9gJE9j/hY
nsXFAKmPlx2IoGarbdnamXUymrJsGZuVzk0hmTDyqIu3Ryuv0fyHdkuI013nYVNMOqfEPNXHQc4K
PULiPylngz6LhzlJeXqrhgxLU7kfCQC2YueRLzKvrvShTFKjAbszw3J07vsabE8CvZRTOiD9YhOd
0ZinYnuuqCEb8nYtIEVNp1SNrH/fZJcfQMso7iDKViIbmuh880KnOApZLxTOYk+vOFFmQ5mnhTp3
lp7sOdJe0eiZ+3F0YHrT1acME1h0uyzxjyabIHfkiSsoa3uvXf9cYwcXfNHjbj7bWBmVqG4X/DHw
Zbo0B6N9Cz1nVq1vPjy5LiW+kToARSVMwJD3NF6SU9g/aOt4kA9FO/OLCDUaeXD286SI/APNh33p
3uONnf7gUYuTSUbwFeA9tHQc8Wieqz3IIkKLXwIse8w7DDCyGm34e2iCxQLShnoQczkEunHkJ2xg
/PfuVxy0oT9HdKaW2+4qU7fwDWkSY1zJkcnBBNwf1FVokoP489oZ7W34Xou5uUiIVLPYLL9kjDHp
rrObctK8AYCsh1UMDJ754+aTNrxRRT9H0eeh+vOOlDAhZaEUX/8Us9vEtlET3inZdyvUnw9FbUNA
7C2h7NuW4/d+cE4Rj7dbZWof3CwlbqrhcW6zeFMt4AHEZ11sahMx6IYCdhm2c7rO+EhJo1nYkSM3
JwijKXNrv6ILmItueyjGm5zSNeMgwgAyUmdT4YAgrkLZKoZ/qgemLHTivYqLhFoqvjjvIRHcjz/1
lzqjcqk9uvDmVvNM8XBI9h8CDYGlh5AMOgWtiyiReUYTXeGHE4EGUV3dSSTjXCCtb5BKLezUmXIB
ytcXQAOBz5MvVwMpqVznBv8iHUaV+t26lJanSHErZXd6huja5RS5nM+5NCcjNKmErePhZNMJnxKZ
thvZxx5hoygZhdCXkyvMxcrbXTA4FMiXsOPbC51KWCMnqKvncehV+Q+ZZP0maI7t8aLLtLrbV8fl
+Wteac+0+TBhg5PEj2MCiswIhaxWuecvQ68h7jwhYa09M56vwpqM1Dx/RH0skayFfOTGVM1RGRon
KDicDPg10pPMgfb2OUd+IA1kY43tIh11P1KVt5KsGcyAVoGRs8vK2cDAuy0HKcaqduFNVs43LoZf
aNT7Rf+uXpmzFOeaWFLnPQndlb8dAMe9JaWuYZK4LvmHkfxPL1+2hwSpeu1wbkbfj51RgMzrFro5
oFplvDmxpdjLoy5iP58JL50HVvtJxdZ3rsP8lgnEp53t0l8HBiyFmP1ESGaEu0mDgsCqzUPxQwqs
LJKWdG9DGAh4TAtYBcdu9GULtHjyVd27C8x4XpNxcqxVDD6bW2qZ0cQcXfZdsKDjqDzL7pyI/Lgo
PNTK1RCjnZKZ17BJDgBEfucGCrkBnFCsOBecFdt5WTmSS2RmyWHpOhg6N3Fgjw4GcN5CJMRdFxlT
8UZ9tjW1lsOHhv6LBDsMSbFOoCmFS+tRYQ5+2Ihe7MLZYiWqScbAI+arUVN4Wlz5IuGZmoEt1ngv
h76dzfbmNXhsPyggZTbfSixKpMbz5WwtVn2jwK57ipV66oDO06CoKtfthI69IBa8YOG17BVahnsY
Jrz7w7OuDbz7J2HnEm2nb1iVCBn2b2uQWMekCJGC0HdQxMnAwLvG0LUvFypPD//XGgsfIDNrbrrm
SVveXunyYhGXtOhXSM9EeLqMpwP1rNLxLxlauxjo2nz9kUudTHGlrhWmIlnrD9dKm9gFPQLu8WQG
1EHIAKNkTGTHxP2Uv+2UhzcS2Cb+MCCDiUmPVN/zZAv0+N39NdGnbwg6v+ZSjfps2zgxh+0cbozI
8CLeLoi0VIUAS/Osruc24/dvxMd0jvZOACBum2SgvcyGBbIZG9MOKO/5Csz/qhb0cLJ9P3o3ViGI
MmRDzY+9jp8aiZu4rdHpz5H9guChpPxrHDZi30hcSDeEYEjB3c32ChL/oQQLm7n2+iH1m+tXh8Mk
5tCIxgE7I7PiWVKalA71pKYdEf0evvnzK2SyFA6HBkBgew0D0YJxcOAkrY8ynsWq418dlRH6rQef
fUW25DIu8j4xWybTnFDQmKLfpG6kKZKYPIGFf2JBKMyOJC10mS8CAtxf8fHPLMle4vanoyuF3oKd
ZyT1HTNlmlj23RMmMfmzijDxlMCGu3v3qFMK9xLPazvL2WArGwZULtedr5z+fEcSzEgSveu00jvw
tU505uqr+xfDoOMwMpVGYt8Kbp0CnAJwrV7rdLXC1XSJXtBg1WxnyiNvn3py6EZ5cqg6PB/bR32Y
ti83Lkpwmjv9ZFSmCoam2IqtWPjXKYgDZAXF1M/ILzeWtPfVp58CQ2Xc5ixJ/zT9FTpgmsjMnqXh
Xxdib8eTxUetoDywbKka2szfueISlqKer5gUjWb38lP57Nr1NjgC5pNnnNqI3Kzs737uzfvHQFSO
QDqkNd4y0OjwyBOgIPCLfX5cvTBqTllKJ9VJ13dcKl/NfZceXDG4cgzyNQstdfi4oTla87M3mRSo
rvZqVSBKd3UAo5rlsiNaywa3fB2vpZyUrfWqmfpZT9g1eG1LLk57bmydP3PiRQtmFmHnD+lhsaHY
tH3s0GD1WmE9Ibg9CMmx2RggtYj4K1ai2VP4/rxXfn5Y/T5VlH8WNUVaJf9OG5SdZhy96qdtW3Zf
2sP+xcfCNoV1ROVxrFG0xwMsQKN+c6rUmQYflJPEqHPGe+OkHeHDCroh9xURopwR2JCueksvgXEA
xD9kMA/dSAIxQYBAiTJjV1A9jYp+eg/uXR5oJ/Dor7qIqUytVKp97l5avH3WMqNiVaBUMi5Qn0nl
paaLWBN5SyDB/reH2hO4i3HDtLCMc5XhZ5oKNQGbm3WR7C5f2aD0Z4/LC5ofcNNul27syxJve20Z
JxMAQVzT2D2nxh6AjW0U6shhabzuUYl63AWGWoiWihJFkOS4TAMmjnjc8mp11vTW597MegLOSLQV
5UL3wzTYKKgLzjuEAcL82PAmp6LxMQnpW1rPOVOQCMVmUabUn/8rZM4kQG+21fMsPXeNopalG3wa
KWgV8OHnoD/dgSZty4YCzR8GBq0oDI5ILWNjtWmcSPzjlkCPjNUGZ20QwMTJMcE1dG29xWIWr3Yc
Guj7BYvpkx/jxFO/NN4SCUVN6frG510hc6KHHGJswdHZQTc8PSAVYlqecyqV09DWXRT0wM5swyTa
EWhklupVqSkxmOwR0pdFPT2EG9sLn/OFS+59GuV5xy9ph/toVaHY0mkoy503RdTA55jT6KXFO06w
5tsZR01PorJURgna7Og3Q9S+IAQNveoR6NyK6zmaG4EAr2lDI/1FUbgPBLlWjgvQh+Y/KRYYafgH
6Ufvb2KkbxguqvKqWQTgZiOTwzUCAnwmFOCO0DpJa7hIBNha2O6nLxefLhVJUl4CC9NegGQRGLJ7
ZCzWI9kBvojlUrFlrvM5YWCvdFI3nOpDH9iYFewxJguwl7WTmEeWm857zdDfgIB9KdP88Bptyk0h
MMw+ov09weBC2xEYym+PbkX0Iv9jM3aEqBH0XfTRRO9Eum3PeRQoi2/zfsYBWwnFcWt1EkCcENYd
y4ZsJf/rcGmN2ebCNSndd3rJX/MHD94boScm0oD32az/BcpgdUKZez7wQ5VuDVzzPKITVPMae2cw
gK1+WjjbtbF4J78YdHKonfLQSN1fcUmhSKp0qgT37mVIVOJRmW4XYFxN0EVS3e1wniDj3qyWYNs7
Jn/gkW4un0fzzDYh0qQ0Mf8qt9xWDfB5gWsV7SvsSrmK5x83kBJLA6LGBoWgLGcNvgQuh/zcz0c2
se1pJE1fJf3a446HthD4l/5ck9xUz1B7/4vQD5tjPf9F37JTe1ZjmjNVgV6zp6dIVjH59UiK+gtD
7kLTqXeT+4AhbjVCuhCrFAvv32wh111MoOG+QeDoFk7ni3n+USd9GXzsrw6HLXYRZuV6bDP0JcMF
xikiuaJm6QqjG1s9i8n2Jz52cyvO+jFx/sWGqpNH5lRqDRywd7PfNa/inHmYnViJSgvAtMUSBymM
bdRT5Uv8F3XROMHERNB7RXq6G9eUGADPcjcabl03s59kYBilQVGR6ScEWBGwWFxvTkfQouj7b1b8
p7h9wB5CctwBqQ5289FS1GN3md9Ykb2tLo/VxPdCRCo+LcanuZ+l5LrlgU+sBFxSReIavmbOdngv
ckyt7BpOJCiFMlqT5ZZwSCq6lvGsEA4rSb3PSAifnwbYlQ8V2ER7Siw6pFlX7Kl5eaa5RzyByeRf
u+7EvmY8V5PBRJ5ygNSrL+aTLSLIsupbKgkPwICppmViiNkOXUyZTyx7hST5Spc88jojWprtV0V7
64bUQ2cthh5OjhwcGsrncbL+Pm0+OeZCzKVAtKseBzhP1phT6DwKrEmRMdmJh9pT2IogHV3le1rP
BfthAW3GTR5MpNpNF9HI9yrG2/RrQhc/ORV8SjJ6e3XkiAsd12ZtzWb0Mdbhr5V67/UDP7Rqu+yQ
7gE5+9Dg4D0LqgSCuG8QisisNqH6Rn9BB1Lxj+lpeixJdodqru/8Rxxtm3v5FwxNtKx1F1ilqIpm
l/QxjvaX0Ugl3YrtkHoOyXHYv69SVtPm8OoE2iM00xy78OthnULdgyBtgr4bAyDUCOYBXZMW81fi
EmSJhjcjq6BvrssPkYy4exZpXbu10bqHvEM5hfbhP1heXRjMyRjovnuOFl5OsHLfFKvCBTY7cBUR
V9E7Sd++4qmlZe41Sm3i0gxnyrWYTTjyZ6LUTuEg43HVQkHLRPtlrQD1PYw6ozEqfJme7FgI5gHn
8pLLAJKcFGNhDptLyUwVgwQ3gaQSnOSJQc5UUX2APjNQ2hHXYjoeO+PqWDaDzTRdvsRm5PvyoFAH
CNpgzP3d/dAt5ihubkBJG6EyookhtCvOySxeBf5dvk5TOOmYzpTaWSuRj0J9QXNeYjTRK9p2koud
ukj2GN6Lm5ZpMbcQ1wyRYaIypKSb2KysTIyXmL/PlHAhQb8JjxXYg7TBGp2eDy1wDVnUGh6nbOwz
w+EukxqMHtxmHz5GQ/eBYO0fzMSMnTM+XAIOUe4+g2GkDhLECS4oV72cnXbRxnRbjMUb8z/6J/FP
ivDo1UAIluhfd53Q09bEHGRqouvNTMNr8x/1q/5Rjl7IrEL9VHkOetayS186SI0r/CXUBSLm8BSl
Qg4Mfdi/Nodk9WVGyQPnl+RGAuTmZ+ZXb/PetVpuBvVp9epc3bdxJ/jcsrSsW33ohp/+U37zrfUT
pLiFXkLprLyguIg3fKCvtEpBS/4+8Gh1CX+3b6MzF6g4WQYM6hJPNu487Juqq6xG4W+GnZXW7V2o
gaV3VQ/ctaf1Hjlc0bo/hu02zmrUne1aoVRg1XVK3UO3wKOSHftQwuOVaHpUqr2s+bWJwtHaoKTK
bss8XEOYPfNAAWbYYjbudoChNaE/W3pKkeQibMDqs0FBRyEM2QKQp9iK6PWwAZZvPJQUQUsB5Bbn
bSqMm9PN9rgtKvKZ+lz9dOVtmJbxDaodjcEy8fdTIUeb1KIZ+jWzFAcRikcKj9QetnPakbWn840P
Zr99tiC6+Rr/fOsQttpmVdJOg5brCG5NG1qZE28K+FM5rlXvxoLoLUZlulmlzdy+Wll7+TEOCsqJ
VdKv85zHG1ecKkY5Y8mkO8linmb9HqiLPigMJZC5RedfdEMN1lYV5xgv/BiO/9JfWtIawsFQodTd
r9zaYPCHkOYx782lwXmclnLVp68rUFkOadZqoh763aNI7ugECBy+3VWBCfNc8GnWSqG8hZW27Cxb
i0fZ1sV88szYz2zZKlgrkVbkpA+0ahh0O9ztBW3kvJpWa2jSKZlHQ5u/ISS83YTashYp1N5Y3Svp
QYjzLW28gOTRctbdH8OYikCmXfmlXp83k+y1eyxJnfUWCuiCMCuyhEM7rhPah9yY/5AwsjKkiYKn
uD/aSulzx40iqzwnJzIhceEciV9MnJ7mQl1vW5pM+d+GMLfy4ekjw7UGsGC7swEc2u1L9N2ZY1im
n9jbPYZTri0bfCi9uo/bY/duGaWDw/JxovtWcEPBmMtkl1LJu79DYJ4/6C1CIbBFagnjbT4vAQpr
OL5CvT132JWFmTwBCH4TrPrGG6hprkD8m+aZBqEDgBoF47BAE/oVrs+ClhdVN4yIY84O/M+uwuak
tX5JWjCn112D3T9w497/UwLoLTSrlfF5d99Y2NyY9HdApG8cf2vAzdTW1emReAgy194kc9/qftlt
AavbpUK+k8SYK/wLZKjUPydCgx5aJ0yz8TZ+wrXSkFUBPSULz3WcWMPtNT7GcWt2umt03SJIdTTg
iV6yIh6Ayj+0hN6e3PKtCbGfOIEJk9x6UZBOIy9gkOb9YeW6Uob6ChRgetDVuHWNIfhj25vMmNNd
lfJCraTB3p7Vp8xJPtkmNkCPX6TdcvCmc+diB53w3gH0jSRowmPuTH0y1T3YdRY1+Km/mhzQnCCp
Bc7fjePNBnlfxVn1rgVbNczaEMs67pFsYTRitAp/cP/hRRn/iL8u++4CnTqU1wUXi2/v4366OPT6
IMQcxiDlgd7JDPo5McQL394FUfsKTL6J/Kj15rJGKZPJmORUTd6UjOZYoD3l/XzDIXufL7kbIrjG
dLRspbigRooOsW32u8YKMRDT67GGG9QFmg7KB2TS18CqnUx1GbAPGT5YQyEH8jbvLlSCtWIxKcCJ
FO9PU8YnfM0WNE7F7zWhJPoSfJdeAydWE4HpV+is19N91GmLakeq6DjJ13hn9M3ZN3zEQGsJPMWa
RnsHA/nPbFP36ABVGEIuvo5v/IUTYHcl5zTBo6lZEazYtC5QLHXuIAQNVirAuSkfH5XY4l5WAisR
yiJH4yY9xQWfhiYEjFv2UDx/OTmal6EWpM/S6jlB49X/ro7YRQJaqwWINd9F4e2dlhQsZFFK+jwq
g9JY6PYtyWE2AVjy0aWh5I6eeGlx2Zip8fCCK4aSY8j7IM72ojzf5aCqVq7Xd5w95AMNqtxkPge7
7CQFuO5nJpronxdQSuvwR/WVr9fhV35MWXcCLrguRKqAswTKJS7DmTsJQtd2RfockVxvNxmV+QLQ
Xp2R7MAH2ww1GJPpP0GHgCaxx5ZX2E0pNHdFcBCbTkk0n2043HFBt9DdPPJ8koegnOPetT3zef3r
KXN6gVvr2G5FZTbL6nredIaQwPA/sSItl+L7dpzbtNx5VP5O0KOtNypYbswKvpBJXYyNquuKShyd
9WPJUeMUqUJ93Ba/KiRheWRE9NwXF9pzpoooTD0Pd2w/Uy725RaFd/j9z+ORQE6L4qJb64LL5xW+
289RhAJZaOKE2PQxexXNM85IX6iF/HJp3xkBauK9+AetLHQr7Mnes/03is3YJbd/HnascTzfjhcD
PFymreBTZ9DVZIwQZ/onMu3TbWlE0ESVdKlYQLH9QD7XRF56gKbh2zeT//vkugWHzrgHHjbUq6XI
aEZnVu2kecwX71DQsTzCNoHvv2rdEE9N6boTe3n3Mk9M1vARFw/2HeUplMCdn3LYWxIzVXcM1HFz
Gw010QWrDgNwTLyHHm3cRiVcjgNoBExBngNn1uBcy5nVYpu2JFnPfwwf3LecVHk6hcNoy8RwS+Pv
63Bydjwd/76hz0gCFOSPM1+z0uPo0UELM41Vlq2Zl2jcO1oxT4CuG6gW5d9XMbnW/LUE8r40t7ws
PRTCdqf0wX8hzZv7Wb8jNCs6ndnfNzBY/nCQ8RifF21hQOJb12rR8VgYOwdpxblCqm8d6FumKGS3
SlHsZi64OSIfx2hX9UiXzBHYRpRE1K6f51fHcaa5wEiwZpkCG5bVZM3TWomwfzxMwJMa6JfC2k96
5HcDuYyjte2A4dHYtajDbCVIKH5Uy5n5EqkRcjCdTzmmrbFluOrdY0YqZNUHx8zNbXbbMwHezgj3
FTN+ykXWbvFQT53GGqKT2F0MKqgJtKOIzb8cZxxQ7LYP4LnU9rSr7GtXy+7UJxdQbYJFmbHeiLwx
XxYUVQw3NiqmQDcsqJUDv8pCbhCyrunNgL2DtjHZZH2GsrX+rITJva8+tRtmSHqJ5XC2B3mcM6mD
hintAzxyfa0VUfYDJdPnsD9TfvhsPJXCTrBJzs1sxkivhJz0K4OOJy281a805EQuoqbqVdy7/nvn
K182ysiBXcvSsmbV4xOQ8/JORM4h+6PktdwJ9MejFYWn1fN2nOiPUBvgium3PZn4zEQ+NQ7ETalb
VHtd/augHb3PpY3OaOccLUkMp2tmXVCN+V1GtdYKan5FsSseV2E360kx+As4cpn31a+Xi2vkAxGa
+RuNAZ3X+Ry5UJ63P9UmyCJ6e2eCV+D4ZxhuAvhPs2kUXis1z4meY9V5xyCHCdvEuaTE6sWl8rQ1
3IY4RbzcJSQgj/0r+12Gi2YSM+IHCbZWLP8HK+eMPhqzz2oHW+N/aJSvDPnkvLAGLXQaTSitSNhO
euCV8u7/zxz6oaxZ2nsZi2b4Qpj/LHSsB0LLNBKqeVZtLR6PiAeIGknMccH4k2/Kim1NiKo0h+Sw
vrKV7BS4slNUPZhHKn4On3LFL/bJFP1zy7heGkcGlif5/jhfe/DlEaaDp4c6Nfkx4432zdkUPYaS
Vw0ejNqupxCibiSUjG8jFGlLVch08wgbMxXDWbq2hCdrECL1KwJXI/ECz8THdcuT2LanugQtiEkB
kuEhKSXoz5efkmFqb4YwyInTc8BQtO8x71lQUqE30mtW7J7E3xpk5YdwNxxhrUrilyIEz2xyRst1
4T40LQE59ln81JV1TknmTTubCrLunbQv0+owJ5ayUfFyTN05dcmkA2SFkKQe2JXftL2i6K5JfT6E
qdXYmUvBtYsLhM7xUB3H3h4tMLePP4v/Ys3+BwDfDKNyQOQ4WwkgW48lrAlEmk0+SnvpQUIXVj+W
iyPCQes36pMyYBvHPxdmNuVk5DpFoWBpU2cDeUzDGq05qpQWsHK1ipus8kMY4AOV1sfbnu1A37nR
GKMN1zHrS4bEbfE+CyAF6mndQ7RIVzA9utv3rVg+cACmqr5lqrA80sjYTInuE3IEiaqH99UpFv3H
roZKjfulv+xY1qlnJGpQ4D734LO0LNA9/Znv8hM35F9mVDd7B53nULxmY2Bwfw0rgWiuRhw2CJlN
PSYB3AZZyOwy0zi5mqK7pH7BweGUWdJOpfh5gRd9bEPAcbs3hfCaSTWQZhv5urXuR5bmHWORMw8D
zWXCVYs8jyhdylCASl34CBtUwG1eeBky4PVN6iNEG4fUph1uoxgrux7I7wd41MSZ0HmsHHBPCI5h
dc3bp9DoF/6Bi+bRARdYLk3bQLTH4chlAtDFbxVMAQ+oHNIzIV+XAWjM3/moJ0KH1nXie+9HlJi/
e27O5cO6eLTeLIOzliTgviD7MiPC/bysl9cihzVaucMuRV1jOS7Y7bfPxU/FYQAjZ5cfIyolYqDE
aqNlCwzqviFHs6X4zVkUmHRMqNwbTqXPE7vLqso0lp3CtMc0zrKPCiKVChZ4xBPV13+yD+62UV2S
WpE5ijzpR2/wSZkmkzx6asyAIjCe+o0Gi/8M9tHMKAPWTooepw8XekubL2msLOIDq1Goly4fFVtw
c2F2sAUWqtofomvV5jjmChl7zdqyYmoUkiL202BCoczJy3UpJY2GrAIypb0xXrYWjKQ7yAH98Hq0
FsnF3ppQslHAZsFEteOP1n/09GQBvQWs96Q3dORZ5kNEFnKy2A46w6NvsEl0DYCPsJLez96bQ13+
Gergu7jmtSd9d6scQv/VQj8xs6KePUvex/arpfS1TkMs7Gwf3CxaG7j/01XExpRBrK4+bi1IyC2N
pV/yoRvP6wV7gWRn0zqWE/lE/EsR5CRvkDjzIop6SNn5om/NmeYO9J3a4GaHQ/AjtMW9EecJq17w
YpKVGJ7mVrWmUScgcZD4NLG8wTGSeKi+vSRLGb52wp0oV4bTqQ2eL+qrfFirGXnUCEuGaS9SnZS1
jQkZQ+wbqAVEk8DUxfv972NwIdZuhzuAz/6qwDf4F49JGd95dl3GJxg0J5Caz6a5kRtR0iBnlW1g
rNUElz0ZcfpheTXj+Yj7DQqI7P06rRWJsD5vGm2ZIeknv35IniXdWTvEnLHckDUOHTw9fVrFX2d3
tIHT/SsRhTuPJaxQmAb+hjxSCpE63SO6FJ5alLpmMTc0UaY153tXGuCoSM+0DH/6mJqJXkLixGrB
yXkpbuqz8f8OL/PCTrfLizVnbnCm7lz7W4CEMqrlRVGs9mdUvn0dqvx2eQJjUd4FMSBhbF0sSWPL
72Oy9urbwOrMQIOhdomBVrbuOiTiiVHq/H5o50D+0+DsShD39AlxU/xbdh8BJbo34gs7tapu0mNg
xcOyfjZIlGuyffOPcdaUghTsfcdA48xxM7Y6qWwP7/4OctuMPc0k4ostTbSeoKKFVXtq+l3h9DiC
Qg+UCumJ8LrANuXjIzEeeaVUJS+8fbyViEw6LGvT6UqJdDrVi9AaRI3LQOj/aTpnlMQB6HjhG7pG
UJCwssaxy+HkFjcM2dGhXy9ZnOSCUvqDTEEihp1eTSGUHl3kZpZWTT4hlpVFBY+CSFZpw/poMmBc
JSOKx7svdT+trv8/WLjKr7tYo+8WJMe1fwEZdwCaXFOIuNyQokAqMehQI7gqPzy1a82rc8CugDpU
egpzP5M89+wfTWP01QCHH+nQtSZ9vZejd9FtK0qC1BtRViOHPMa9PM/MTL9Ae/J8JRMd/uVTGr3M
ZwKDO3bmXSbbEzYOQuZDVlHaGlGKcCy/HxxOZl2H2ej701Ilw5/wlNIWGdq6LBvc+EiCcLK7iK6S
W/JwaaXYt9TX+avo/As2Ua6FoBRLVeJgsWGbz5LJXxVVl35KY338ExGjRtgAdJtbs9sH6pHN0Jb3
7RLGi01sB2l62tfpMc1uMT8OgNm1nvDpx7LdYhvKI9tSa5rgmuIYUaRLPA1M38le0jaycXjIdO+I
RonnJ42eQVbQTvL+Xhsxh8OAUUlgPWpEzO80Rqcjk8tLjFeKBsF4fxKXEQu/WOsqO/dBozVHl6Hu
OanR0KIS4JKYfhU4bQZ405KnaSZbPLNhI7zqKc7MguFUlVJkcJ2NYvjTB72veRkC/depnSND/S2l
Oi/JyV1+TUsccJ7g2JbQlUDGu2yr+lB9NOWgA7L1zE0SHh4TOfiaI68kaYyVWTzcJI2yleWUS5WF
bpKslBbymbwrB2PfDF6W6ErHuBJH7MPreDRXDii95SFWbBmSPD9ter150yp40LN/HQexNDWL5cp6
u+CTTGOvN9LM2bWFTDWcS8axiUhWH8OhUc2TcKZuH9vmqZKO/ZK0whFjVLUe53r/t2AOr8ZZaT9r
uW0oyVp7DoPEJoPHoe3uqnpbmv4Titd45WR767y8LogSWnCmwQ7sRwPzMEAeo5z147WkDNSDZfxH
roB6FiwRStZmwZbFv9NdmRk8m0n5iFJryzPdvae3t+BsaQlNQxAZDbzpMVfZTM5oqBYaWPneRSxv
lu2flZ1GjisDDkSlXRr/Hua3gPMPDCWW6gjTahTkg7Lz+bMEH+dP01FTusCmKu4pok8upb3GPejE
RLw4JxTxLHI8JPN5jjSGa6jfT6Cl9LjUX666nciDPkwrQb1qlAyurLHADZRzA322ZjlI/MY44maE
8YGy/Ck3pvEBmeBTduJFfTv8J1DtMN4gYq6UacUDk6B6RPumClUhxkGtI051C3noMHee20oqNkA0
3B0M7OIqkIVwVldXZ28A2JVdhovCBx3ZSLDN6fTUtgAqh00lcfDrYNwt7jsxe6U3z5X0jzpVYNVp
TCm5fBNKBhOYYhlBT3gYWozkchZJk1VP5zqWpSIXF58kSWXF91Jc2lj2NQvtIgeX5kpKjwaNKpMo
E89/VWdrCamRNZVSw3tiPd6DqTM37AZwtBEN7VsZoYvF8DEq8Qz1xxqiwr7AwZZSDWApSBQ698wa
SmO6PczknIPcRSNUFzeu7fFFxk2tYlVG90kNZO7cQTNn20pRWLaiavYhinCoEbhUGprkwpuEf9ZZ
AF2ho3vLYZgX9KHXAAc0LIGDCo023DuO/pAoFUTcCYdmptGQ+8PHS353I1FZgY+MtkkFIaEYZzSP
RJsbFWAtGYz0do0o1Ct/S1rfZRqI6ZaadLpy77Qr0aM8fiJD/c2qSvnOIPTusItMJWAz7JjKEhE8
FUNFWknaRRMl7XVcSkcvIHluGhdcNe50rGIHMOkbcLBFewEGz3PIw247HumXT4WbbvcpzRY8OM6U
oMfpoBNNB6qXqwcvnF8x5z/qd8VS0xn8UeWCIlNYXQ/08NuKCO5B2He+pSdYoBGXuHKDR9TwkxQT
c8cvKRvg2oPGoAL+T3hBe4Ef1mQyeHcZt7N5H0d9/02m16Kn/aOOThWZlM/JTVHYvttC1vsvCkXV
cqjZ+83FrlBSuMJiWHFRVIAeZf5JcfEPl5SaFpyQASnHrXS3ypOOpBhaHCHDGaPNw5RHspqIkzSK
Y09nUqAX05AZC47bU0iPewYTP1MxhrXZDFka7dq+EHwLhAHTE+Tdt1hk4FlWl+wwkaSiJ95A5UXs
3po7dBKczXmg6azxiltNSq7CNWfj274JHswU4QAzQvkigjseD+rX5mbUh7yVrEwGdTa0Qx6NIDZb
mAdjfjsM4hpaB+CsNQCbxjnh/9xJ8GtVzRBoE7aLO4YimeavQXOgXgjfOgNpUG+37XFlThSheZEy
qt4839PhST8kt8gu8O8KrlHbLQIz2sn3w+AES34PA7Nxv7ebN5pU6/Ucv0qaK+HB1g5IjnW5hDIn
YcPpJ7ZTBTjKJDIrUoP5su0oqVl0eh26Ogt1XdZekaRavhlzGiotcZrTiiis9nWoCAtM1R3wBbBS
X6dIFNppDqRR+N7/pOJT5zbi1/8nF8jgy1Lbr4RwZcI0Hgwl8pLNz1G/T3bG2Z5kAoKXd28FnJdg
lsw9JCUJ+tCIx3ubGuf8BrxbIQSf1oS8w6qylMDUUfcu82TcZJr+56J0XKGeGqSCERTr29F2AMcz
0stoRBJzuIK/nrOqReiMLJCNCNMG//wXGUKJUi6AYvETyh4A09RXwOdrMyxKhSA2VmIfgPwBQTlk
u4KmBlO9nEcDOpB8vIaDwjkZuIp8jOh9zTXQ3fGoxo2LVSDtYa8ai0o6qQepmpX2u/2lzptV07pW
2OXUwdjA0dctwAOGaPKsMnYwU9rfSTJwgC/+yeqceflcpErFtsitHY4NPcSizCbIX+7CCwqLOLXj
s3U5WZQ9HKbN7BjwS/wJuVyCnb08KJ1HVma2/YVEUd4rZ22dTRMSZH/OYHB4CAOGao+OePzhjnzN
0T1H/bBdT3gpi2PKBJTVSPpuLiHNySMM0UTCkkaH6eOo+/G28Ip6j8GRkoyuuSux3f14b7+xrm9V
I50gu9fFzS01qyQ9/GBTZiHjq4TO8Pg0Xokd5ASp6e0LCz85BPTzrNLgbUl373XDes8Rh+Ahvt5R
decjhj3Nxb2LoFT4OuuFMdS1YOzj4jSj1XlrjNitOlr5GE3aja5jNyCOmOI9EUcz8hRwVBUwohf/
ZMQdYohA1GBpAKWT0nS552IVBh0mcjATsfDa87360nT2qkwkEjRalcA4e4duKoqrxQSzYExQO4c7
9bTTGQKj6XghH3jqYP+KVIe+2ZGZkc1XcVAL00DH7SoKxTeUFfZ+xPwPgOboZfTM+H7PJKM6a9xv
q57rudom0loZowVDfe6x7zRbmG26WLO37axvw07oud4ziVdVOd4YciVXh0FR6430iqbp9stBqKPe
r7Vb2a/dz7BLBTRl7lTMTDbOWnX0G5DkM5IA1uB63gQLW/YQnRQZCIeoqLEG30cvx1BZSAlCRepV
WuYM6FbOyH3IrrvTEFEqaLwbO+83/kB4wDMRssqXp3ZG+dSq1wxePFGkLTTnQwxl+Uz3GJJgbg02
1yxo7FepCN+b10WQbSWY/GHSvS0kheF07yNN/2lLp0AtS6GEV8VyH5V9Mvewr98vWefNq+x7CXle
DV3A8PGuQVopS0MkDyVbwuCLTWR6bCVQLmL5qc6GSeusInp1nsVnStzsFcpofXx8RD+RY1eAXtV2
QVSJej5yUSmigW/3lu2C2qScx95qHrVowExwCk1xcEP8QNgmQZUwMMp6HXYEl/M2Lfa7nTU2dmGh
rlkUgRw2daeOj7S+NDB7uMm16Y3VGrgDkv+PzTl+JsudTvOlVY0MJPiSCvNE2xpwRgo3+dON8iqc
GdvmFaJI0kTa82ZDH9qUDKkO23+KNjdfQdAoaf6nAWyIVLZsx//uczoLVGbb691rTyeK6VQ2WTl2
W5sCEqMULVnFBFG5D1sx/6ko/YoCnImBX32hmlgGLGKHhNMgUCcGeScqyJo7WUDqY0nlFXebong0
PKVhtxbk+TlNzgBj3sF96YgLINxuQF7X4ioykbsHH/UEpmN520X5p/dhbvj7vdceYRLAV0enzSUl
jZwoZfT7DFRQwLw15p93j66W4QvW8Je8UwD2fdqlfnaa9hnSmvJCSIRxHbHo710OomSYOJ0tn/9g
H/XcF6XewdhLmS7im6y42KxVOsZEIyx13EVZXRIHbQ6J6XeOGW43p3awGjc9estH7Cu2qOWgBVF7
ycdg533SC2lfJPI9QauCI5ftiv7Tkwcxs9P+cFUNw52YN7qz4bD2jeIXc+1lUKSwbi/Oj9gqGiOn
XlXO6cNyYmn9H9dLDfIXoH1wGwxaHoBklQmwnEX43en1L6oVe48BcnvkbPElVuByUPs4kdQC+V4N
iMZssDwaL1vQ0BGeiVGWTpiTsmxHxnnX+iDpZk764TAY+4/5ocqTzfvmPlgG8uIlGvKLV+pqUJxg
HFARoxisbvXuOXBHv5p1iz+EIPaKAq6s6D8MrKD07qZvwYL/eqEJte+Mfm/acLTzkLwovWqQqpvZ
NQK39yU4ptevnHxm8Mw5MemhTm9zIl9Ku0zKp9cRR8TzVj7/Jx9qS/VFodF/fi+YBXmoKNYbbcH/
Gz3VSC2GFZdEKmbnVxlviS20PNPPD8uxtOtURQEPakF965qA778hWYlHpe6skk0Tgwsz0sG4b2ov
P8V1of2BzMw7+3TJDxWdUOSASCVWOzZXhOAXC4zFsF18qRZFGhUHMpUC8dojxtTgTREMoZk0RZzj
xlFlcKOBJK+YRql/E5LbtQkd/7kX6oMZnb39iskgKwPCtZ5UiDR1vke95ttOxrFrIzzTvSNEcuvT
K3vHsTLOD8jXJ/Mw4DYvV1OLTxrCpH2ZkArJelSUMgJrLPhi2t4SkGvvGBc9PbI/ZzVMSbIAhmQ3
25s1ZyxT16ZfRLrdbOaXfYxrcqlGbmn0j5RUw7XChE+X1bmdobBm9znGF90twVUXKqrSID8gdkOS
exmH7OobFGefzj6eb5FsImBGnBH9rN/Obc3Lmkc3n8DVcM3Xn1Eedc1MbHjkDfP0uUbvJUkP4VLQ
uQQDmHG/WvwJwnUVTX6jQuQ72aI57AdEG/2wG1ujRCU3IPPTy1c5Y2k1woDln4YD1ikC5BGI6h0C
0quAOSQxh7V9ES338ftlKeLUgFvMNPXy2SyF5N9NQa62kI5UmttxviNxdxnvVLtHSsKmk3kTN2Ph
TJ8BFitKleEaJXTs5CboNDxNea9vu5MZKg8/NqHR7TUMBnd03XTE5D5Ivt223r0281+Kh9xqHbKH
3vonU7b3sAKMyMdTE0hHUaF9Ertaew25t/FSl1I9UgZNjwmVx5oVLGAG3zAGIJyVsTVXcwK/eYSi
ahNcYcXCYepILQTjewBon0VAV7AeMd07kMOsxJCQxW3Pooyrc1cDFcPncMtEXslGb+yylFZsnMTK
Xf1F2VlWATOicfJ+23bJWwaouYh5btldcesgOi6ELJknC1DPeV5dkED4Btr9u95tPMTrlk9QgTsR
cEyhzTJU/G0uirT8VrT9wKDnuxP1T4tJmb68elBpxpAcnIDj9Hmzg/9CacWfmRNz5I4MxYidK0vD
vLmC6cqrXSA0YWBXT9URTQ6Wghi/vMs4ISmMvrAw1Ato0jyXxatLuQghOxo0DgULvayGPa1xGqgL
C9fI9xDp30UZSTJhUKk90EWYNFfqps3mDlag8xCf6rbJvp/QNbkljV0xo49UFZFql7vfDw6ZvYgb
50sfTAXgD4GWzHeKpSuEWIxKli1fats3qm6bw5HcFYr1cu1do11aTkG3NZfkg9QDXL4pA6t8Hjpt
b8UR0WtLNWpqxlUJ97X0Hg6zIFQZ/32H6PSaLoltFPWAXYmR107hR9hZbCumVBhxbiU3TxAi+li9
JFSlzw05xKSCsk8RRSPVLwPO5q7Qb6ZbF/0AO8vrbUgv3Zt6DuBCCYi0L+rjkbxTeyy42C4+PKxj
V9xC5dNWKmfUHZgwhBPC5B19SU5TFHA5EYslj5WBImIb5VusyAVV9vMMZeJY8uAq3bedVZezVJmm
vwyN0AU0ualuHR7iCEBcsU/IDx61O6eAdassK+hb+9x1ldhozI14x5PWqXdz+CZjQ727SSaV92GF
9lOHLOyPqvKEoI+5zm1vttoulgM50/+ORLd55xOsTSDFmxNXe1q9QGRIK17Pdu+QF/ZpWr9gUgom
yapGrbWZQzGCXdsEsEhfc7wwnfXiKCS0tvBeqtVIj/VXM3dXEOU0CbGGXwmgwtfD6SsEQRJhvdv9
fgoTJVKBtOye0ElmLdUQNEsIPf2rXwvoREtGuSsQszwSqhCHw+Da+f2FFKCY280TkrEEoAfemrta
MUK9AmqVnTHjHQtHHOwCVqJfxbbBcMXhwddfQAE6Zfi9hKtPtd8nUQ5RMcnhvKQKAW33Y2BZK0lX
9xop3LDcdwHgYk9nYIxyM/nInH8YNpgwmXqFEKRda2IlziiJtg9Fi9VWGjqZeqE0Tgihr94QRouC
bBEtH3jT4vK8+MhChRwCkpW3mPuS8hVPc61+Vk4mAiFpCgyH7zj8pham44fioQY8fuO0SdqBrhSN
YBM9ZAb4fBvS8JqUezbf3xjmeU/4ajukvENFidTMPdCmN7w6RFBtLyM2xrWFB66TU+0uIL2ooUxM
EgZzrmlfJsc2RtVcwLb0jECwBYOdrmtS3EcguldQK8qH4baOCQsGJlXBc7NSonlJpo6VmeLt4X4q
jZjV2Ar5lQQq5u2zEiF8lZSWz9Bp7gIYASrAPtvxszvJdO6u55NU9J8Cd9jef6vrHIBF57ZZD+81
4QxdSzH4+tJJlcqRGi9X1atPZnSEbb7NmukYpWgW75i5QRTGFB9Z3mCQ8y2EGjwaQ3TvyIza6CON
ah1q6ny//Yfo85pxDEgA2ljMAiCmrNE9eZfn1fLcULhXPrBrZEcleJ9FoZ73yb3zC95Jk257jSVO
yqf5TRrhqcUROMOTCSrBPY7H5SFQKdBu0yWJWDiy3aAl8038zHVnm9vZKvi1Cs9nbs26RX/7Q0oc
d07Yq6FNRxqclh0Y5CCjpzsSVbdzseENOtM2VKDuF/wdLKEzwY+QI7/2fPGTLg0hhwuRiEhCIs06
2rKZcYsHHhjVOkUsH9bI3ygZlS/rEsotIJtNZ3g7UXL5/BBexAn7oZz1ZP6kXs80jeOplheNdGBK
7Cntb9JnyX/zLfNSVhl4zsNTxdiDds5vveiBbd+EGDt4ve62S54GM6KpM0qT16nQCSt7ULXuwfMU
U5AdCWAwpNYvTVLp5s1YSylUyiadRzu/6vx4BOwbDJ405d1q0rL+h1JmWvJ62HmyuXBRSuLgkrk0
3vAAg5e8Xt2XGOHeDwCdSWBpuicpREQdNEH01DjXNnUqqCfvdhSU4E73pzifco54nGQUkpRtKeIh
bL4n/ix/tYt9Ywfavbu60iZ2G8TVaIA86rhrz+76o1I5f7fnzwxNBIjAvD/IvjZ4S+654KxJLAca
JCS16tEQbYk5rR77J4kWKzLkiY7NHILUF18L8bfgRdtLZ0j4pdNm5bQhJhODMJbbkbfgznvAKkBc
m50NXGryVXCUMggl5SxFuRYKffFqXMRWhNUpLIIcB1X6OdSLtyEhiUCaKTjJAkoFUfmPqgAI/W7U
4fDnZoltRPx6c/G+KjNSsgryDVtQTtiBWudtO6IjNH91JHDJrMW7fO+JV3d4HWB6m/zTgc6a40h2
H740gwxIRXSMAyo8RK42ocL9gykaeFTq0+6TvcV47LCX34e6OaVzQt3++a7fEIgTxAJPuMcqxr82
JHsndyccRA+rt3FSG1LRLPALQSzuf4uh4De/ccy2M46YOYUpjwMP+E7yz7ihsFNf/RQdQNc9cbAG
gmFwemwAdjN9KSqR07CKfxiOD5DfBGdxNBFJOityusHu0pcV4xD1h82uwkkA7qSH+SkahoppvL/M
r7QX6ezT82+GuXNbaN/fjhF36V4ZdXThWwX1YDnzcV0hejL6p2zhJvKiwf3JJP6J6T0xP8RcPaaA
xHyxRpxNklQro2FT9MeXfdyaj/JZl5K7pBqzBO2Pmbg5RNH8fl9c9+f9j06f1hDO+t2EAAy+QzWk
h288Wva6HzlpjR6ZzzSG5oAtqEKG0HZFsTc4K/PRk5D0410k8N11ow3JbYQ1hvUA8lByxaJXtuvC
6au0JEEi1jOsXaMciMHHSGdWfkpE9LyZYURHlrl2eirI5SWAOyhVFQ9zPY/PPqbLkKW0tQwnSDZf
cwBEJRlz7lUkOyNF+zR/r+LID0RKMIQ9VJ0lqGlE7u1yINpYmDr9w9XAwmUOpJaNHFnjpQHsuaHK
G8n/3dHWKF/jsuYC345PHWv80cLu5F3syPL5+ppzydB8917RZZEWlTMp69BZauo/cU3rzB9PyNWs
Ku7YDrJUGXe64S9kQzUUVhepmpc751kp/YiKMYYuwWrw3DrEtbxX+DPLHO8beBD7NyRexiY0x1QL
I4Qb45JE4ReJjLIoHw47wLE3rQrKoQBY5kFCfZrTTkOVS/TDXZ6zlcP6c2Ca/pjPR+yY6iAy7/f6
qO6uFvD/mUGT6Cy9QE8yycwAtnd9YN4fevd1Knkr4CJBmARLPYMtxjdXRErPGICWPNAbsTs2A76z
aEFylEZIkjqVeyTIz/3HgI8l/4KAya+nfysI6wzRnrwqaTum63d7m9RZISoEfejeL5FZ/nxirUC+
K5tZpMoOLwrUBeHF5dHVd41Nso8Eq47Q8jRR++eSAnyjTRHXGNeIR5JNoBuoaC9b1mquklHelqI0
pGtAxvEMDINj9zN5dIMhsMh3kgmvlVmgYAaoK9dLfO0LgRS2PJdw/19qzRBtf2JcMrxDrpJTmGfk
wjgxbZ4KJJnzG8ItxPmKf9uxzEyot0z0Z2KKpz9B/Rpg3oxufhJXuV0jsHosg4Dsagp2azPOqm7L
WKti49cveupbDTYSK1jTyWoGmetxfvV3j0qa4Z47RO75sPggeFECVxbBXioUkLcDbNVnw8PbqUJd
JwGfqAD+KfVwj2uhg5KDKAhzhDusbiDWrDPacfvLrXEY11OPAScbIo7Ff3DNSZfeuA2mpZ09HPaS
E1B+CwUExsK3MGocnU+jHsZ+gH0VcP2ZDXHdGa1JLZqOYqdvbN64heGi/IWJmTa2HZvDii4/bsTn
3c8nTiTBTJzOiCmSKB/wVdAR4yyYKbFV13qQQWek6tGlMOypmhoZuc+QO7Q6Ul8vjJoAstqDzPYQ
tF3WZV2S63op7Mz9rhz4I9vTJpL+xcpGmtG1O38Oi3A+cdFswenBOPqkxW4/8DRqmJmWS952xpbq
eeeMKGI5QVZNpUCOZv8a5igI8S2zLSAqDpqJbbNfvp/il5wuxh4zhIXCY8Z2Jpxz2l/jZ5gl5EWX
DaCAU6+fOUTDxa4tnfLIfS2HRh52e9yB4RjXP+Oo3JyFu0iE4z5atMgmM96FlaRCBZQFE/twopZd
21IUIp66ajwVnZIuVao5oY0eOsMAmEsKFsKs2pFg7Uf7H76OkotttJ7a8/NgmujM6bE3wPa/X4oj
dU5PJh/zYUpXTckPdidw6XFDigEXFGB05BA9f9qkI3VGoFuts3SPqt/rEqWl/pobB20rbJWXZcf8
VKAiHxXLz+S6UqUjs3ohnZWOoA1R17emwuQXH3WYWEFhNS7DNDTTmD0tJatWUcFVJmzVXscwOIe8
5YnTmAY1vUEJFkPnaSCLhcan1pKF0bl4cyVD9GFUrcpnGxjSw7x95I08w5svB7WsfIay1BwjjMhF
ipHZhu6ZbEw1P9CBxM1NODCoKTvvYdAbup80QUK3TeQR/q9EuqzoO7j7LVhYZFN3ygX1vypJTm0j
vJ6fCu84mOz878N9699Ib+DdLz1uXw7AXvh2qYsUYS9Po4kQUoC+kT09AhBTVUt74jCueXznav1a
BdRVVzysgwMb0hDlE3qNOB5IRqAh0xKByj1JLaeafvAi7GzwgZ9HD06VvNpRUs6uZoN+AkhlKEgH
imQWSeg30cc6075Hs2fVqwd3kYgbiKWxG7oMoNRt1GPBMHVJiAAvA9OHhzSMjsqTibf9rVDf+zvD
rISgzo2a2mDelBtyLPfyA4JbNh3GBc+K6V4s4qdxOPEkT0OJtjH0jaBTN+tWZVQYo1D8F+Y2eynh
WjhTGxf5b86WEvSrOfzWN1GgVFQHFkAJichUPe3PL8bTtSy3NFwMb+utaoMGyVSbJI5WmtvgTmYc
npWGQfrtmOzrEc17T6ESMgi88WVuT6g5iLk9wsU/usV5x76i5Oj7sR7Ew/j68We7ZjCNiNhes2xC
hNNGDQ8IS0fAdFHJYMBXlUnhb1z9yrXef20cvdX5bnmNjtPyWcGh9lpPCWij8HgLm5uAsULZOoao
ujBlqz9lb3uI/glhUs5DqUWNiA7F/bYMS098PShrh0ecFAf2n/GTZNiX8qjpetnEf7jjUtidWz0Q
Y0XvWJuoTaVN+GHsEZ5StGGYIHvg786FHTODy6eLOacpP2+mEqBp4paf1h+CLACjYQhSLckVa+yp
PHdAxinT8hwfWThn3SD0C5hKEGFlflwZORaGWF+EtzlGg9D0NDWDMnU0u1A5QPDFlw98JbkXmg84
s/deN4VY32aviMQYIkP9mdTKiVlsfcwRrth+oNfLm9hfdv5pPFY2euFuU0CLUQ56LiGmDqugaYvq
Ot7hhoFTif6IeZcHoh/ObZKMerABkmcmknu3bfohQt/ivLBQog5lig/kBoU/GJ9aarL9KfOjFyp4
yYZL1A2VNPBNkzGJV2wsLT8fNyKoADBoGJg9jcnbWx4dFzVBe3OSeOmpGiaETgpvyYcng0TtYwjB
Upg4V/Yx+/QFPnJnqHPLsL0hZ1QecZPmAAhB9T9CBdt3u0fymfmWWQa4xYOT0qugWkjIAtN4HTEA
QIH/iChdepbp26o36BNgYmUYB1p9VlXiQcwFESzAZgywNxhlGWlu2JMcMMk6T636NXgVNJxLUxVA
+dADBAY7/XB3p/5kxZg4Dq49mSmcoZz+1RVQoth/HnqxxBJl/cJ2xywLd8+nClQATDHdKwKTcavC
N4Nm3RdMMLYHOwyuldIGt0Xw1HZxLHO1cjoJc2uJUmuz7JCmO7RCpj6vrjt+Y5086fyNEEpMALzb
+mZQg3xaPF+0BAy0ytrrzdFu+CWnI7tJgSygmIiHXEq0iKEpOAroN11BbYtxBJ0dP5ud9UFoI98L
d/BUPsOjnHl02jE/UtCHF3FErG56mWcO/x5P0G6+acwJ9GCVy6I5eIVLPjdDba/YPWyHnF4VIPai
1iK8Hec9EtrduZrBGOeOGm1StUuLjeVpdrAH8xrBG7k3ts3x3a75Qvw8lpaeg4DlXmkuDS405n4N
OGkMrh28hHIuqvbAgpNuvJZCd9BvJpzdz7N7p2tE+p4ZzBpClAU4YpE2Fs8reIarAlkhhfQ9KPpl
3kPTukpk2NOvnP26WtaeOl12X8Fgrh1mGB++etLTs7NAg/xegtEZF8vY9KuLc/vfpVKnyGcGrma7
WjCwk/IyHNUeQ5VthbSme1tVd1hBshGD/zyCTC7hENNx7aqP+WKx4xDpWgIVjXNYkPmioSe7ue3x
LgMq6R4gFDj47/bwDiFbFD4KKcCllj9sLj4/LGUrV9BIUf/9sTlojd0HpJRGlioAqgR695uso7aN
AsHTF+5cCpSu2EfNI4Bi2VvoIb8LusjMEgCLYjikt6naADFEcdbvbgN0KCenL9tqqj5iVZ8QCLLS
VDUyFXW55CL5q5apzy5YWDyCWtOBqrhsTlh5qIZ3pGp8JI8OLUbfpLu3tOBregRvS81JTM2eO9/K
FgrbEZ31uDh9U4Bhr0ZPPHLY4WMd14NTDDYOHMMJXCdr76RSoD2mO7Bs2NaX4f8pR5JkEIKnkT5Y
VYC7l8Uu0QsJaFB5yPrrzaI1QgtUZDsFoL8yA72KEziFH78ZgH2FMQfhmSsQDy1dhzQk2Fq4nSf/
Gf0wW80PvszyYZqip/IphHV7xMzaeaSs+6WSQ4kW9bCeVWqXuh1txcKycKrGvPNd8ECl8mNDJKeD
AwX92AIy+ygHmxei+9h/6zHomEatCLYiGg2pmi40d9zJHHG79GB/dd4J+2Lnj1RUbfAS2VGwlN5X
JlalycK+kjF+4+VRP944Uv7lEqppb+T/52Tx0v+qmPNie0vYUlG18CTcT7gSNIWBKmGHT5FyDfBM
lmj4Sb0sgkTLpnlY/rhTGTsgVkKBOKvE2gKud4khQNtTMG+4fzKJ8LbWE2afqA7fcHED+IrZStTN
anT0zWcMVb2M5v+qC+BdIgchWyj4VDPA6VJrkFJsritacgTfofYAcQSp4M9XHmL5j8ECA43sLCsO
7ju+fh9AeJaJRPGn/6/nJcsxkQJB5dh1staOJLW25uZMRnhoOrYw4HRPd40adHMhBiXEkrCcItCp
Gt50mlTm2aQDKjdogE7xnk9BbHb/m9yO83B9Q99jaHpeWCGP2+irlISmAob2bndU231NRg7bumWk
yKgGv84i0UQcvU7GYPeqRV3LdyY2gYNR/mUxirFWLXA8qBj/FT5TJbks0fDvWemNOUCIS/K5qZ7M
SV6KYqw4cKEE7UaIWqxnjIbtZQtvX3S5/7xVAhOHIFDHvPhZ/ueKqbKNueOGlOXWzXYBnGYqQa2e
1nNT68iMpQVBJYzRCwMrMk4MXMFlHv65zriD+ESVsMphDhyI/KwFssrmyRqGgZ5qrnHFok9eDZbq
MaVBHkWg4VfIQspJtcIpg8So0SY5OjE6SOdFh0bOAJmziOKEaYv+5yrAiBaEMq1FXuZdagRdWc/l
LT1UZdqFuzV2OnzXtYQeepEJRUDB/4dgzAVuOEI/nRxsjeN9MeDIqmmmwjjB8cnEqCqjnccsPlgR
MoXM+0JHy7oBighHDQHk7cWG1uzRnB+20kucLg+o4gmuT22/qUnVvzGr9XfoEl8UQRwmgQjLE8lK
5Ehi6dDL5rCzoRaZqlWHdaQwvcPPIGMvOieQKS01WwaoN4R+fpjTHOknlrgvExGXEBDnwSfyhmg7
D5ge6ryCr/iut5XLhqbKbdNFAF2vVz8pXdYE50IG/J3xRFROUMk1YkjSEzBRW8ywlYdCB9FS4UwC
HEReQigI77BDuHO/Q8Sxmb2YN1DoKBl6WlN/rMrI3bspmSE7GeVvkAS9IYOKen1jciogY2QWhnU4
qvgt446vxgXvrjPCqJZyeXFhJTkl5WJF3hir3JfQ30zP5kNTL3v5fUjTpJiv5PTLpo2OEqmR0Hkm
QhlN7ECYf+XO1c5nh/kFswhjpRRmDCzBK1AnNEOrMyJGs2mYm+YE33jpbhqK1CxuMCalEeD1fK0U
MKZpeMEUvbG8SiHfjxUxJONHp8jzYAOeNezlb1pl55OgRx0z7+94qL9KQKt9yyVv2R483jNQOmQf
dzjVy/CXEcsgEHifb3AupIX0JS/T3/XBINW80zRfiWMrWTLhdHk7cc8N9P6mwexajSqYmWZLPjQv
ohIo35Bd7qb2uXtDckVQamDB5qyWw0fHxhI5JpJzBrMr/JsJ+EUcVVa17IJZrR8To2zea+BgeCbq
osfafTs8AZBapyIHrM6UuCX76rBLwt4GXKIZCmG2hK3MSkumZEqG/pV9iApQKL2AJNarzsQSPKpy
4LE/WIlHp68xwcA7OIyUPTQn8e7oN+Ktili3TixRRpjUlUB38ixvRV038LCficA5R3NIhoZYy3/O
5aRB8YNACiB8fRpx1Ihn4kxPthocrcbzwNdyvWgLHITI5g4V1XOE4L/yweIOUAKXBQVXjAWKr5Et
MlVU/le2bJfaSMZHLwyoVt13RAB8a2WmRZgkJSeDBfCiV0IzqX5I/dY8twxMRu+ZZGoCcAHCXsVd
yJGJfdStQg11/gsmHjt4n9qZ9M7i3nTPyygPVfDgfK4nYXBLZNsx0/o7/fSvei7cRpIKRFGeLY7k
FCxPdTLeT772BpXC7/5yK79TNi2fLiRo1oTD26vOuXtjCSTcAVvxAG+rVaD+MLqgZdFms5Q653nB
/l4dTziu2vU5E7Ov2H+Zq1zKyZswRFMBfJLscyIqFiIyEuqV5KZ6b8SxGuSRCmR04bozpJNKvt8x
+cwc4rQq5unRP/4PAKY/ZtIUkj8PMtzb51bqa0iWDb+elOFEjeKg1kSNiB+faq/1/exgA1eefDdk
qPpkMIRPfp/fiX+WSwfRnnh9UzHqhdgxEjQomiBVBIbVKp1QAalgLsy+6khNGhz+C0sSgL6k2wBO
gjYkIk4G/BJ3Jqfd01LGqIj7TK0kEjp8LhR4TrcHn6lmv955P4kNTd8ErlXJJF4JA9YSxKkeuO3W
YuvxsrEHIx3+jTSdbf2TvISbih2zBBQNncpKGgeRA6aOWlJxJi4D9nKXvO8ZnW13Y0icAesZmbCY
0UG2UFJ/CiBMD/mN3IgboW7/zhVfCgD5umBjAV8Lt651zZ3kyZEXvrissvlvR7znON+Pc6mhscyI
CLFP2FxLGUbrO4iMHFabyvpYmdGlxaabmWrx6QAGBn2VP+1ZzGxZt/Nh0JVhj4ty4kHqb2BwSvPh
l8S+lELnx4ApKTLlz8QBqDBkcSSdRH4fvc4y3hHGTwNB5ky5QcSdnoKaaG81kEn3DWPyaGc1TxfT
+dwX7+K0gPEZpKdefvDKK+VRPifa+SOTV/4vUqeAOQGv5QIrp9T1WQedMIPrkvmcdo6W4QMNxVbQ
lyjaji+6ylrPeKr6qfSS+dJJKwhXbdmmr21By4ANA3PSCCM0rrRV9xZc6hGpWmaUmjASNUneTbXK
DSeiDysQIaL/j/1HAlKugITqhe79UvnlNDRqNLWgN8hIw5t4dAknRwoYpGt/g5t4lsbrweKjaJtO
fd7XoVXk4ErSAGV5jdOL89dvg+tSiuay4fR6BI3e2X8Hfy5t4cz9PxMfJAg01rRUAYoc/fMrSytW
IA6OzxmyYRfkxfa0t+4w26anlVZqGjWfK8hoFENbi9OZkSqqYAWEnPM9ppo80omo0o4PalfSPYJD
HxeQfjo6iOyScNKbEna7sT+tPbn5jbBGcYQx7yZa1WU/tzNNMWUBYMFoTlHeVSUi4B5GbUwbHsMt
oB5FPoJf6uNZ8382Z6BJYR1PGtHGmPWf7pUG4RzjzYoe0nrgzJGOaxikepDSFEWIzYV//LrYhwsE
KbwTFQA06xCeSdmOQTPBFUKelC55xShGMVMQiueC53BQYgv0TYvnvk430Uus4mSmsEKGriWdB1sU
sKu1T0D0D8toGJMy3IhbOnWfkeZDF3sFG+z81Rhosv9SINF5SAp+W44Z+MAuwqnF2s+oeTrzBIAL
3UNrAI6MgIkk9AsU0VS5cGr0F7YodgGyG/uDBkqlAFRMPC1sljdWVwKDKdavUX0xKi2f0mnKoYW/
d2iqeqz2oEYBcZ1Ed7Pk17J6Ui2EKwP7dci/4g82bBobkx3v5S7CS0FMvsxHozOY1ZqjHW87yCAn
z8ZoFC80uDka7yj0955Z4YJYTh0yo+9NWdacduiSJaz7TRhFfXIeZ2rdkB5RcgOyDWvc5QJhfbRv
Na74TTdGc6UbX4e/f+M20xLu77gBVUrzbr0psajj3PW7Nj8788u27DhKI+512Jou3y+8owLqErMw
+qF+u0oKvXMMe/QxL7AdITLUVo322za+/v6a9mK/gRJDn4/ctpUxMx/P0SBzO5wg23udOJjo2+jm
FfHwPi//8cjXJjc0WtrEV8NhQWfR9U8WY4mBMKzuwvw0SVQuDM1v2qKcLLiZBgi//dmfEKSMPmkz
fghBAQOAWJpqHZ+1BU/SJ2QVBYkbJJqG3joGNzRfasrgnG/C5ge4uwWs6N42kCA/p+5saNZWxyi8
jSY7iGibLjvvdxMNugt4ZRbiHfCWirgKL3cly6soVhw5QtO0HAA7XcJuchbxpfB3wv5ANYjVi2JL
5+bGoDj8G9JKPYYENinOiJhRAclHswz1729sqNJGRjMV0EPMfVL0MvvXtgGt2pFGWGV8ncwqdOYN
jl9LpscEy5VlozHfetUteOCUOk47iMEEqRLbGYTB38y6H2Y9fLVK7r5Ik5j96EYotCi3r7HzbZTq
8Vyb9lCIt51MDyBGBLk7GAVm3YeN7nUFfJ+VBOwalI2KUuKGfhA+lwQIe4tRwoocBf8/FIv83PeQ
+Qgmn5Gn2ebrIc1NgU70fg9rbsAeMWbiLRdBcZCWFpdKsOxHebSqO9ggVhd7K+5fUPPL5gxyBmsS
ALgSOd85wnIfagem6mwpqNXjzYPh3ItYfxRtsBZZ3UgOtuUqDfP9SuDgWD8hzNJ1JkMPfqGgDK2n
pbTQt3+j5hmftf/1hhJ6q05RfqGh5NIHHGtHqwzHqen4UAgugPgialyKvayIMkJmxHp55IAp1P+U
zVvt/OxDLJu+csA4/TDPJ0zKSLQRSKr0n8xzvJpYLZGvLZyPa30kK8BZxgJV4N25dlKyPiT4PJTE
LU3kT23DWepi1j3pxnfIh2jvLh5qXwR7PV0K6Im4J3GGvU/tfXdH97L36AfTZL5jXOplYzW5HTWS
pMnCWsuzXHrL6NLxf071A0Kb6a7YwSbS24VceYE33JmQ2hJtptrZ/Lt400jkzukBewMInxFTU0Ef
pxbN+3If9hkZmFt/2k+FHsOokG0iMKTQIgASGeL3BKsBDy5e8nyufTkshXH4qdygHDNOt/RtdXCC
MWUu+KbeqexDE2N7NyvEP9XQMiy75jWZ98GDNX2yxDMduzuhYD5E2AcSRJ39uCy4yzm3kAlPkW2A
bExHsZXGTDLa9XZASyOHzkyPxXFaePsmcc7pgMQoTe+fSIjFmC4PwG+Of0+wmHRweYckanNAb131
nNRUILI29/b7xrQn4pyz8URETSlrGNnOxDbENIR0o4YmeHquIJe4OZ3CdfynhKVVLgtQMDqbDk2i
ien/4scl9mKl9VDo3Yvo+4sN1GwiqQcWY4h+zYi4qbkSxG5aNU9SxXhyaxkIVxTzz5KKvRXebmdV
Lo+gt7yNNaEs2lpgAKCKXOlZ7xWSl9/PrpE4UN+4Ii+bTU7x1ntcYskOhhtSpX7b+pC5wUfYjOL3
gTbVG6AF+Tlatfh4N0JS2Q3JfsopWzfASBtI88KH27Y10gICYtCvsYhtzwmnl/tcsnZjzGSenKAP
i4578GUXjl8I08do3nmO5FV7kCecgyexK/9Pr8IfvpUciIv/SVHyE15G8BZXb56JyZUyHyBqYodi
Zu+FCWTJ3PhkamoGdncRzrpo20V1Jcr/jKd9Abyqj3r7Qf2KQqYO00LFsesvHZT6ItH+P0vSZLjw
mlqhfaB46ZKIcfYGpA9FTy9yQA+VME0JWrsljSnduhlkQHNjbSFmGgD/ekcrtPVSROgmXTCDoMyw
oNcsL4xSyVqqUZcSHwTVLiR45Ihry7QuLJK1H7F2NARLtJhAdkQ6/+mj9HYPsNU903UdaWTUk2JJ
tgCIMlwbS1YyI94trVNPz1SIGomYHtzcViDY4VJz7/kTaT+/abo92IpLCpYhQXVP2GTVKnwW7xdw
yWyRyBxt1HQJIvJx2IUZKLpUX5gVPWjdPRXolH7ZN5n1OrcoznyggvzgYLsEPtm3sMiukOoF+ClY
HlNoWsTpJz/XV12TF49WzcniTX98N7APIYy7UewpzvkdEVCy95Xuw2rGC7ru+rOOb71e22MJkUmQ
r1pR9dWnAwj+gzjmnVT1c8sAtSvamPIGdsDINDAnMxYjrTHomGiRqOZZft4Df/Nf5LjB1RMTKq3p
JHYd9V8D5DTHRBLVYYtIHKFS/ucMfRuMGoLYFwv+x9D1EtIY6Sj0BCqMmS6Ez1rgPXmPtIw0QV5q
BKx3aoMPzPv1lhqyb1MrLS9JI3RA+dynoT4Vo2W7hLFqKJWp3u3U4lN8tYZt4rpF0HIUij4S2Z6V
y0Z/Vdd3GCGv9HyXaw2jEvaSRmWbLvyzTRou9Bnc6JWys1Lpfau7h28JTfCNh7jMtQPmgDKjzwmy
+0TpRRYLX4GEA2Q1wDi4DaI6l9awLTpc9+e+PDdtPe8gpKofrHseO6JwripCytc+rSZn6akVu6nT
YkDBIYrF5qEsCl7kD26DTdinrNGbhjox5qu+mFh4tvgfTBg6G/xe3n8dkIjM5qQkoAcmj+TlN3cT
zFhQoUFRFMUS5rVDfcnlJ07NMvMd7Xv/UM11XwwS1axmhfTt16oEm9qvQkDJdtlO8tmhI3VizQnG
afw0qjPK07NSBRH3Ot8SYWSOsPFv/2vN5uglpbe1ViiugHPTfqzu9SXwj+IcChnAjOEZm3FsZDma
RXLGs7KGd2qiCPESJNmR3u3q9NH4n/jG6zHixGYb6H3JNGy0lacTNw7yf0zVnXSQFBJdKkHd8bfT
Hu1qn85ZmVI2HdrFaHz7K4wyQ1b+szVe2QTtTIcO3XfiAeNoTof/4pvec3gwYk0TiqPa7g72sPxJ
rEIVoVauZXPUv2HCIVjkdrX85es0PpcdBF7W5F93OIgLiOzEtZiBHJcSBkpn0JupPYIsGynRI/8l
MZCm5hnpF/ka/A4yntQkijkEw2laCTYo9BmUJrcfCm6z6sXodmgK4bTU8xRNIhN4d+5/odSo//11
r5y8Fwy+e+Ym4kAzPrcql0tdmySO6GWuA/vleilVZyku14Fxp52tKQD0ljqUWDTEeZvi9FjflYTp
dt3Wa905GwED/7vrb2eDFoVjpK43jVYuQXuzolQKE03tRxojcnS7+5AFI5WothEuH9YpPtfxaKDi
0Yf4cT8LzI41bfZGz9JMMWtoLsFUclaQ+faVn2EN38EHaQf5yKktO8Hjg+60SWuJvh1PMpTeifkP
KUzu8X8JlhZPaopYKT6tpGkLnHExYFA2AmAE/Br3cnV9ynlO98pKU6RotUmxiVUZl9XqHLDcSq3y
LzEBNs8vARd3N1XN/xJxKGXCTv5rxAdLSzXUs8P0V9xskmxyaS1QRs60OkqSCkD0SglRSivMhplU
ETUAfv3MbkKVQ27hqxuYo7Zg+Eq416LMZTfRBIYBuE3GOpTyTlO9XCKtT3XjmSTCb6bwukg/StFj
0guvvSK2+P7jgVz2RHeWUYfoK2g2bfXNwDsAD6wGCiKPXfLD450nKTJmGqoSGkhKFIQF44v40lLx
WFtsWoTytrOKnOcKNOsGGOYAqjlDaRvryipHLcZk5wXbehNhz9V3uExdX6WLuVtjIPcJapw9rf9T
it8ZPaZRH9fuGpPHIp+h4tNwDa82Q7FU/lbW3O0diyaPi0xV2ekmKvGXvnyxz4m2tMk8scWmgOgb
hFnrblNEr61YyoZtpUsopcxDiywKp+hoDa2MtoIx1V7FRq3b0fAxR2q41X2YTn6a4p7FFfsHsUVU
5BZfp+z0+GgwYKC/9tL0DM9A+wLB0WiCcIQMHjgPwcU2cKJfG1rOu9noGuZqkFq03M9wtCfJ5+St
CB9hfDUAbuQeCM8esq2TRi86XLvM4xAr7K5Ic3pvGSmit8Pl+tPhrccTKq9EEp0c00iGq4MVTpvA
fORXKGCYFxQg6IcJjq5Cju8vuZaW6YVbpjuMekB6vD7s969HjJZB69/MRRF9pOxiUTxLJV/eBjI2
BRGdOnekdaVtuKvj9KEWwr+kBvUys42zzp0zfzvU84Wq7+/JusfB2NsBXFzWGPH7+t3WN0Zo6uAB
z9uGsRL5VLOg7koSi1YovV2FRiO+o6oUZx4EqSHfBFOARdSjXL5S9WhVDiny0XGSP1g+cqo9jzU8
uNg4tR65r/BGBHk+h9RX06TGCaPYXQI0YLeTz3nbCj7NaGkqgp8SSnJe95QN4Un+TX69PRS9nycq
lSD0oEZHevNzd4BrONfuncE2quwDG9ag5gjvHTEx/evV/LZYXdKzDw88FkuynjQZQ9SNeLunKLym
+gu9zY3v2sjNNjwGWcd2a6xrGGdt1nqR6G/m/31AeqJwrAfSOViLz+SI4JYbbhyMXMMf25eiCsO5
cjkvnzhF+BgTJWV22c4oIyByI/AycIwhXf+c3tp6t6QZsVUqeJz859d/XNKe8QHAzpuSuf+CK20f
XdVrioKPj/0a7HePLupF5fwa3hbGgn4nQNItWvqsPeBnFp7DlSY7/dk7/ihOeCenpbG8PAMrutlQ
1A9LMeHfeyuKhqFtPMuI2BGB2CQgxlEyXyU0Gtly+RxHse74Y+r4hrhDqRAiciEQrzQ+MS1LdAZo
cMEGEFa9P2tpXIF5+6TgXHx6yODgQZ5Q5IZhiZjlyf0ZgAvYy2WInhpYDIWReBatF1m47Tf2/DsR
LigSk8YYypGCTEuCk5JHkd42unMf1J+JgQb4VxX9Y+0tnJn/1b9T5doN/lUvawPIuPJafHGm6rfR
Jn5dr73Vp1mFmMVd/sOJjbHad66oneZKyB21NxBSCxnaV0V/KsERJBnnYbbHHQOOb/SqnWyCdWKk
GjZOE5gNNXKVnS8nZvQHFzd4sJIN3THDl/BRL42g0nnIjiFrLuF9h+CsIgtimiimYqtGUSajFBT5
KnSNfqNxBMFSPDpKUlMNytXeW+w2bCsGnUqZtxzwxkXGJjoHy4h6jAEqbDH2cIwSvyUrg360Zm69
07obxRmS5s3Ny9kLg5k+MN/vt/Rr/ySz1er+ovBvbShtpKbyrC1ktVyNRdKzdF/kiIsDluZ2uz1o
X+pSf/nDtUgL1LUWJdgIqmRar+NCRLGjfbGyZnAwPorVBlPQkB+0QvfItDNdXpPbS7ZE8W/7UgFV
eK4e/G7v/1p2Lt4L8Leo9d776nwmMQOvA7qhrbh7sw5nDXO4yuJChTJ6mzC7CVmWSsbBcLOWt6BV
XxyyaPDGzhH/HQTo6ALWPO8lmZvxc36Y93uAp3UkvZcqxCLdgrdaUI9tMZ9LGjS+aeWkw+/cVMuQ
6xTk5bsv2dgSOykbhciR64/ImVrgchOUZkztbCfKpJzrJpeqBra77vrJcdcVbcg3XeUDHSgZJoAr
o2cIxXFvDwMwZoj5+fGizV4zmcH7Qvs/U5ujzxcsdwYoOIVtLZ1hBcPDpjo6+shO/Vy1EtsRJMQj
rwLWdGIkypcNOU0tU7ANVvSgOlMC98dSOMdK3nhkUlTar07P4/lURNPohqEPUuI7KjzApGv/3S4Y
8JqTpbntCpa7IZtrHAJAMjkqnUcy3FSUWI5RdEe+NyDzWkyU8hYdqlzdfZTtW995tLH03+PIbsta
izWU+PThiJv3hIp0qwGwisHB01OdnKLcjWmyejHnHB553aMii2WpbZDp75I2Li3l+bF4SLZ17HYx
0dgOTjGyVK6iL3jO52Z4Dai0IWJIcnDhBlwckah0D5ykJCTkqw6mRK0hkbIF+pB1s2TOukdfmmaS
vHX2rimFs350162bRm74MFPxY6PIt59MGO/ljAjjZkf1WXl73F5KYCpXu8IQPdaxA+JulgGoZFyv
ef/6BX5MjGnXsJ4204MkLWtp2f3ZNfqVflQpUg+LAYE4cGk9/AceDNQrSPUIZvoQQaq71dh/BrQ8
lYE82jHjV7znWKfv+U75EJOGnyVmZsu+s2D89dL+qbIkF/E6LCx+6mVT5K6IAwLqgoKZvULI4iNg
mqkhJz+CRJmZcFUosXtawUMhsbtxkUH2sgnXA6W4oY6tYRdFYRnjUnyFrGeG9nHQbZj+fErv8CIP
bknUTegyBL/4gn5/VEKZcyb/zhWTnXJKXBEEie7+nVvfDfFpv5zyUI6Jz/22YhkR1GQcCc8O894Y
UtONHHiWXtmZ6jaJ8Dtvq7pfnRTFSvmek/L0b4es/4tJGZrwbd39LYTDe0Jc59qkXbaO5A0JAyfm
KceiPP5lFg/Npa90q0TQUlH23xSdk1RSbhgPFWdLsg5DeD2/GBCk3Kxcjq76bq2ZT/hjgE/uDHWF
4JxUdXUj6TmL+MYOZf8xCRQywJixzj95gF7jfoxG1ZrkpNogFoDLHZZESXcFTSlXYJzTAQwN31H+
/ZIVVc8VrhcQrwnYE6jPObfOHmHCH7FuJkhl45H6d9Ku1avyOFF/TV+AEo3LtEm+Hr2XW9mEW/qZ
CA0Yeu7qspSGAnDO7DfHgtDei8JDi95X2ETrBUKPWMrJN+aSH6A5mHeneLDAQNjlMfzRDw1xm1ql
UhXPhPmSeH8c2THHRKni0pvahlagHBDX0lOb0zHr7TrtfWQWtc6mv3pryx22jlWnSMrWy3lXIoyW
zPHW1yVLQYUL5YWrJ4AgzjqIEkPlm41zgXRepJ1Kbz0YrkrZYxBFQIr2itcuGjdLVL+MmlmMb+qC
cWEtBimlXl7q61M4sTudAPBPTMoFGapW+IWd2XJBlMu8+u2icLBOKq0JieQptwrWqKWDpcmm3y1B
w8iVysxaKDD00/CAr+vOXcurWOEjXFRcCG9CmynNqk6gTI4+1BA3thM8QvPkr+TFUNFKzmTxNECY
Oma9ok7BJcoryv1ZzeJ6m3ITPFoXzXbZFDgZ7ya4FeDrsmnY85vBnCYlOTXtTnP2imlYphsrZNe1
4Zuso3tIxc49y5ub0F8kJuxJEGbkPHvSPlDkpt6bZfKlQtSKI0b2AYiF63XEhmzY2f8ucw74kMrt
uEcBtMMCytmYAeKfUuIr4DN5eHA0TXXwleeoKdYKBnO6RZUatndb8pEmM/uHJ7hGFJ9tKsFOc+Xr
M//a1FEOB7ddCz9dmQOtvPIycTUZDQDyHAuFpQijryGFc9a5lNqP8brU92NLnetQbfjnJQZO53c6
rdeaQv12cZT8nuneK4VxQdW3Ml5bwZHn293yBrrd5ZPerCjdqGogwT1QACmDkuvSxC7o6uUFTLNz
5qIapEQoIU6MSaUdh6is1m7wRriMSnv2IDcdznfofLDJS+4BCLmi9DoBHL6NItNAsWPlHK+mrfDy
uPKDVZVGwtAWqYX3PdB8zrtqfn8kPtZBZVc0oWNqJgJeHrorfuyQxQho6i8wWzh7Xb0+pkXGJgHT
CcIl96556tyJRKmZ0vPyxO3N8HsAdUJhW2C2cv9WBMKkh+dGmIW/UBOA2x2kEnYTp2KADMgxO1RD
jtMTW5e6x9aQcduOs2wQvlHkD72U37vhZetupNu/ZqNUdIp5oZRpev4ATERk8sRGP8ekioG+EQ4O
pOP5fdirEzsCDilNRYEeEEhQYCJkdPDdjfqX8vrmh55nFMdL1yKeCHdKEiaTl94IGa5Fcz7+eNfW
EMi15N8zifQb6jWbNVO+jGAG4sAptICuHk8xf/esUAhhXf9THrtqiOkxdM8a50axkM8DQjoT36M9
KVvHTffsXf5jZDXxoEWFB4ZdtFs8AiNKnZByx9wJCGbTfiQBdsJyGWN0JhAM+7+x3BUIRCMxzJpE
lXizY8d5L4E0Qt+qKWB1D7VZ18rUfT8GqQoqE3V6STdqxrLc8MS12pZUZmXzkyQ2zCblSYE2VdkX
tK8NwYJnbwQkMQjRDm4xVmY/SLsaBCtsMSbpyILqKFbs3WiYZCx6/slYzkjjtxSxzG0sdfViT1lk
Y/pAt39YesdE1xxXJkAg7ZQ3cVPKmNxKbwU/3u88yUrSpUZ6OgS1bhjilXe/wZzEWqHeqjxWfjdO
w7afunVm4YkaIb4gmeaQcSYnfCwIM1+ol59s3plRrprxvsOx4UIUruzwqM7rrcdJyxfFdvoRJ2Z4
x+ccu2rwZYEiwQHZAs/KnpGgrQaIEk9bkIRWwTRYCoSrKUgynoMEZq33kYjzzwtdkdH3ck09W2Sf
kmwMWhq2JVi4FrvZCei0kkRvgXw6aOnLU7oZu87cUwxIO9p2xxqPPiruI6Oq14cvBBZCJzVq8CGb
MjdB92rjKfEhBuC+hS6xDVkBzv/pUo43SkzsrssVRdPLlzaHg2OhTL+0YbX4MiiICoIVxx00A0iF
+B+VRWOt/7naJ4BFkSob06TPW3HRNr12KqcAg+JkZxtQ0a+S4jq42fFYd7V38asG/uMj37AHNVlr
Pf8/LT78DQWBDzncDZKVgBO6KC8gGWNWHt+hBKCRLz5BTtjEkyqDLni69anSM9dxhjJUkEJz7Sw5
mlfCknWbLb+PYiljPzdM5Fa2kCNV5J4hHgDkci/FSLLk1U01LVI9yj8Zs7qE89aL2YTvzeKIMuNb
ifWORRYGHhDtk85MDT+Up7FyylqmDeyT1V8MNt0S/eYagCgJ1XBWClbGoa4DQ47EU0ImEm5TJzQ8
Bp72y4DtS7Rl0326JGzeXvBAdhYafQK5oYru83Vc6R8HcJs05+DV68bqi+g1j9wK+26J5ZCkEdKD
+ab8lTf3AIlMMbTO3HghBKDgmM9tbk3OA3cf87BnUbVv7pYGDKlZyfflaSj3fz9v/YNwWCeU7SVc
EMMeAVsBqOrO2S5+nKqUJT678pXT2o2AwWD/5VatgMBW7alNgy5p3Md+rw4LLPSBgDQtRF0zGKQU
/3Po4Ees8co1gWiR7AqH4GB6d5IHBih7foeqoQNUSbU1/GhxV3VJX9f1Whr/h6Qp8j9Bb1nhp5Gc
VCxviq+9moPsC9pdHaIcymPz0DiFALFIjPtElyKWeSDxorvJvwIbhvVC4j1zZYPXuGvO8UuXLzvN
6aL1V36GXWL6geomxwYtJcS4xh8gBsoGtIDiM+gySh0DDy3JRjI2PsKiBz2Pl0f9G7kFaY9r/W32
iKlpTD1H1rCUypvNtfHsv+TRFkWJ/KFwCAMHxTr4zmdJvae9nFrMpPe8AoWwG/KAw0kCEUg3NCCq
GnYQo8aFO23xeSsI1P0MGxOgOsVjtpISPeETa4kvjo6nm4TaVmfZzdcO7OOogF/VYRac6yNNjYgv
YoLLWWWqND/8GEJ1g0t9mkvzTtyTvu6JmTv+JCarfJq6pQfPv1ECdUDGM1yplud83UCMXSIgVPHv
rGNC6SJHva/qoqpN/cjDScs7eqXoTaSepRJKMuYGzvFXMJc+S9Jy9ekyfxZnHCHJXEK4xuCMl9Xn
+pIjlLpCbowh1a/RSaUq1n19hiZszouNbc4rEUWNLyeGsddh4KELYGsAZ2NK5c+iIby6nVoA1gNR
Ds1dQOg7WcICbhBC7D3GE7DEsNBYibHg+Jjrg1/JaHIw0A12CF0ZdYFeKhuGXVoEbMo0/KLWOsA8
g3t8WVODHx4S435Uvnmh8JnTgl+i9Ic+3PXOqKH/i+k6dFsXVWU98k8wSBKB1iV2q+rT4Xp64L3Q
YtlmwIEWVjvxV8GLGyt7otOMIhwEmcDYn0YEbEx5l34liND13iw2E23hDRZGAK7zpYJBbXH6rJP+
Y3zjJnT7tav6ufIu/cmrYsuFO/7Ah1sxpl+vUlYVY+ak37z45hDHjO9PH9VxkkT/AMkTODthfMhP
aPXg7YbP1CXJLTKWfrm+2mcKf29TVVzWf/+/YpKD6Tkpf5ypsHKN7eiwukiABQzplZW0yebZpgfy
S/vWe8+/K8BGWTfw+isuTOWHm04k9mgqmpFY6Lide8F9kMMIsDlVUWpmKoeMcZYGoTWhdh5UiCyT
JWapCmb9gWJXshAqe8CgKzqz+ZKwYlOx915xCaA4vNreW0UczWBw+ujd1F8IXOInSNqymf+kPt2Z
iqde0wXb/gVZ0rbf3zO+m1O9R2fQ4vghRuHd/hF04OgY9MzyhjOALaTkdnHBtN+92h6IQYRB3L6F
35xasEdZHZ+0lR04hZsbwXI+mWbgec04jOG76ftt/VCHJS9/bcxNGMmimSO/x47YOcrIV3UbOXhi
TNlL/guOqJ2/696TGR87ydFeLaarEDMqu3zAiT7QKuqR1uEQYnqREykC9t00KkhZXytjba0fQ0Th
KqL5UTbdT9LMnUyH4solcehXAhlD2FyB/lGArPF/2bKs3dmJ5Ou+cWOLuGWA/dVB/mmqs9hRgplu
CclpJ43lIW5laSxQuf9bARYF5t0hUa+r87EDl4hoWIFhBevxg7ilMQhMiAdRrQ1Aia3AolSpVTj6
HFz8cD+qJdaE+VwlPguP9w4xyH0VO4fI6+mr7BsAAAtg96USPbu+SoVelo/sngeSYXL/cC4VCdA4
M/wA37uRgGqZb3UTVPZiF3aW2mCCPJMFoGkgQGRu4wpfgXl1W/HqJq3MArIHfnlFrc3jjvXDxI3/
fsbTpMS/SPWqtUV09wlSeIj69rAYf5GMzZ4RstLQuDzzVC21fcXA8N4lVKltJXOO47BcZTcD0nnW
E7uwmWfmluuxlxbb9jRCcDt9S+nYgEMBe3AO659vxUmCwFEgHpRO6FA8pSWIRc9rnqW/J1YhIzBS
1JjxeSaAcaCCb4R1kwHtQm998b7n8JpscgwKOCG871e5OQmrWm/gtImCTOy0WiZRmtXkywYTJTOa
bpNHaN7HLGVgymD3mthFjSdrXGc6cnU1xBwOretC3yP4B8ebhTMKWUseT63u+gXeS0IObP2eoiUZ
6WzoVgdNgrLZnStnjbkOzaN+itpNZ38iq0Cjq22tBS9sMN6nc30ipC8zplrorPO/P2/mCKGJGerm
Ta+JBPI/HYn4qS+4rhIKN70bxcR9C0I4kEIcBuX5pNKvDmeLFjmhQOXpv0a/QfAbymVtnX35ycdH
405fqkJtM9YXfH26slAULImLWV5DCNQmXgeaVJSuqK7j3OTfA68cBQTDjZtsKqqO76XgI0sw+C/2
TAJGyNObkc1vJDcAFdzOgxl3ymrY6+OkxsKh83O51vM3f6jMl9phyQGAFsp59duMaHX7yXvd3Abz
K7GjreKcdnJ4yB/1X5c4zwhGNR3jDAc79auJJbidGxGSvtEit3bW3Ckcxhm17dCdGCjSZUT9gGQG
/3g46iHEYPz38XiStWLX9IaFo4kJJKMPn4LxWoT49saxaL+nIIpCf2n1DJLAoFOyO7DwDB4BSG73
5P7ZejkZnj7lb+0xH1hX09kNLaOMzfhOguXKgg+yU1Mh4XD/ut+g93KYPDMcOJ3V+E0EAzDrDs6r
KRJSph9jXrAVbn51KeFObn0neUzakO/nBtYVbIEBLOdUfgcf7ALjlkYlSgyddVvJENza7mt87PP/
9IHDAuDvqNOqhxXuYyRB0TgdFAFwo42yqRUq6nhAUH7HSB4udJiO9yeYyvZw68DtxzMTV8wUjgE7
E3SJ51yxGC8lKQ8l4UdQit/zEzzItEWnTh/yLAwjt3og9F+pYvG4Zv10YDPYMeTwecG7vPY4qFLM
T3ae1knBIcKgIO4osVIJxFqPxvuKawXALmDKiKQ8UcR/d6c8BFcZtLZLPJzXak/bEd5gIsxrViqv
rk12m9LKmeg3bYiKNArIl7GzbGdAeWCJ0W1hTQkKeM4ogtKGddYPyPP1OkhC6Y/wESt2ozyFO76d
H2lWY6Bo1d7UEnlqmaDlsLV0hDqBnHF01DRiS8HkAl67Ut5ApLERo3nJ9NWsAZ6ndUUFjI15IdRr
F9QGbowjOv2H/adOODhTtuOr38pKosRa2ncTMrP50M0ysWv5lu/Tx6DnQpdes0oTEaYDIKkFFxOm
mVxMC+WK4iUKMLY0Sk5VmussFYE7VK2S+/+anL7c34oU+bjP2n6hU07WBUnh6l/XgOy0CWa8pROE
lxYDPnCvdXZJl85hyj2VHoN6a5yEvNquzuaZJ9edjxVMxuQ3S2fWDTYzu/dG4G6xhh7bCRpWZaSD
ava0j0lY8MaCJA8Tnb/YP4HSlr0mmf5GGLF3J7W2T8lC40w6joAoJLQNXb/us1zb4m/Ay5kjD0wT
fDJ8Q+njvlTLAok8VC5WtBt1ntyj3oaHdHPdhQDm9n4nLucXCqFFM5ZdtquZRfAUiWYE1cP8eJhj
GUGbM/aqBI4RWwBO60sBdVaEnMoCbKxMJ19hW0976unNDHfzB+QGUdxxHsHknVgGdo8HeKWXcJHs
HhJ6tC+YWsMWPrZlaZa/Jo7loYAItm1zZ3A5ih1wEJ9MulO+pNaTZY5kAcxcyVB9VXJe/lJMU/MF
GHa7qdwk9nDMXrKlDUJOPvgqFiDG7H0BYjHLE9j2xGqm6XekpZZcnutTkl1C/Z+LOl5vLGtJEQfh
MidZEgAIyyGveo9LLap8x/HBV3SL6bJ80FixIma8eMZKZHfhkUiMapSjxscyGFSRyp/mvdZYk5Lc
f677lDq20+QDpj5KRNWfqn3HDD9HxBaKumLijJPETvRwoi6NpJpzGOePhUrVvkaxsVI6LUf2feWR
guZg3iatyJcZzeHO/C7xwFRJL0hzXkGgRH+8p5cfvYOR/L9LojbqJA/VVKZNjA2eNIlj8dDGTP7t
REJpqaQjjn0YjYyCxCkizcl64x4mw8+X7ZdlMiPYHNS1Yfp/Nw88rQIs70psRDc/eQCNW4z0Dbj1
dCoN7IQVD7G5LN28rhE2seKliuwt+K2hi66wefyCFl+1RaJ4Y8g+tPs3e0BXHVi1h3xczCKTHjnf
nk83CcnQ4oM6VWJEagVC8VSCEyJKD20WPScBKr1EK6If0tHHRer+v+iaGrfrfdEpSSbGhGnvLEIf
WIXZJIQOM6Mf2obkvdWrhW8J0GRrYIyZ9ueHvzuJ9iSMLgJWEgwq4p4p3bLqTq+1XqzAIo53XKz4
ELZYcBwWl0qQ+O6+fbvZmuz7HlNHHx+kst1c1glZtGdyqCdBvslD+9z/n0X1n/Mv1bAJ+9d7UnHp
HRpBlDzrvPGq5aXwTKo+W+RuljWOOm7X33eIC31xa6RY9O/VEwJKPhJQ3m9skJnuTM4KSA4yCvzL
TpI68oadP7vzf1KtPIBfHu6N+0KXSw8sauiu0dqYHDGU2cRtCLF9jP39S9CPGwnrWk00r40+S8Go
duIuKQdU9LE3cL0SazPt8TCTqeQgZB+sFvGs+dM/2FcBprEHuMUMdtqRGIwAkAgj7ZMzPSbf3RNs
YfofJgjlUZ66GY9X88T8LUeDhHTK4MfPFSotYNP+bSNSnh8LccsoFXpz56xscEy/wdwUPWXhdBxP
sNgNqCKLZ7pOfIUOE+MA3O6KKTBk7clk43Ai2/a8AfvLjaOkrn2w87YJOS9mrbOTPKLpxHwIJWJT
BiVxNyB/gEU8d5Rhc1+UBpaLhXDPDqBK5YvqKXyW/ZF/HZFq8EttW/lt8sq4XFsGXxVTTrv8RjmD
yozAXA3dnDmd0zOn3eJI1nCyX8ZHSqIMyWwStSMbVmMtvsXHXyvd6E1d6VPPNAdp9IIG3dhaWrrT
dPaaLwrfFlIl8VXhp/ghquaQrF+BG+1qToj7I7TsIvabZxbrXeFJEv5jupWCFOq0tX0HT/DUj+Gt
sjGE/mRapiG15BkOXFla/9xQ9XxKu7wCuIaj4mQoUIRkZ/fAf4e2fCWHZoMJjjPv5DGlKv983BB/
b1jPeGVFRvUCZtkiilW2MIZjUOU/FezKeAWTUNkSn0C5tW5IanVKeHSNpL7oZkVilMFzUQ3y65KV
QYpRSoUi+/Q1ukIbUCiU4LXV86F2zuZnb+aNxRZ11Dbn5riDH4bQ+rrgBdrxzyIOyEyuUL2lDxUx
u01xE/zSwNcMkDCqyIY28YI/K4XRIWqaedtYuCSxxln0zvg9/Y/zDSBCPtDWE2Cgs9MqHiA2n2+T
BgYTPlzMOYfhZ4lpD3CVZHeVZF3PkNDp48yWLJM3hY84hX2RwXQ5yztEcsNUXurLWocpmHrQdTLZ
tsbB1gaUTaIswD3x83TJdxLiOwoLuqnt7UtV/Vn8hMM+mcJas80uDNqo6KiNZ0ixbKuSSeagichl
W9d8nsE5VsPBd0ZIurDn3DrY6TtsH1hwmn07YP8HdKvqj/N3olwkiWAkOb8cH3INGOiuUbRs9mjV
ZOXR2yYSXG2SsfIyexCFWxZZzs9Bg9XC9mIhQ6qQ1CTRwlZP1irXeMfLTb8POXuN3UsJcWSSxEoh
aDLIf5UqjjZT8AdbaIMQAPCnl064Ed/MkcDyiaYBsmxcl5I/xj6wflTtQR5WsILT3GBPkiXKe2CE
UG6OnoLulxSkX/zR7tQFQQZwOYKkkJlm288ie6yb0y8UuibpTXP9cPUK+J/dMEHck2NX4MBtPgP9
17YRglCsSO1iijK0RgFkYJgErJ3G4PJfH8uhTW+nZl7ZGUq2JgZJ2GKD+q0sDccKZTTCE4uwDcMO
H+Iy5/yT3KKjWDZQrBNsVrchPTH1jzD9UkXFD3wL3+Vr8S4FG05GUB9vV7QU51bNGnlBX9sQwbvD
9rwZ88NltxKbccEqHl77lJ/brgL7/3D7Yy1ofOWEHEjKtU/gJZvt/m3OQrOoYO7V2G288xQix/gF
EJ0cGgD+g8+MTTZF8uDaMuVe5ZLPBeqU5rYIZHuyrlA5OBlD1USZrBXdN2aFhUN5FMq/dUd3h+C+
6SrijoNKTXuBSMPt4Cf5ZXwWVmvChSauMMSxA/QdadRLWPyP2hGRlBL3jWzTFx1Lq8WTHskxqb5o
0v/BtblwqyXEe9F7FpvmtoDch+qQ7r8J/JNFuYxphZ/yzts2i7NIk8OkicTVIP9MXpGuQAWk1uSj
lq1Bf0rYUXj6Jok8mWyuXqDPFaLkJnP/atoF2bY69QsdpYM4NUGlfPeMKKd8GbvyZvPLt85x3ZdU
JbLN2hy5dFTgMQrUlbcndnGszJ2x+Ol268bX2XmSZMtJgGIChYJTU4C0+Qx17nS0lNiR3FU2nNkb
Vg+yNigF0k4Y55ejWoV9nxpAABxQj6bBoF9zi6eEBPnwAJal7BnusWtcMX/7SGq7N/d1pr3FwpSy
gQfeXtqmxQBlgB1xmFoOMSNK18ryQR3oT+NTy/aQa9XjUO2wbmTHK2tgJ522XSuaRv4jxyJ1KEFV
8AuonLlxNepGVgjiY4NMHetoc66o1bbiQo8PMgCdkDTHuno8ZOFCENB9YRDqTGApTErGGjMDaP8X
HquU1/VxqbQ8F3K8MY/jGkzcZC7p7l/gy8mN4fabsNyfZHA/+tGn7uVF9dGNJObh98fItskoURrF
PasdQf4KFuGpmSdvTQiJHt7v2Z4UAZB3CvWoKxOpLUJkxln37tSxTfRamxDXpXtbS7cLC0B4C4yR
YP9ZvDNYPiDgzkxUmL32flyo5TIZtvSwCzQjZg2b6L1HmKnFU/opI6B3TqfW0jCxbe5L1EdxC7VO
aVQoVfLv3jpmnjmvVVTR8uCWYFVuamGAZnDscYty7lmXzRsqi52sg6WN4zcSvPz3Tzc0jMGlSiwG
/0+txTa7Lo5Bd9KGNpT6W7dnUs87Wr7yGGwGmP34Mf3gNRwOLuPpi35j11ZlOO8TgwfpTzFu7M6E
4vc4WaxEsPa9p+q797UKFeBN01RAbF7tLQY3Y4Oj9PRB8jY+kCjC5bwKNkL0wROpDqAMkbnWFuY/
O7xaHHZRhlr4+byb7KIQHP5kyn+dNE4nDRj46PCIDZfnuQ3NPhE2F2QKvaIdvegmST+lJxvPTwbe
Yh+2X4b8vGC+UJIXVAVZGkr99u2T/nuT6yWmdNcgIO3ycgw5x62OgITshB4PO9t8FwIuOcfnX9Md
SxVClarqh7ZMqkvomE0zDKbyUVwbCiRg4hT1DLx13KBgZGjPph3p36B1n0einT5WjaE9xYD3Gffl
zRVSImrMSk3O2VLw7SY12zgy0z6MJMJ462FhBFkcJegN9P+5cWXqJ1cO7PuaKZ0jnJsCgPYh7oal
hlqE5V42RDda7s99GpTwyScqnE0np9yAgajl5MJAyjyR4o9dRsba9Ok7HeqXuNYO4zzxCpYLGO9R
shuQBbvrXmqV49HVztULHtRIlLdR2kUcei8QsJ68DwoxwYFzk9YJvUFROf8bzK2bfNyP8lKqpy5w
Nm5i+E0cxLGE8gWyv5Or4dIt8zpaNqMY+j98whM4U/5F0TCnifJAqh4bH0OaiCwWoAkpmKXwudoa
dlC6r/Yidj4TUqyCT5diNPqwFZSyizrn8bOddRFxx7+o4a0cY83LbVRARNHp4Cr6W9Mo36uh/x9g
/975DHV7sOkRnAi2X53Vm8dvT9wWizm+I+T/sDmH1oihAfqWdgPlGbm78LtpRz7CPfuKqrUZJ4cm
GYIjVDCuIUaNrTtg+K1903LMhtqob9hPEA02fddbykvIH2b9XflywHQKCzv1OooC78hRp/71C0kb
Huf/j175ZqHce+ItGtqnlKpP06HxAmVc5MIGH06jdThaiyv35GZAP+bhnwQbI3tfD4cxk5lGqKkb
HAO2/CAxqmcTtz63nqlG1W8HhJ7cPVo1tz8mr3vU+fOm2UXZqvoTtTgpUMCsbavtrSuJK2V70z4t
bB9rjETJE+xHIqvNQlciSgrccB5yz+mMcWEBsvBItysgSVFmwfjJQ+T57uKrdcfLejUwgE5iyg/F
eomqQwv61PUXpDdxdHcmh3Zo9uZ6a8aE8bJHN2O6acSwW6SlkLrpJb/Tzm5rsfPKS7x2NZZi5yXg
Y7ONGK1hqcNyns8KwPOWSvwfPclUIM4X08Xa/hfBUyR6xjC1QINqrZTZZFn1P3wlTQHIU4ruCFZ8
TdF6dGM64RfBlqRsr+UgZEv1tezzhUy6G4G604FmH6whqY4eKaaTgt1iGZB9Hlj+zyepPf60ln9G
uya9+aN/vdGxVbQ/UYIwnEtUPpBXRwJOd8Yhf/HHmc6d3ycV3xOPkzZRdreMmhMA73d4tJU4Fd2w
J4a6YKCosMh4/xedfvTT6Qe5vRrnx9Av4AOw4a0SDMh6yzoKL3qAzvpuJgMgQaSdnmf8NmUFjDob
s81l5IsSZ4G9YTWAQUko3yi/zU/XI2Cds6kNiVV2luPDRVvj37a20bhmCSMGDuZmZSbJybajEa2v
WF/FF+4eYNJ2WGG8QrbC7YB8RMyUACTMuQVGFmF9INDGdUJXFPFCphkVPyHRqQOQ1OFFyOnUaRxZ
L/4gJNgMs1WGln53NceWDeYWTfQMFDSSIhuaYliVRrN+sJDhj1J4JUa+PObca01T2yvLN8Gmwa/x
0YHhb4WHAUqshzzvSQCe+hvrA+YyY3Gm/s3Y6pCnwKMZJCEuQAcDeecWl1cOu0txkoH6BQygvjau
QodcITI3Zpfd+KGrTxdNJ0/mbzQdVai0ODUb1E8cWW5EG3eTk8SYfb0t9MdbvW2OgR5NcU+rvmBU
V9bFEZi0ZXSbpiZKRjSWiP+YTLnWmrNGF09g3w+qg1Uv7UcVVAENXfKC2nR+v49shPAE/PSA+aOb
H+iQxJzBsaDgI2F0AyoiMsXaTOg9chLjUhQrYbHDQiT0Tv9Mhqm4Mzg7cE2PkVABZGm/03crhXLw
GWyVJ6OQ+dhdUKy+d4K56e3c0RJ8k4waRY1RmyccDwJGPjOnLkalR5Y4pCTPSgC9NzAaJvZTEOcA
qCg0QFMrFDnaVjDll5mk2sZcWfgrf/xNnonBe94tsSDZo9dPSv54BcNdOTiNf2xkLqp0hHUN/VDr
In2+wm8j/23xhPzYmhPKQXYIwNvWfCPnilfxuCERjETigjf8uL+DJu3KxFZpDWlN5USsIfN8XkKL
H7iLS1wSC3mFUE//1wHGVKWTi76g1U3v247ixZrE2xN1w+e8+vbUd3vuq7mC3KPbcwuVbt1woiLG
tMN0RHrMywa4m6bjzT4S9ndI9eGaQocIUs7JcRoVUiwiDVZiSaBOJzzMkYeko1D915gOCx2swTHY
d9ld7SJL0NdTgNd74XaSWaJSLbFuPXOITd0DOTd+lTOrfUGBgkcxE45ZEevCUSJcBP4JhPrP7bVp
XrGhHZEuYQpVUJhStNdmDyOxDg3fz2JRApQuSZejW0DYPNJoVfPr77Da4MP44Y5E8wqS0q8YLWYY
67I3gCZ5rNAiPA8SEyyz7FjIA79n6D8dS9r2PiaoN6RTVoqVVnEjoCdOWSob5gdzSzkPhDbFozqb
Z8ssMT9wxF5ZLQyPS8kZH7gK4lomLVkq5cU5CoLjS1h3at/cSmCbWSM8dofwKn8WsPkkjlQddvtg
oaE3Q+Gug2O3hoD/sH/lCng+9XNj8WsTsOoOlNsIHJ6+craNu62yCZ4MnksJOiHvAPPYg2bXspxI
yBL84LBXckpUHFnlVM0zG6VHQpxAexT1F/qoz9bO39a7c+7iNALznZ8TKdnchMeqYoVuDXS6tDrF
vyQG/Gz33Vz+W9lZ/mkHmyPnjC1br0awgXeTmULc/plj3VR5scJcxoBXonRKVNvPC5UgyBpYUglP
J+OR052To1DFeY24sxctTSrXHW67bYzt9gOhyMGse0IGXwLq7X48MC9LoYwAs9Di/dMxZyUFYAly
6HnLfDE8Ee0pvfbS2kv1A8h41nDuuo15YNGGDU5GyyiGyqIVFz4DTWJ8qHsoTdR+sR/foAhIsfnu
M55N0cJupCBWUjAaGkAzYcWQ+vD8Gz/LSPvkN/yUJq6WrVTJ03vAPLbRi4ecX0MBvYWlOXOr4Hpv
yE7PBWF11fLmcbu2dB2TEUjOOdaly621d1rVsyKwKtsJhJh8PIVvEKh1WZr7LXx5UGmjIWkfWimz
mJac7KtBi+YsdmHad+ehUKk/P3v6vyOB1QWXnEzUdYBlJR8/xrrWLb2BTe+0SXv83/EJEupl1Uqz
ef8A1rZoE82Y1nH7TJ99sGVammJGH2HR6qnbv8wxYkfywmWz0RuTG1/thsD/NNfW08zcFk5RbJxU
TXeJ9ods0BoMbtvpgD9PtrgZBMYtbTWsba0udGmc1PCgxhodYkFm478zD5TRiT/GhTKpTV1DT7Ob
5/ABfXsWU+Bqv/oFOSRngSYfLA4AoppdRNFd4kI/WIiQo9qKaRymvGNtKyXLyBiYygLDiMJgIQoK
AmmP5rBFPqbiHTpxENg512XnOYHqt+dOk/6DmvTeIkTX5DrOpat45bQTWtfil0wcOiFONPvnnIap
4GCw76Qnpg6uq7vqubnQG+iwkzEIwCKaaODTf5laetKYYM8asaTsGWBQcgW+AunjqO6ybm7nPX2/
zDYUX+YbbHEi0tzS3IPEpCTsESmbaKLwU2xHkEyumXNwdoNzNT3bWp09ysnESioM+bKfY94HCteN
9N+gsBKVO5NHI9jDNags55UZhZw4Tw8XQ2QHu13tIfaP/Wii9rh0IMsmjSq/V+GDkNJu43GjpZRs
rhox49es0rI09cg8EJlmeIfzTNPr2IihtGRDYOPs4Z4sEoROnyrfFNwCh4cVApvfjnox8gcFRnKE
WzAb0lMXB+CLT+VLC+S/T6WzbHp6K0gYo92ENg77O+wc9NsY+MNpw3ILfQoFU9Z7T72KfCtvx85t
28YdZARBqxC2X+Unb9+Gpo5tkp3Ydj2hnVkuZpMNpxS5mBeHqK+CDvrQ4UjU2Z9retHjQ5Aw4y8j
dxqBigsRQsgL1zNEAFRvx6Tg2/Xc6w9KNRLHc++OKq4Z+y4/Z7FJB/llojZNa7uR3BiFqX8Ypp/B
cAx+uuEERc96u9js6EzlEny+9NvOHbbSv86WRhZbx6K+w+KP/By/QVCCU2wO4o1KgKz/29WX9p7V
JMFBPl2LwHZ/dmMjm7alownW11iOV6/AQqs1YSBV0jxq2qxCrWYNEH+ElGjK/KbT/HKba4oTs7JG
U2ja0BGWy8j1X40xk7vebbgBh6kdpJRbBPYYKk/nHzQDckg7gr1930ElTN3RbRRLkiOYLyYjEJGl
rghORXB0ctCmXufDrZyxUFZqOik0L+Fd36yI4KvyPVxLTUMzWOL6vUpEoJuBAJAEIfi029Ajrz7l
30duHIAECheqx4Xhibef/9OLQGOGkawZx8mf9hswij6/h2V2/tHtjkUEPyMdenApou+2cGjmIPXk
yI7azJaGuF66XsGIZCmWyiedLphTLTl8i2o9yVo3VjGApB0a+/XKOHsyboEB0CMyU8shnWsXUsZc
3LKSPpz8SlprDDpyKLCsM04KQNhkuZSkscVitB1m0SESjkyI8c4fkB3Xhkf50UvgjG1Y0x+rSB8m
OyA5p4SP1b0tWVgUQH8bRw2e6FhmC4JDpIqYzromjKK4rWGePo14xRtdgtzqxAjRFZeXkNMOxMBU
+5oFdXVCvMoHa90NrEgapYi4BCnD+A4eJkugsVfF6UL3K31Hn6gN7sEBvZEgQjaBnjLM2auv2TiH
Y9Sj2O38+u2Td/YycBhZBKgb9itisMgIfKH9nQJhQl6tF6w4KJebAmv4Kv8eWo9yRWC6H9VATvTq
YIN8qp00mz/0t3ov9EA/fKrnVmJZNkr3hiVzQtXI1S3iw8e15Kd3vmGnrBLQLEvQJ2IBXcBMXLOc
kCXXwu7KrNDZsDlfitdjQHHPSkviqXCQwZUfT4KLXHc7f+oawkMMN8ZEx4BVvz8aDgrfyVJHEJVr
A056UQQlcbdYH6SufMGprKzogsiKGBj9DGEQT8hj2AwCoN8kZDPm7DCMFRAxgs7D+RA3m08vVNSU
wsr0+DtwxdR9GlIKs6oZTmYRv1o2uSaOH5I0TlB8pk80tsBlx2kRFhCKQYWX5fej0EudEFbHkM2q
Z/fyw8S+OSWvb3pFBr9GyZTRuxE/Am2DVKadpea+pDoVlTY7DJPMbrDN3t4mBTyVTXB7rRqcLXs5
/wfMBhBi+tAUA/H7B9oGREgv4G1QB2j2Tpk0x1DPQSawGnDk6xvPIktQBJ6s3ZxNzlApB0Ylkkq6
lX3aUwnEweQ6ofTBasg0kAv1lHKolbCemMt2Ikq0Mg7zhnNzxgbHSku/MaIzUUVhxcOBrpopyno1
ZIpf+gRQBCBIo7WW5I8WPRHo7mG31S/BpliflVznIui9tXVA/O8EOFQ+IPBbLN3z3dpF6URtoajk
jTuKyaHMg8VNOi44yO7Hszs4MK0/gGJI+tH4N+XB5qBvykOxOskx/db4Bt+U1uNrfDC2zN5ZG2mh
YQ0h+Ydc9hPlM3A4GJrmLE3+7r0xA+odewlKJMcziDcHCLHj2psSBluZTLHs6EPX054EujQN/4XI
qZ6do7g2CgIi7NbeqSakmbbkO/ODi82qtdbB3Yrs8o3mxtFKDGRAQzH6VQErrZ+MUeGGc7KQ9MxL
QLQemB8LGui2XicQ9Y64Kd/gvhhxBXDcudwRWU5Dzc48JmzIzOTjwjcDnaoE70Hh23ttV5RvU+mK
8zoRDEQOC3SoJB48gGi/hndy7PovDIHoc2AeNMJ3PmHPSGPGoIdiPovWl9LlLZY4zHa8VCkaFVfI
7YL7uqAR3TuDDV5+Sr+guEQCuaHejF+Xe5UqZGVrtGCDMj4EJSu7fdZN6GC0RfQhHMmZy9o+XjtT
ck7/2F8DvpFE/hZGgupKG40igT/PYvfbbEpECCuIUUKqS3LbSV+6hdTj7wVzpBmCPfVhGLTHFuu5
s0n6kNeatptCfVNfaCL0yWe41aI7C721DrKCokqNuPqONxhTCoX2KfihsZA7GltBd/KxeimyyBJj
v0aIxGIfJ0c7Psc/5CZ0qrWzbqI6VaAUaJJVgePOUxbZ9Y9H8fBP2Pep6RLUa8YSeJycrVeYAhUU
q98e9FRMg11Gh9B4Z+0bHJjGJRjbWVGRI02Ewvu//6tpcIBVUj0eF9lCXsmoQURykF0Q2eLr+ml6
8cgImS8BXH0OcwaTFo8GA9oO2Y5JMye8C1+7JxyomOzvQDPCwF31ptApFvnf1o41IL+TXK7Wx4yn
MBDigadQcT90vNGmhLck7mvvUJdEJvdV0e5v96tZOVdu3lQMOhoasj/U4KOdgdDqSGW+3J0NaFZ8
pC5NMqL/dVvTW+eXzFXLbLh/G6ppp+sOIDJ3RSONZxFDQAYnaxxISivT7iTJu4Uyi7BF51FKQZvH
HQ8lRG4upNiVTc4S5+oCZ6j5FbA1SGZvyS1X/fLyoCvukYA/SYX8vrTrx0Ih9n0dkeUY3j6qSfm4
DCuoElLUPhKfhhoryrCmJon9ShdnEBf6pNTwn7Q9U3ZSKwlZ5wsVrDRzDQabMqYwbwdFDfzW3Kt/
FGxB4/vuI5WJ7rPPW1cAzq945wJS65YWo4BQtTpCtHF0RyXGSHN4XODVi1Uby92zXjcjF9EH4s15
MpITpDQIoh3Jmvm5Nd/w+zq4TLh+iqvXcpEil+feYG5mxeNcMSFQcupw1o21O8E5cVUnp7BGyUHq
PmVKemXbcTicJgxPccgi089wIGpHMK8mTZEBkP1iHsUk8WHqk84E1SXavwUuudb8m4hzlymGV7KP
V92cNtiMXjHSsftZBNumsmGiJ0qMH18T1vf3J/gohjVL9J8p0Ut91oa0Vbyy4wX45c+Z7J9lI/1N
d9IInk7zKsNLcwUhuPccbQ+bVdSwETX//zixRJIyrF9U/Y2NI98qi9eZtfVVIur5JfJiIufHTV0L
jEGpD1zptLPNoFj69FhrUJHV5S96reqJ8oulnkVA9605KwgK506S61YWSiz90uMZxQvsUZxlUfoE
pZBY0GHq+jRyxyHi0aazIaMg5pt9ATmt9mbmW9pvjdc5Nh9PIazFqoLyIBnisp+Bl/xP4hSotmRX
E0Hd+1W653zhO0LWWbb2pPA7I/RLZI93wwLbn/yylpr27XHs7ulaPl0JqE4zFBhjufw/J7LV1wSu
+/DSjmnUaVNbB04CSiYryM/MDR2fgSNRMuq7HYy9OMRkrxVmQFaVLKy7An5EyUNTTiF3Gl+i+lH2
/ZEZmYxk/KsHBNEL+T9lx8Jyp7IL1LzZp6a1IDGP1bs8/IgMYVFx30iww3BLYHVBKSkj1LQpHOZS
FX5R1tSoO5hq/BOSfxs0vFDQ0v5ipPZRw3V9GI0rom5JhJ97XPM8Ut294a+64DHfRL67RrLUxeP+
bTk7SdhM1nbBAHmQpy8ESTHxVA3ogk0Pp8m4OIKRr6OYeHz6ebNH/vZQifGdhthzR7x6QDcuRI/L
ovyKOnurcMvjS7yqYKacSkE/6Dw2r6i12eMtpxSCD0NCwlgEgwHfGT1d+xabPUM2AlUfO2VYqVFR
TCPXDcO07o4t6L8gj9aZYXXPHHxCtDQsc399zAsaxlA41DnWwyB2qVkW+5nc+OxfSFHYyZmte6we
BdcsqVfWZyGYbZKnHV8VTq3NPtsZK+PGUMpfBPSxe4q+6/9blwrpJdsRoOng3+TS7Ea2iiPeWYTg
2FsepzQynqCB71KAdG5FV26g7YAvUMOzuRPndwISeFkzelU4RTf9q8UWzvKt8L3jEhT3XAoj40Fg
fyPQWzt/72UNEgEdfZFTCqKHUnpbLdRAlTsUkN3klcvwHUxPhRlD7SyJZf7IYqhd5LUOid39Zxr4
11NVUKy9pZ+ni4/Y8xi0IbRxwfCXzxkQ3ImdUqW+KUzBUyKhwW6IchMH0O++NY5TP8K7mDPecbGN
/R1+wJGMBQ5R8Qs3nUEkOUq5TEeyozJXfNW//cakRz0KpSx9+ga83Kzp7sZieIykwX37NOv2nV0P
B8mQldAXpWTaQf3BhWzgoTYfOysRPKij30qb5nIaZ4rbiBv3+w/ZgORpcLcgbPMUjgrbQt5SQvcd
mb8nHlgRgK1sFnY+Q9ngAK1U+4dxM3/KJegEZ1MOZBeAaKqZTqGaTflVQuAh94ag/PRWvN/03zUs
vaLuRhBSUuZuuggKx7CHYa4rxsf6XFjejLwY50M/gRBbRorDDk77AWvk1/jwtIbrhZ8Bpfaibb4v
W1hTlNfg3RCygP/GMVD0wRdUQeHIKjjCss9rg2LoyRBrO6A6y3wAYurqnsmCA+fi3tBiov+oyOqg
EgfuaLt+HmVPTQwfYjz6XeVrlgw+ZG8LDnZ11JZcMTPag9N/GDPzvAjT9w10mbEQAHdR1kYdeKmZ
DFDeQPwgLHnf9aNgnVRFKP7kiooUD5ShDDMLe3apoS6ibTrHai8wdu5nNxJ1ypDESPf+BKg6YH0A
1+tQXSVatqNrINt979kJY37yZfa5Cl94e6kyyZm1/hR8rAMCa9ARGn+aFyVHzykZKBIqmJprP7W1
NCSbmnRc/sG2umckk1FeJR6UhkQV4QQi5sRcNlitwyaaFvn0G+wy1e8tegVy0h60bTQCww4IEoxV
xpyPgXM705DByy+YKC8vQiH6N1dsZQRntZiJ7XmG0/saJ7T4lx509ZQnqpIISW2F3MYEWuhRbBBR
oTh7ple5PBDf7VcO4/9MSq+HKf202sWQhF8D2/qPwjRwduRWzqPsrZfQ9gjgf1R91yNaVTv4a9z6
sUwAWT/w3lniPFtKjLZlztJQk9YfcEUV9J1aiKmz26gDUQUgWXqq5bZLVhKkWtK2nMVuKTZ1oca4
NQeXQSdYw/mwMS8GSE4KrNHd7Sr8kW1/BnBpWmawOcZKeA5lGcD1kEKEdSZMvQ8JD94d1UkqncVi
3wIGaHLGTQViV3aYj8OFCMFcgk/CMTaMOE6+3jK0IucLj6JsoqxBlGiABeuawEaZ98upeosjK/mH
YHRQY23hehmqIIR97xvjGwhGMNUMRjl6YkrP3eggpFjLFk4qEymuvyLPEVbWwqmbaiQMCgfcHk0D
B+CswAqW3nQSpC2dMvw5IabHCH8j5EI8PpVuHWrbcaPvQbpGSygDbbLpKwTqyASqZ03NSLnkA9Cg
0kx9jX+roK5aiJYNtN11qz9VQVDQ3EPvcfjH5nRKclyJ7cAZoVsbZV+Ns5hjKaAfyJKH4Ww3TMIz
Z1xw8JOIkDwxWgThAVMU2as+0lJ/8+WQ+nIfPRWVgdUbe0oUij7Qly3W4KShWTxlk1rdoC/w6Y0b
J4+8DZlQ11K2uGYjBZc+rI63DNw0zrxSV+teJZNFFpTDoCrvCMRrS0Kujz39yGZvToKkP1RP1URN
CQiZI622DQv9hAG+1pW3NePd3bIhXYgNF1FXDUy8g9DxORc5gC8cjTaokpZ73fwg7z5F/E6Fj8eI
IMuWjM8yxDebun7z8ZRbDk80q42TTrN4WgX/FvhvVr5dSIZ52js+4s6E75MlYelTl+w9vO6lICad
IE+IAVDqc8x0Z2b+IOlOBhV0kqBPesd13n0NCgqtn++oeiw3vaUyMwFydiyH0vglXN9QW4hAm1y7
2EEJav32ZN8BzjTFEFbmiLFhdQFi1HKGO3b1iLcek6Fm4kvPl1K7YHDltI46QY8h79Q6cJavQ1bk
MGgmAurNoUcEPAmhs61mjVlvpv5Uc3Z2kwhtbKR9uE6Eb/Cyy60OfF6j6ZitOPs2JWJlf4hTeWMB
1QQEQ6i8B1Nfij91XHeiWjkr89cS8BdGdkvN/vU2cv4o7aVsgCJU4VQF7PtC7vW8HS5CdtqBwguK
A76B15A2X+hmxXi6jpwfxA22/x6nS/Isy4rOLaAVCfHxV814DqdtsmJwiyiKD4WY6eZeIeNan8qr
7fb5030+HcJSjXynfrXyc0lWQaIntiDnZ5kQOjMXGGwhYwJbnUxpXd5ufbgTNxHYrUuzMrx4Gnbq
CtaR54fUu2z/vciI4U2CNH2X1IP104vhuiz1kQ68SBtGWnUzgaRggujqHvSpxhxw4BojS8QF3Jyx
KbbGLHP0Mb7bwU3Uj36eAfukE7z8tSNOSrO4uqWwswSYCeFZgGAJG43/tZ5tlJxd2Ej7gx43Gks+
NxlrfRecFPY1KDzvKPinEVYt+Ystcr0n1llccnvQ3n8NtOCRRoaNz/UjnlegKNJH/IaakHv9LyxL
qsZV9jJA+sZ4+hHmbuMOln5kjYYEaXhTWlNh2/J0ha26ag6un6Gal8fr0DC19eYbAuTyA270FucT
EMXoDeHXudWxYlylk5p0HjwyBnrRTN+0IiUw2J0CLNlmfF79Yi5jyx8u2MDza9iHzfz5iWBFsD0N
r0fSSWCLt5Qi5pqV2nIgR8glKBIluHgGu85/k3aW0L1IAzQOyJTEeWlpBzb4nFqIzBxIll8zQw5b
ina/co3x/ohnljdRx4hAImbmkXrr8bJLsbc06lmMpR+UXclicf/sVBxm5RhBtF8Y8mY/hjhy2WuN
D+j/9CSZVKbyLPAa6B46F2RpKX/Ds4dJc9PQhe9YQUP/zGVqpOLIZeUnJYBCX+7g4oNjBVEIyIUN
owyG+lDLHidsgddJNAQB5hkg5MChW33dZ2xOsImRs0ZfQDRckoLF+iXp8UeUcBdNLUvaQ+xJbHuE
OcCEDQjzA+5a1k/YQuJcvB8t77KjKnKKnEnAK7SGgFnfq7HvUili9CXoY/ugi4cghZssGOxo6gCZ
yBtAwFU3CzfENslzCJX/goylJS9NkYKRP5wOv8IZ3s/CEqipN+jVlKlrwqVsznxpoBZCgWCtEiMZ
qbNaGOsxClaQRi2e1pi5k4IOLzTcPNPGwdROPkjR7vod9vzeGi19ysTEeoHRahhOq0Hkgyn+SUqg
gXGJ7AyCzXVM+cw9/48enrZoiYv+BBC5qo4zQ0PGf98gGy3xPz25uomvko/c+J8ifCRyWkx0UJMg
zNnWqnKhVCjerSqhgs+v4KT8XGpw7zmJIbgAfMnxWSTvrIPI+sTvzjQS09+9HCxYIxvg8YyctBk9
vUbJU90ugnw4MWtakr5qjebs7EUWjN9BSH7LOPQBqwh6flaQnyNjdcl+OKYiGsBuVRcC8FRsb65b
PXY2ceaYMF8i9pSrTmUGAaZkGiowlhD+5NkqWSYmLkJUqd0mMRBVRfqydsu31Fwo+njgrnkZ8NjS
uWHaEQrOXuw1xmgWT5ZzGJUDsJ3Han6G/H0HbRitGDAqxeu1N1xaHvknI++eI9ZBWobq/q+z8IIs
ItdCFsFzgUZzXc2MMDYT7TQxgB21nNGlh7PpkNKqpWYvMNxxqCDad30/vpisSSggIeY7Ou587UpG
xuIMnMayde7xleCs1u09a7l5bHJWwtXvvx4lq+nfRvQyiMrmqNVqTmtVTCSORcW5DmwHJhox9EJw
LBTYFZx2HyVGq3CZvnpFeOPkr++oWqbd2utAnQxACcWJqbmpyVx3CWp2fiaUZ/fOkfSKycg2eVWw
n2GX9QirvpQ4JnreR92c0urrlLbw4rks00cIl/aSBYhQj6g7nZJ+iHGXwHew1xGGCijEal4v26K6
h9m4qVBVjLPCMr+xBgsYcs8CNGNzP7nBr5scTEtW92UZA79fCgRWazCW4Ai37qvnNuR9ElQwa+GM
dUAK0kIHAJ0MVmmnOfPQJLPazo1SOjlZG/2GSST0CqEzx3aD6g1Sddn0dnAaWKJHfbqFXksjVmJz
4t16Ukk8Epaz7zf+BL6dQwm/Qm6H7kKH9quK0nealwl4oQVFRlMYrbAX6Aqsk8itoanYqCMNWvoz
vuvb48uc7DuIH7QD6GlOHVMKE02i2++mCVbmwNXPQsrgHulJBSdbDi2barYcVaPmz+smhhSJYfmH
YV8N6t3l3fbh6uqITEQ2ksjSSH/QPVyh5Y6oWlF4TiTT+cfXabFdzodVHzvn2CV2Qmtiy0YHUJC9
PpfxrNT6q85ay9K1sjCEyeQVqmHzFuS+lyGFkNw4JexeHZWjsangqA40yg4D+LMdX8+NQIQb44xy
tkU5KllMsHMcGlTEqRijoGmDd0FWbKgp/DanQtEa3B18kTpcK79Xv3Z3eITS2nhG1MaGfFFITYuA
jqOXrXFd/vlOsjiAe6zXCVvcrXOB1MV2viaulywUk5niEPkdu4kg/rERsldHEhop/3RPVHi0UlhW
rBthZBPsQ05fimMDJ7U1T17hHV1YzSUHZhWDXPJuFyxKm695o20f9kpDSDouJvKjZlNSpuH+G78Z
a6VQIcuhPTxQTYF39cDdG056F/adG6hw99cOTOSW0J1tUhS1uDyhuFPP32Y7/Hc2VK+VFtjGMJGd
HfCjA7APBH/6j0MkNJZrAbScw0kqWEp2vwd3SDu6z34BFr2F2KjnYDQoFomQomgkxhRmNb8KsLZs
FjHzfwrF1fAP27NL7hDEBFzguV2cNn6goBPTgIbiSHKNCrcnI2YVFMDt2/JqUubcYvFUAQ+I9URf
wYhlI76ruxhqVrV2ylmw1MbelnZ4H9Q8bLh5Vg9DtOFOug2b/vBe0R06KP3St+sYRRrY+WyFQ6b3
xKjwTkstKs+oB2PuqeyGZqBkv5uxUnbp6HYGTXN98nBVBn82bNf7gMI+FCzNXlkbEyCMDB2i4YGw
pLYZ8BHYidv6zo5mHEvzfdn6KbGNHJEPrMvIFVTGwGKovIPpVoPThr6qTQb796qwYe264kqzSmZH
C26aCD50BYooKICWzxPp/PJ18e/BMaiN7i5dbC550w7q9DFr7yA1S0WwaVbeHmVfOCk357f5LjVJ
kicg7vBrz+Aw30rlpgCKayABKHl6X6DFbG7A4qvRvq1hh5mngiBkI9F4VWZDUjfHq3JkKAt9+LNw
XStSLePJjAIpsuHuM+vbnq6byVv89q6RBkAsjp+Gk7+SC99Kee9wQWgn9DG6rC8Ev9NSOixvHxPt
e8POyjILWwz5BIZZCNIEIBPnPVenIYOiiRqOtaEsWsdd5l3iHpa+n7muA+0HC+b7YRIjsJRUc/UE
FvsbxTpSIyeUWc6+4mmB0HjceHs0c5d2zPUYp60kSfqnC5Mfeo/IHhA5uSBzj7t9FeG+pvaeYdq4
9pxhHHUyAXM7HvKgHtaK6ciAQxYVGV0AuWaPARstpQyr3MsUgzcLMy27leDiz/cZ6Jv7fkeIC/hB
sntzaXlsKBhoArekSrpcItvra82Z0PFytHqC3K+hAl1BUW+dQoVB2pOmXvX4N4v25ioG3YGieDhZ
EbEbZ2fBf/XXc8vjD6MukrcZFbc+Nl1sK+Tti8EkAgQ9lrQQat/iJpjbZ37W2UGYGQNmBVJQ7/rE
2/t8kyLnbOoRL4PM19MqtrS3eWkhv5Z62zTH3NdhUKMc3/rMyHpyNFlyxJqk00cQ5DB2wbdVOgwu
WS0mGbalOwaFyGlGJ3zkXqfRZ9gAEpfxGtA2MsdwOSJbcXmhalFGHOHykDKXBDbGUCfpYRrtsJ1j
cs2/HCPw+6EBVNzteYJL+fPLyENYbQk0Uq6zt0nmYueJpV+hVXRVPuFDsMBNlN+3AIZYhnFTN+DT
IPtbvH0zp6SZJiNL1hwqO2vBvfWCOcmZDKS8gY/dV4GYEcQQ5T9pGvOTnQ8CcVCXqF19FFr+flyC
+yQSl2ArdMog+dHSl2cAPYTy+9FGxGRH8ZwMD2a1jfeHX/kJb3RXJu7wZaINOI1+I1ePUXGT2zVO
n6XxZTbudkdhYGIJD1t+un8+KfBNTGvzqsxfka/5tH/SO4W+4CQgH9/Hd9X/ZmVu8FHjIJ6wOmLa
erpTTQLBs0qENrH7AEJ9p8iDF3e9XgZQey3gnCdBTIMCeRGxGFAlkwrKg4KsDXe0Lsg0IF502xCQ
iS88hK0AlKlpyWSgrer3TCWlA9dD8I6adRDddbEXYKuEc7fucDt7JYuLR9ptMuAUEj79IZHVqvyF
GsEqJ0B26lsu/AJcNN8B1VpgolSeUFPTqgQSv7JPD9mJgagxW1cN9fE7F0GwwbnQd9dOKePpQj1a
CASgVnf11KGoeqH3rCy64Con95yi0++kX9pmgsurr1imGK6oblmlYUFSx6q22G0l++fbyeAU2LGm
gWQa1yMXS45HHWwwtLqx1H5xXE3oBMholsQqN8POqDWuVBhLi21b7Dr7xJu88U5lG5YEUF588gDI
5ljKZdkot15XPA+4+sS7w9/JrizibcvnSMH7qjFUE7qlqhlffpA0cL4RkjMQXksIhXTpx8hmIaVc
aCsae5xFzjAXf/7Q/zmoOeESsKzMqZNLwXlcxCcw28fC7GoUbqkKiCwEe9sNdeIK6IZ6TMeZUl4S
nHyiCSKmExx5q9PnBlRA8ApfUstyJfMpXov0uNOVB7TdmlvRo4sjGsr9tgN9xkL6LYoKcgQTc97L
acomNVp792kOcJk5gH/AzMulTQGXUeuC2G8RJIfycIYjiZTTNy/p4TyRBx0nLiymv//manZMo2j2
xE91IAFNd0pEPWHrKCRbAb4YBSnYtUlxbznOUhFOJnMxq8CHPozKlfG4KC7DX+IBYa1fAKjNF6rP
zlSOq7qXPFyyJVMeON0H5zrlHQ2wlbTD7YNzoa4poTVkfM7Xs+XzRJwcclMtmJOenN/GV0YMJgLN
q8Q8M8lZ5dQTLrmh1B77t7cpWjG4dkbR88S2zgPKrehqa+zpGomanX5gDEpL20flm2WSo9PWBqs6
aBt/8FX5Yr1DOMw2xz9yJTtTLKSDb9ZMdGJYSGAj1gtYuOBUwY3DEju5j3cd+a+7yzzLtPFlFIeT
4VGGkSL94W8fZBPF5SWr+znC3PJDTFF40UP8io8IbN+KLLpC6itP06O1B8YOma871a72oDCTmmyH
ekb5mbSj6BUQDzcuSHg416rXqa/pmX+R0HS4PA9/a82/qhaGQNejeGX9lg65NDxSyqdzrxDCCfZv
1TQBBmNDb+gX4zklI05yYnwf4jcw9XGRp8qCqim8hiEkr2PM0RQrWL5b9sAf1OwqGO9X0BRGSilK
hGGLvOTIV7ZKv3y4UsJG963orLifYCjaTmSkUBhAc7T6a+f3RWJBOBk4Oxsj/KfJldOamqQkqDo6
cQPqOdPPa+7+Ob+2A96vJf6jNxSnM65F+9ZEQ1KsbbvCh4yufuxb+5ETIgxTyghASukiVqD9IWkF
uMimPAo/8bWvtNC1SvMywHifj3MKeuzcFvi+FfuClC7/mLmDUw3JZoQw6oN62ukH0pqZRTxtjpGm
qTyo0AcyLjyhoI5t9jC0/NTifI+03QvYLYm34SzqFD3GDcLHJ+7yCURWcePzLsZgTM1uUuqL2r2h
qTXje5/emuH8eMPVoxplq7KxIXPemmHI122n3B/ywEYLtxSmkDMCKj/+ZkfEQvFnL7gGLOM9/yKp
fFY1Vr15bUU3wXDd05YvdQMv1VKeBCw0f5VqNbVlvekDzB7SNyqTYvpBDc0RdpyN/CyXfotUrLFG
7EuPxhN2OAze4U6vAybClq/go+IjvOXIGe+enjPM2REWHpQ7gwsIEuh9LkRH7zJ7wKZEuDj6uoNh
EElM7FbJYksN99xpeXcOVZ2SIFdI6WKtJsG/wTBro9z8dDw14ay5IQODgFieuSSmz6TUznLlo1Mv
YWT+4+mrwauUcwZhUpGuI9JeiK1cGUKTCk4p1K0iL3Jf/OikckE0WjQqEXqVdo8z+a4NvK92VrM7
iYxyXd8HzvDzUuYJJrdTLdVdts7PiFWjRl/LHjlkuR0EW0aExpv2DFv1Bv73YV6Z9Rg1GUzyo5I7
wfOSKF/mXA5fDSGw7/sUjeCa4f9i+FsVgwRhVsCUiue3YYGircBTkfoQ6sHGT7K+CQq/ewx6tTTa
D2zfLjvQCEwfYPBzrBCtY26nVCZ5Q1Y8qR59VLrlfWOnqszRWyULlNZ6/MWOZvdDLvI6VCPYRtbV
AgMssTQkv8gaYg76Qryua2FOca8kBALxvZ97FMrktgLv4Eo2rT3VVjqqg3iOXSUfTJitsRDOoxoQ
ShqgTlVn48LljE2NDZ8Go/T/CwNwfS+vCQRpOzeVKimG79KyLap/1kHxFyjqeu7y1qyk1RTbhPuU
Su0m75OkZ4Z8RbCxjD2QVDP547wUCqVwNA2BkvbzB2Y6CDZtgGnsE1SirSTnqjOMEjJkdFrU2PAB
T6O01J6IZCC06yiH17anWbZPv5LKzql9DUoeLqQaejCJiCHy+CRLwnPq7wO/ehxnHlUfCr0+V/88
G/XXj028Of0MVIGw6lq7MXGfMrR9tpK0EPJ+MVyR7fPy+WMH0HxI+YTqYZuIqZpXoMsHM10cCKjn
6BLxXhJHLuQf01+TevbY8p3hE4RtkRWUp0H1Rpx4v5QnwDIqpNd5n+g478hMAi638SX9PF6bIWox
kF3V5IraGjWk9Tu1cudCsP98mUkr5YEzqi1hoK5cNBcAC0GW5vPVs3RBOj8whquvldN741WkiVDc
SBtDv/fyJVR31byPW03tffB+QL6Qr6aUyHpTvDJgttD7kFAYn2V5M+s/dB+Aykbj+LZioq+5eogA
lB4uk7vbzhYARTR38foxEl8iOfB8+1FSdR2jh698ovURd8lmqZx2UI2m0/yWAcz6viPp9rBzRGyz
XwB58BQqopiPHH6nQaBgsbQXxwOpdffbMvtyekej7K6UXRnSGnXNg1EBgAxt9CJbW4Szv02Ekm7Z
V2FQwxKhOIBv63J8aMzUPnQBQVAm02/WYk8i02z70sLEU/NxFmVZLUTDJEW0Li9ZBG9f+VTzbYRb
zT2oCiynMAs6xWvpa1DtspGsz0lzztXQZmDksrAbcEov/X2fHUzwKTSPLq5X2AUF30tGzlR6bXKQ
IvH93Ey3P274JSGIF8UAr0jKsEjWpxtaP6vSVHS7OK8n7Y42vzuMC9n3d9BBqB9fhw1X8dkZhz7A
xgOL28WhAhZ2mlH68+sWJNhi62RjP4MAvsXIypeLIGeGjpwNMHpkW7lm8vCFYVbvYAdW8PqiUmcU
qmdwZdvIV9X3bjr2RufPS6h9cwdrgrK6soTAP9m9Hh3Cs2ePX4YBOqIgJnJe644DhUSqFbgzW5lk
biaYQ1caRGSdGKKzBddenzOZbIlMlXmZN5HbssPKyrooTLCPg80WHlAa5gjcIeJnPjt3gZaWzZ4C
l+W+nbZcBWwUD06ENrhhYKGR47se0BCwvKI0bBU2AOevw4FaOQsYjIsClDEOeg9tkPCeJe6CbCQN
oiRb+9lyPh2jD89JMMdxnJVIQfuTHjHCQUehXcnK0XoMnflkvw7L87jK3RIQXPHY4Ot1aHXz44sZ
gA6NWrn+dRKirQhp6Fq6fjNF3kqw1C0SKssmwLWQobustsmDVXMMLROQtIzJXdZ2Yb4uwZZfsJin
vY5ZARiAN032wGd7I75tqtHRVLYbURZ58zDaFXDaFgXoNAfNlxbhdvunqRJmYSgec2jiUgXJIerK
LQXiC3c7Mtmp2FkiVbNtEnbPVESjaQF8gvAif4FyJQrKu9b2J0wZgPTc9EmkpTW9vVDceyTOk3AX
Ntx+Pmekp1t0dSAclvevv80QMmoM+l4vVLDAPdcAtanmQzCDcoa2LN56WBPy/nqRLYJFwAbZBcgz
pfOMjOm2XALQ7lTZi7bcNHgAipOWw/mXKD9C6C+q31S5mOHFMs/mtqSO+gItoGqKJV8m4C2DZOoj
GAoOOWAVdtPFvI5FYTK2Qs2kf3rakkQSYr5cMf3pr3A3g3ILcj5/t+LRRxL2ACXFPT/AZIXVt5iR
u4h+NzqD68hbXYVZDpQREhVZ7QjXEfSnxbtPEHrXq/ePGm5jhvNar6jXwYTSuZQdl8bk7nue77TW
p/yN0pNEnHjUqQ+zgeFj5b5rfEFJDR5wpbDh3Ovl9DP1rqjxR/esYdjf1Wqxdz4xhBS6bFRyOun7
umNKuh5rANfWNi6/aYO4wdm/mjuoA4ur1vojDH5zW8Yf+YdOLwCN2xhatR0ydqGVr2lS8JXU9wv7
4K1tXNkmzasQbC3tzvVcqPxkjtatBKHZuibqkDf82txRE8uzqGyLeA7QTxP4dH85Eb2aE/mCuw5U
SPm8TDdJLRnbfWnjltfFHWLFpyZsXM5IsiCv6mUqTB1VrzKehrkpShTGNyNfkQnSGsCijCKfxG53
vAOliCt+9W6E1KKdL8cp+CiFVnQ61yU8nmAi1HrmOIlNcEtKm2IjZYwBc8eAWjITlb9AyS5uzfrs
jWhmsi42OZ1kuJcUqDXsUkmI4SiUuKLfa8BeqSd2ZfrKHC0mNK0Y3edvWdh4YSmboudDxvQQOlRX
8O3tvaAIhr4JFTlO+kqEbban3GojHqtfR2tywwlQWeGChrCT3LwdDwz9jpl/EVi9YHK5eQW68H5k
mFbOYuGb8FbEuvZivWHUC0nZsFCeiClaANz9QxrWbcY7CXkF/AxmtWhqm7f0wgPc6/zS5cTqo/8r
SRw8H25xdlcAqMHH8q+tr66EnPKPov02Kvaqt4orB9rP/w6DccZ1gVFHCbZ1i1yOOMjVRS/yKpSQ
CnsngjI3SnnQzR/XWHPZFmuKB8K2S6cz2fLj3kkqLoTc2is4to2jz26sDNOBO1M0SZqcN130A52I
DyqLmauJ5y5+X438/xslQuThgIOlG4h1UKzADKM6N+zEO9HcCn/qI3WklWWUWs1phBNlg5U7FtTo
evR41omc3AIGFYGmAyJUyzbpj8Qp8XzM11AsVEwHP9IINiz3ZZuUu3SlnxWju27Yk1Tr9iePlUgG
LKjKfdWYoLL7R2vvS6gBBOBs1qyVCAEJNWCRDG9Kw9S63KDzbylzZ3Ok1iyTdA7TMamfYL9mMqJp
+qmszkVrMQtuPwq/9yr4B0tI8cfMqM1WoCxDBN+VTYqkHTiVWETE24X1CXvkhqPjYnbiviRHOlIw
wB8kL9Q2+MSolf1Zsf5jla83NfyoDGLw+L0YDroXCxgvbjYH2f0go6y3aPUaibWYfMCiivzTx3he
2hk/7j4JIONP+3XgShkn0up5oZp3nqx/degAVENFoLvGbys5kIP0BWG5dKy+6FCQnvcSJIvSYTNS
D5sFIFPRw4FAE/qnX/mJI/FiiBQdJv4t8PKJxDfA0T/kPL3KA0HmKoi2ej8OM/f9l9l70nDEwkKa
GTijFk5uQggpNV1pJAKFQBv3Wd5KKYgT01+VVLidnA6qPzWK3AWwXctjQcvrVixoNmybt61M/Ui+
r23T0xRbJ5Qn+Mqudvgo2PKb4DIK/iL9+qhHU1REBzKlpSU2hOaDbjiPneFQHhIlyxY5CToKPCh2
VK7f0ae2UrJ3f2UypaMONW51fUlOEm+B1rJle8DoGrWsAaykwzTY3qcMmgqAdCHBz1Q/7itFK+0t
2+CN5gVlUxlsMLJSHc00quN4R42bD1QU7d90yKepTKy+ocmjvYDl/sJaz/6Lvb4TObcnL8cZHynY
XXnGUoFOOWxArOclGr5f6pHhKzqFOvGH2jIAFcatEFCJgVXm7r60KRpiY1uPGkGFrKKzDYeuBzxp
Vkh49xToFe1G2hXXe3wiqKweHTEkP2qecnT6EcxhwQnsblJXwZIBfwfHIUzXzJFaiZL+Dswo6q+z
ltWUeoLTUyaqJAYfJeSBUlfDki2fY9hROUs9YT9CKEFBlGaFrnldJz5sft61vZ+LPO3OR+uWwoSg
F7D46TmJdtPUSXwv8WkTWuRA5A3BHoJRHVIm/QZztcbaTtgvMw+DUCaVzfBw4/J72rQ0mLI8NMkZ
GTIbWSkodo2CASbS8Bh3lBRRwvMLuTKy2wNCHLSHhgaDz4fvS/dYh6BleqhEEoEGXOD1gfw7/tWw
tW9yo6rS4onnWEIRhcW2J86/ArGLWx3uOdiWk77O1kUQZqjyautsPoFYKzhAavCEfEoUW6OvUC87
HEstC4a6Q7+ehrQFnsBaYtUYfeAd+PMDziaLnyccLXPfJppBnghYSGlFrshiqNjyiane/6tkPXRz
ROBn4e3yT+qEgpANLYrD2EFvmV5WK5X0zYsTwceSGgp29u/sT+4QOOn9abstpTMoSB4xZURfAZ1Z
lKdO6UKg2ox9AHjnqa10ri/DYVvAHCSrXO7c/AgD+WzLHGNkcjTFFdjaY9nZUERScfy+dmJjSHBZ
Dp84zD44+ZoS0X1W/11Jf1J1UkHJDwTx9dojuX6j+PyzqBAZTB0IjUfdM+WFuUJ6kPZ7QMjWsNE5
S01Wa/s8BKOXCufEZnp9rw5xJeyxuAgrEaNa50qyXcjPxuUemZuydtNFQIvAnzeakx+i8NSLJpF8
lHlTref/bt2661R44tN5XLwIMagNXxhpWSLhsDOwFVgPCIobWWLMUI29IIPQ0NzNftb9ZHieY4X+
Qxm0yXlk2WfEWExHC1TK2XNdUjLw8ndaRwvZdtb0JJmMYGPLAdW8DpkfarxJTWU7OtV6Mp8lDzlS
AK2+q1qBnv5UpZp/JHcg9z2clgi+SQUMTz9rUlWIYZGaqhT2Urzq8p/WehwyfRB6VBfF5ZtUMCBM
AoW6PksqyCo6ZwQ4FNUdPs4RuZB/WMljIa4quHN3v59ImqF7+neJXvNcAm6ZuYbhiS9y0G2Dt2GA
J9I005eaXIFXsd5xYchCUg2aQMvn0OIskGsnSs/Pz0q/Rwx1ErAZlrpu6WPcLc3qAe2TI2RYtydC
7Bnm6ade2N59IG0lr1D2T0ugyuCeJg4ePMwulA/gRTxLYzHvzJcnqiZUVKXXeddKMGHBagqYr6ZS
xFPacBf+b89tJu5fGNIG/gFZVeqr0a4peXtklu/CkJcGjgYhMnMaluxz2c+X/ffVFVlPGTpEE8a9
K4C9tshalDZqNFdxyB/wgdzCPiLIvhk4TcnsRSs+NPxn/rz+cvBFloSnsnDn6dYlG7Sk4qGmE0U/
85U189M4v2HkO1UKp7OKLQpnjI6hLlj08lQlwJ9cuLJX7Vn4V/qgwZMaw1v+lo/k1S/aRIxEoR6w
G1GcKlPCEmjITIT+iamucAMcylgl9iQWSKO/kQnzhfSHvBKYjtNIhu7fkKgcRy9Qrr6sCV4EjZsM
lpt2yVcxOvA78wNei7vSunVZBpZ64u3XB5X43kSTfFoJ0kXJobKfZiDpQzuKvkP0cQkobHzK26jO
GGQPSk3JoUW1WfwYP9eYJFuFne1OTtT3mB6b4g+Bh4ShP7B5YlZ1d6rkd6ZmVWs6LjK69YMHs3+E
Ug5B4V7tfzv8mDZb/4yKaue7ctUd9DRkEOITcdPVpGsACK+xcNG5Bf0het5r/ks/x/LZwds/bNBP
DcS0T4zvCTrXIdWbYbpfqZglo6hpfVxu1hkZbWimjWxjJ4mHCWlLDh0AT4iAt5i//nWPyyhJ9vzt
lL73kwCpB6VVD2DO3R76UswuR2lGeL26YIwzKZLK5t7dyKdLoF2QYjZQytWny5RRmjQQVZ4prfN8
xe/O3td9x3Qq0k2wYP6NYRmcUEfl+9I4B6I9cddpBJqdpagd+VwifISoBcKLTBpc9QSzHeGiEI6U
ySwLUD8URPD8YN12USxapzkrw/1ayZA+FXQu2D8VFdv2tM9ULQkq4r7eCJXAF6U34rn3C0vGkAsk
39dXOoaRttoRbfyImG+WvM48Rz0K2OXDXCXUTn3YL/PJdpdOvL9HHzmaTW3JBlq6fzQ/nsHGNxIV
qg5VfXKO3L2AgY+kpLRd75CyELn6Op6tnpxoMg3nZaVMXKZY/sxptqw1I6HCJkD7ARxPVLxjZW1q
NRz8o53omWaaLoSFiLoq6BJmJ8944yDRbr16lt/IvCpYtre3/cP60pgkN2MRb0lpuoQ2QJdYauGL
BUicMnurG8D/7E5TV3WMtVOhMMaf/uN65UYtyNzjdaEOwJcErkz37uOIh4LKj4DnDpGEcUGd18+U
j4lucgD9UvciX2cEB02RgVgM/Jo5yXtbJDDlC57TFhSStPgy+ZU+TWuzQKikh7MX9+9u8qsZS42Z
4P9P6gj1iRH3MUUgyZPhE96noG/7hg8iuAHfu/d4zuCzKPhiQPeerHctTdvcU1BJx2Mp/UdwsZUg
xI0jYgjrHtcQZwuOiLdT8Pgug0U59+HXj6ebWCFhqOz3NmUiGshFr5ytKvaJ4PzQR16amenX2r5N
4ZVr8lSObIkcOThleuGjCkHX3xlgCQxoRZf2EOZcM7b00b4NP9OBiiCz6SkocOv2EYuTzBxyTIGp
0Iz7GqpLk3aZQcxNxJgta2gBOZDiD2tMR8TLEAQg+RB2SRNmGnqo4CftwyEyWlrn3otuxHAU5yRy
vB8VfAMiyn3V/GriHQKq7xBGl4uCRSgB+Yn3MwkxragT//5W359xmwr01Iwsh0/U2ySjGZ6BcU7g
d1dzrqaZdYERgtwEsjislzZ/ToOLgAahZHcbu1QduM6oGGuEzC5+/jklv1PWuSKl8Oh3ZpMci9O5
AeoIcXmMnHzKZVQmAngRgG2XyhrWOTCD9QG+EOD9AsW6znmtrv5U7WyZ6zpFXqAZuCJ39kNdQCEU
WFy07oiBfFoH4psF76i3kOct+a8pgFoq6mWFPmbv13ahidU6de0xqBs6oNb04Y0ESZ0XSy+IJaic
+fS9RFfWEABXxk/jomsEZmv6pyok+3kvmTv43NvbBgX8nio0jAHLCIq2Opd1B0KxXZv34g2N+qTn
zx1GDaqNbzYxB1kOznSVg8gwY3Yg34jQOkbr6plYlqRJVG9nNYSoiGl7drFYc8dv+ceFyl3Dxf1n
BuoRm9Q3iyyiuQe+to6cYENbU2aVfqZY1lUXQyKGR06fWJDJuNB7NqQdppi2ZjZjpDMb6qjGBckQ
2/TBD4XhY4QKwHpkIaBAlZwtUtvF+5KstAcuKMAkQ/MHnfGx3aoTmw/6FVJqElSSwbIoVSGng1rT
5jt4rjp+n6yxygSL9HePb/hD6pXiptrdWnsWHF1ucuSTwXcWKI6JoOLlJh7sVp1PXhKJtWVmUnbY
NoMH4IxUN96KU+56EtOK2v1v3MWNf0nEo4fKTHSKqWIiRAQd/k0tPF/N8giiLgNgrtf9JjGvtmVz
Vz7/eCRywxy0LlAMJqQYpKXTCO9TBuZtzCS9fZbULnIlgxPOKAH2PGwbBA/ALZjcuzOgI2jHWKLf
KUYrWiUbrAC91FnLze5KtgnvrB9pTNXI3sv/ST06jeLlbfXTwuCGIYNqAvmNd/7Xc+b5yzQw+us2
C58xyD4+bKrs4oigcA/WLTZgPnIpkVfr/VgN2MDleG/DHVCeXpGRJnpKjvMMPd8LtbAUrHVMx1j9
xP6KtV9eA05pKs4WnN9TnoAhn3LxDc30AVgMlkmKn/nB1WPzDl/y2lIbHKa/GnrSYaMWWlKH+uXd
KKQyQNQR0ApCyLPDAOwjSM6heLxU48eh+NAOA55MpkzZNCyE1W0+ezsPOqRMZs2dFPtd/buQyERM
VvxACixNGffq4rZj3iITiQqyTvTiMmFzho1nx+qDFZSyTxFxWhYCsbmUq0pGUKj7Xyy8+YRdqiYI
ipkLydMxPxr7S56i+suk7WZTVpZ24YxZxk+ReU3/n2w/Dip9uwUS1+Xrl4QpQbEU5rvEeMqA+hEC
KuyYlAbxNUBJzDyjDiuDG1i54ZC3Hbwl8c4/yCVffeV7qd44/sHdNOJQffJbDr4eB/BNy1EAdM9C
/UuX2nKg8lhL3y8AaMERpzdUZy2sLpupmxirNYC+lHLNfxrg6a2AAlsbC4RlFilWGqoznx5GqDSf
AlVtGt3i4Z2OcWC8JKrczzqCAAK4YQZBZ98/OMAjDRPAKBbuao1/gy/hOYu4m33wWrxWMfdfrsof
ZuA/nozXYhebOMzQhcbcBpyLQntFui5lM6vw8z4X+X9rxoMngeko6R1bxtPCGgzp9C0I4YJr98Gg
ZxL9GUH0oEvbdmMHgYVNyfwCtSqT0EHhR2N2RRaayJLz5oCgea1Pvd8jteVxMZp2WRIDZY6SMlcE
LVaZq0e9ncCvPNhLxQDIAThYVtdVvTskJ6RjYpoWMGSTQJ9yzw08ax3GTdfCW6yWK1ckFbSNNAVY
8B/NZVF+FSNwq7oJ3szP5lO8o4BwzUtcOJsmvBJMeRqNHZOhFr1LIgIhbITcLTFIWL+UNDXuv3WT
wfcfalrIuWWcbaUZMQdkp4FE8w0inuHnFk2M6kigQxJLy1KrYceJVhFl0qaSklkWValhLCq7J3Si
GdVL4oNbwOvhZ4XNu//4ZQoEZKqybWSrIoRLiUNuxfWuyZgntdz01pZziyWZ9pdYUx7lz7yh9Zfw
0PizaQrNlFL8edFSozMpbVPJya5TnquyAMNaowQMzkRAeg2xjCHu5eNbQ9aYyR550/OCSC8SnOJO
L35fjk6tAdbdm5ZejtRFWVSddR/cr8VHyIh9eWWvPhW9xVnoBEEufPAXBkuwuvevzzs5E35xnsir
0hlQcQXKRfAsMztJZEj7NHOphpDlm3RZTwhPAy/GqeP6jsvFZrUtNz9Oe+simqFME1HWyA4pNEv9
47aAiUMtyC2BfX8X0X1fdwBo3WQW/uQ4KFYoLeqDWKo+NKG23p2qpZPdxDnLBSUjgS4E+i5mpIZb
hH5I8YBAHTwqhgYX/dVNhHCMuWzg4tDs/pc3TpmIEScHzZynspwxykw9HM3Xz48GZDc4LQzgmqnQ
73pXR3AzX0HLI9dNUOdHqFYFIobavSC2hUfQVJOQo7ahvEaR1Nra/9yZoOFL+2eLl4j2JizDg02V
MdVr8XTqZEbuFVz9IZuQCWTuXPfjstvBrfuk/VOfWpCOhZ5lxWmUX3qc1aMKLSpgL+80YpxWXUB5
UDSdyQkLN1z2ZhHM6mU0qGoq/QaTWsZ+CP7EhZSz4GLUdTWWZVvLl74M2b8AbobwDt/wWv6q6oQ5
Ream+U+b3mRPXzIBzs2Vh7JM+LTRGthw22PdvTlv/+bHZjAcHxodzE6trdF4aJFVXQidSJiD2Whz
PbZf10GS3utnYv8kKd5p3rjmq7uF6huYac5bXZYd9B2bChnjr8lxcJn/+TWVoyWvj0B4Pv2+FpPX
GYrQWSLzky/m6iGJuA1i2A7PPQLtHhpaIAEjS5XgSEX2QOX0dewYkxVHe0lbZJflV0BdvrCyH52v
IoDYlGLJVSxuOd2/sTr1u/CCBrURyDxKSQAt7cSoZYkGM1VLjXIOzZVbHzEC0mZqZ3D0x3Xwbvu5
iKj4f3823hPzDHYPPAiAzDni6pVDXDbURVAa3MB7m3KLlrjkQb5RXL3e6HCwf5Gpoxr95BTS4n0O
ItLll7r75gD5+zKN5swWUTWuujsQiFLBmk0mSmhPzJ1+CrKw3QY8d5A8bzzRDt9U1MO3zfzehcq1
gyEpBIw0TOoXc9ZOFqAU5c0SkIvjh1aieNt5MgVAExWuLDF3yLVX9awtSLO4+sudw7kiiJ8XQ7ri
d4KBZLzddbJklsZFpTYhrrqqaWnqAsdfJIZFJGF3CYAN02ALPi5mv8XVLT39AfHB99xBxanjaMtl
Li3TMKkL20CrIbnVr7FHtTuxVka61SqVtsQOXhYZ1dymYupaXMIWsJRpYaOnEsJm3y3xZ4lEAqRy
xRsvp0OxVNpYgmvsd7HHh2eBj6xAhL4rpC4Zg4wQQek91N/S7hT87r5M0D0F25Jnp0WDyZmHY50L
WbIt5qXNB9/m1Q5kbp2dCyC7/vZ3ICroHG7nsOKGD54myRlbzqsZKYc7nejetKmDgol9tRi0hvGV
bSsdSyprYUwcmsvlMfqpxB6/Rpd2D4w/lj2/PMyl6HDZIEh1wLNOaDeUX6PrvTTXWm4X2KTY8u5V
ptYVBfWI77IpYHDlfw24thzmy7+YQ+DQoSo8rzSqTgs1MhCRWa+DSXu+GnMFeNit/9xlK7RFEFK1
rxCZ+xjyU6J5IosCeGF8e2d9gIWCgyEF+ruqFvLXjJjvpTDCwIjujKlu71DHFofhBzo5+oG3CeQT
3LCBko5ya/06BmJgrmSC36PmvL8fSIphZzhR/UtUOuJlnReeuCFdz4FJOy/RPLlkU4fGU+BOwAJX
smVxHFs3Z5MyMMBp/w/MQzyeuUPp56S+0n4rY2chBFClNBfKSQVwUM4ifoeYceGlXMPXoFmcXguY
ivscXyNSmuioXTQM3pxZKUOuIxKVjMDH63D0N+6/bkUHGb4zOc35E1WB1LTdZulZMZJKvurZQRl4
tCusrlbh/0X1AZ5wdE8W1vDje69VaoFy8np1UzGpF8EfQiHAx8WU6JXLY6beSohM+xfTylkXgUJR
3WK4Dfjzxc4s3QkJgB2XNe2fjJY1Skn/pJtkBWmyZOicSLG0pPkbjVxZplAB6KpeRXMofaXPJjZl
5/iC8I8RSdglEpFCrXiZre0FpcXASIqGu4zj8o9lCC51KNJ2A7u50FE+G3eBDacfc4kW4zn4Qen+
lw89fl4BOyjbVUUW7/h3niOFEmcdF/iA7vfPOGDtNfHbyJvp1SSNcwGdJL/m/b5vbAGC40eFleyD
iGvaNcb/SGG7lWlozP9JXFyyiHZo46/fO4ua3kKhv3iPImbNQ7bQR/r7Bu9ynDw+/bwW8ptSD3Rk
1wzOOhdr7Vly8xPXuKcrjlRR0/ZkjU8slWt9NgHyxPK7+8L5SZecg3/3PYtdMLlzIPKswqFwOYGs
2sRsH2H2w8m+IY+S6gCSjLzobqsn+Niew0wpEEUHCFJqStpxJAW8d9htG0xdQxFTPnwnCzFWfx1A
dwOhAmMF3Sb8vsow+dSMGCd4SLuJeBC2gOW6RYaVXZ+gkjCoIMClw3popshUcFTo2AfzmlF9JA2d
JI8QNJKU5FLzAgaPCtnB5ur29SpHame117hUTB5gj3oEyyU610XdPR5w5iBzebSrZ14aOByHuYCQ
jTRGHXdvCZJq18a8XDLakr5G4TL8+o+JBHHy85T5du16wozGtnvGd+7lGgjh/T4tnlQ/QVxhFgTv
oWfj1FH6UX0KjlFDobcQCTRfH618kNR24loyzoLfUuMA0jfDq8XHW9nsqujZjyjDY/NjWJdDUS9A
wP1c8np7fz9lPIA8HlFmtRThFwkuLYAMjm7tSKjC0JkCeN+HNzp4K2vBYRr9EX5XL+Jda3aiRKCR
9+UnNQeSxbjJGt/QsG2pKIUMkEyrw2S0fEj+/+rkwI/e1H4LscVG5Ty+4mxFTD5YZfW7L9PhFjL3
R3aBC5e1MrkqTtODeWLlND0qDxN8AmsJG0pIZ1kCn6u2NVDBc11wSvOnny7mP+wJ0WtbeekzHrYM
UaqDG4y7G11+NQwNeCTauCT9eZtmiYu0WSsmx6DL1cb/6dsSyz0lZGPxd2bgc6/JUEnY2ew8o1+L
aZR/m1a1Gg15s4Rq25UFqc/T86vywW8Ba+IODnc0+1xytJBuf4tlLdzjjdIaDNwjbkWOV678ADJF
JVYDQc1EgcVJ8HUWEkfKUSFWvqCqdf9IpO5hd0xN8PUe7NzsWHBXaWoZ0mVrTxRMRnS3UiTe3EJy
INWSeN+g5n1Fu5/08OcUj6FMOkj5TaE/+dyyWThbTAXtEYbynoO8hCaN4FWBj3DO2yQQ+lhoORRB
ztcUJMuHGKnDDumVl+eUog/gKXFC10kMffveboFz6GQ64IXDbvDJcfnppCFBkyelnzdihU2jJ3fi
eZDB80aM5zoJK70KmePb6eMN0pBNNWgAvf0X4dqQ/7lrr9oy7wPACkZrg16EPNmnvwL5RJ1DbXd0
iYav9cReDbjKQzFn6H3g0gjljr/k4TC4aN8vteNR6jEe4I6BvWa5HNJCApaLMoCEf+rKOOrs0hh2
n9p+g+LEiSsZZ2i/UpLP8XPYDmaeyHi5uE9TI/5ECOqbInlxw7eoC/vTZDRn+xK3NgoagKanJ5Oh
bmUEeau5KsUj1IalmuxRhdEhMyjhVZcDKCRcijwGsAwQ2z54yoyKEvOPPT9822m+nO3528uxa09k
s8eRFd+KvcQMrSd9CaBWZblrk4QauAUjUpR3KFeLWD01kPsVP2CyntSS42Uk1YgltAOus8UoIs6P
vtmPPo9QXqOfk6aR8PFQfCA+/te0LJIUsu0EDnsXYx4LbJ5wTQ1iXKHVlBtB2PBfmkU7zHI+X2AV
qXi5OhbiFlE//1HS798V+3uJNkIkFx5+dLSbnQLWUfl7CI90o0V2mvp/1jXkNHp+btBdagsfrg3S
QEiOJG2zGmo0d4CKX6QudZFFr4lBlhMSrxb5elZ+/+16HcNKymIXyYYNJfS0xXDrVVSuvIbZa1pd
eFUSYkgbtKjCq9xGC3Llw6A/FpcoaxSec0pVgdAqPLZa0lYBc7o3SqoE/Yr/GUn1gxMNys+HmZGV
/0z51zkI/1PBb0ViyXNoSA+TRIqZM9xACw3RyNwB/OljO+02WYtWT6pO66WR83tUru0UowTd0m6Y
1P723MWp679AhH2Skf2eE/hkkdJNkbS5e8AjueJZ5TbBP+zoK/KiayRkhFOhvvYutqWMI5O90GRi
WPoheG/u+Yua3X9CcsxIJRaJY4EMdYo9gwYkfTMf3GdKNJY+3xKPecAtJNqbm6uzGwxzeXW0iW/r
hQkcXUM+v52nwE9DHFiK22o28BsGgnU8TMoNPPLQ+ra5+iVV2ufPhaAjPuMyv9cEslGrVyoP8lm8
wUrIBNCjyOuXK23shXJV9zJO5pbzxzZR0Qwd4AiinABYRiVZmfr9DO6vUfHoAfjokAwPB5QzgyrV
k4D+3HtBp2lkdHdzqRTKgTXDN4MNUFJyr4hBGCWFrwbCwFjgTwnetdHX4L92b0QYi881VYGnbSHE
/DCuzLUhOyirS8KcBpkfHZ5f6S6d1pqP5myF/Clqfqcy9qLa9N6EOxUrwV0YS2JdqHoiLX0K+gxG
N3M2+eXBg34QHL8HDgjym9rHHYkcTM7KdHwbeOoYvv8A1Hl+Od0ZIA3Wl0rJivROgxQ+eMGP3lNX
wS4Z/JRE8QZm9al2IJhQGELBsxorL4F5VBe57DyUp+LWgv/PiKJOcdIhYEx13w5zhhLKUhGHBI9p
ZDe+P8kyr2v9pKJ7zoqBB5RxbHa0sFqcLpr+y9xqZHFWUJqobATTmPJu/gxbuabm70lGkxQCNV9A
CSRrIu7IvOeqw8QON7XJ+2gJra0K7MXq4iedBvSH/DxGOOrs8/HkymkC8wAUN8NSrTX/NxVUfHMx
jo+gts+cOJQcPb1XATWFQ2EA1GBdIn6rKRxv3Fk1eQhr7xCGaNHq7aU9oF9rc+R/fS2FEDNPvWex
F7d+2wZex9GkDfng801r3BUbIimKo5WAjv8WoPcxRiy820VCrEzMuSdQZLdVAldyLOs4Chas9/Ih
/w3xDgXKkdEr0DbU4O1KAJ9EwvNElqSBsmxNLFDUCnKF+OrXLIwqh4K8eJKUGelCrDymsdGbYDB9
PMsfsd74owu7crYMfylKgSW//N2SjZkChON8kI6vs5bWzhm8rLFUTR8tnM32K7krAeYh+dZv2o2+
F8RX7AfBnG7zY5KXAhbUX9cPZkOhdyNRB4jv1RvJ3EtH2h7GY8qshow6Rru8u//KZkEgMO1X1oLF
2yUnsEEhgX7VfaVuQfg2ZD9Pp4knUMvEFmGWG9bg2HHjKyPKaZfrRx5kfEnyrwUWWMOFLDm+34BJ
i9QTC/reZIvv4n40RW6BlMIGWgAynezaummBf3lMT+Wy2jCUoy97LAKpvqDGZ3c2C9ivgTrPTgtl
n1AASFfEFpOiiLU8SMxbeKbGcKj1pGy9xxgUttpp9w4ESKTrbt/iOrpBdP4OdS1vU0r2bkQ0VJUx
8qAbP+2EOgk+1nBkMEsvfQ8G7dMNQkkzY5JzPKUT06DT2imIBvXYoBaqzMzbZPUqHXE/XdJ8y0Qx
QBGyedwOoy2P8t5Nogknj61EP70h5nsTu7dS6u4X+Vw21rnwu48xyUerCRruHcjznbzWZ9bRRiI2
Z85eVeRF4mzE8GVqrmtCzHIuw/tHazpJdI9MircdlCOzmcBOfFamdhd4Nd9z69+EQSPbfSR2Lju4
FC51COk61qDxHoQGvZEf5XE1MgC702eferYH2oAfJtdWS1yQE6B8nTC7LnkrTWuUzP78TZgqT5OK
ON7p4L5dWk3bf2Whi/Q9y9tGhhQPq5db+Vz0tzqw/MR/RlLMb+K/OusQDu4sg5F2DuOWuNSWAj8D
25KtjY0echVTbQwLLW93yZFVKN8AKZ+4mdNn61T+tAFWIgPo2GPC1yRcnLZ1dCr7HIBQYXLq/bhl
JhwARYQW36XgxB2RbCZl/2MdNPqt0LMn5ktTCjaPtJe3Njcpeksg/pkkUQHI7MQlv4cyYbCNuEy6
rvJjmYu9fPKUbeRbHTh5E4zq+K0Jjfi61HGw9PxNq7/vFlzn3RWrejOCccQ7nqArMFCsjpqysCSg
0GsMwxxXXb8WfHlVIm1NQaGyqj4SYiJo8LWn4YU1KkFBwRsPlMRIys/aQV5xTJk3Wjzzd7buhbX5
PjObRJAdbT6blH3BmxKcUjEoZQoqdmvXYzYBVH0zDjEUD8vf1sY5j6O4PUgQvGe7vv/WWNntPCbn
F/rE3TwqyRT56sZ9Y4mchN2GUnLeel8adw0Yd4ndU7WhY3WPR4eOj4Nh5e1J3DWXBWlZ/HEFJIQ5
s1qm1YP6Xy3gFQRpYkFXxlDgZhoaAcir1pnCkCgE4NpgNtJtN/L1q2Z17WlUNtLYL68Mb7bkeodr
83TXBgsiNUBm52w1dTg4b7HjtVuShPJnUcxZ+o6f6poBnFWsOUOI50gRTApFYRB/LGE4sfuPSiBc
uQgHOufJM8u6X082HmMiOhqDTgKb9NS2ho4BbV+jBEZF8wdQUhlRSG6h/+tOPkRbYwECh+kaHZ5T
41xkKtS9766e0n0bm7IMhno0tMqPOxT7WI7acIUiI2+BDGQPW/Qd7vYqBNGtiamd1YSYcVFwdiD7
vKDqkomJzh5gzbggXdDZTroMnCo6R5lrYErjxNTKJZHbpwVC7earlR+njc5ZQ5P54xBpuTZKEGBK
2WNClJOkyKQ2eR/Xq1SVIe7jjdEbyS9OU0ijCHpGPcHs/+lvwUljmGTTo6W8yJQdI7gLhj/Z2uzk
kA3EqCx/wwnkokB2m0MO7WZu9Y1uUg6Nb/TNlFkwTPO9tUwkXWvsZvt3tDYZyDqi9dt55V8YOzVY
mZPlx9WZUD/PQcWTryZSUQY/cN1Rrj33U783EqMINs22bUm3Aw7yjfIrQd256MJcp6BzlkwNQQej
gACTOrLCTRL4JbFg5cua8xAs/ztiKsFR3i9cVI7aL1yvGMJ3h7mJA/ER6miwYPdIcLIPKBV3/esg
st74HvrT40YPUJQrrWzc5wL/Ij3hzC550bahwvltbTb5aCDiag8nKi0gvHGcb9HRSjEerqZqKuHh
kTvipj7XeWYA/cfqqdM5F3ZAAdo0bXJnc91zEIPSHQfawn4Xf46bfCfwPvQlybJ7iyb+RT64qyfR
f48dgPo4jp/h3Ggp+dlVATU4I1nH6VVXO6d//wJ2GJglaEfu+7knmwI6iogQmebtMGg22vqWTFkA
0ryHddK1jqaaHWVLOlBdt7hc57DzSHBhJ/xpH3s2NLHFXTVFVgg8gNo0/AFEuzh5+agINSzUMjyK
fJ/CoVdouVkfYe9Kw05o0prHdHdxnw1ktGRs0yYPqQgd3sStO6bM/XaVNqoWs1/AfOyRb2Rp41Nb
HJ8t4JK2uoBkm+m+18jD1obIIS89cEBgPyIBd9pmpN75vyOEo+x072BnDFbSJArvCO45uaReCDMV
I3UKyQEkSmPYS1rSFM6fBg3pHc84+CERTdNTDIcXmEVLCSlibu0iS/zcS+4g4ByEgb4khkxu68SJ
DLpKqsjqalzNL+gKgob8Mw2ElRnjjgpxuMW8VO+ZY6d89vLHVCg25YrRPhivLTgZvszF4YTkWKaL
B34FJjyxXYY9az4TGXa06GoyPoBC3ql1TUShRivislL4q97aBdhnJApCIK5gyPNK54gyKgVuicMG
+ntcBDx8Lvg8/w8bNZ4IwgKC9UJScmrpSG132JWuMMbiDLdpoL6MSh/kIxpy+iRWWKQ7sc2+/anQ
oixvrdvTZipBBD8Hg+ekU4GZ+sSsT2V/PEGc6HJXC2RHgYgCyx9lSVrR1Jd/08TTFc/ZawHVnv/K
DVmR2I0NXHyqU2ACq+Gf7PDvq+scqIa7saD90eLNrO4+eHRbJivBBaNZMWUk+KDQAEBmuuKjQNpL
hIfVAyGxLMkGs5AZ3oVhMDGVLrTT4afr9GeAN7GU4Znq8iQZGrzvhOy/x04ryHA5bN8uGqfvamTl
6rHkZZQ0d+uecAfxM6hjRsL2bG7fk5yrG5eTFf+Mu0E2WqUS3KTlLWYxH72FaWL+mvp5iezGb3Gc
uIw83t72zA5scnqvpxdZrITQgi+HGRg3X0KOxnRer8o5nd7TsKc49FpZVyrxyYYISbBUx0zigYyG
Op+QHc/symmwfDtJDnQS4bLAFT3MJXd2d6qhTseCvfzjsnbT2uq+J528y/RW6zNrBqNdUm135dv9
f8NWCseF0T28OBkTvUMIhrB/HGcqg8HIKkF6nnv8pgB7SBQt7ZyxSjTqfn7tNHmHh5f9f6U7rfSs
eWZdLaTi7oWP5Uq3I6uPj46gUom0SyYdVfEIqv1QLBxOWqk9rFi3H1T6Ij5JkYwSNgMD9H5O6ehn
c1P1nZDvVwNtl3Yzj3jAGpfRtZ2CdXgSGkraO1h1x6WPoUkT2aB9WF7e4yPTZWsswQ3vLhaspprV
5sc1BHgoC8q194dv5Cj+j60EIAbgNUE05lZpAbuoZCx+5eIK2i7pt8Tid2kZT1utDNVVW78vbikQ
qF04uen12bX9w99XzJaEWpGTlCCbkypLgtcTPfeZ9cGZksEprVEgovOfKy/XcTy01hp8H2u/dPum
iwhK7B3EvDqDXtDjjvWs1AETFbNdBpFfDIZrVuCMLM+jrljfbRS9A4+z549M2LGfzKZ53Nn+1K7E
WUEAy+mGf/L4lDD35Fja6PldkZugMO48RYRlCx9D+AwkM+Iy/BRr0JYbG8vePjODMB6GUb6693wf
UhQ+xiIevV3pT1oQtcbUEzBH/ndMQcyILzOUJ+NNPP01zSGsBWvghnkR6yiZ0d+29l2w1rgs+C/d
nSPxxqqm1eOnnHOoW+YdPgpPVP6OlZYwARKuDulKZ/PssM+ujzBxY1199MoLBxlqmZTyaPNu/ugj
ybDKEDTZvK7JxSsC5SWuSjTpWY0xYd1S++I8XlRkqWUZ4IJDmC4fU9D2vSfNxASaqSxzWaX4YyOx
OwBPfkbNA8eapeducC2d5qebBfyD0EJsZyXvmZezfnE1goTigaf0H1AUpqy9eMiyJCO4KNYGSTb5
3Tqd6NMNDcfWSj565IEkXglkjKfQXRskUlUE+DSnF8+XvljvSwsuMy9y8a/S+hDR9Jok2qwXfPm2
7i4T9/CG6cwtR1aLpXc+ccXvFzFbfahssDsBMdZxQW0Dcx4ZS6ScgAx5u7WW7T8+RFikk9wVKX98
/Pu7K2KIbjNEdOt3062oe+HT7C7+tQszBd3T75wIJSUaQ6XGPsoY8582oiiDHb3w8whL9iqz2UfO
AGm8NtrGS6fpB9O805+2NdG1mEzqPNvBbT2uApXUYL9AJvXo1SlH97+jiXWmrxpd8uLdC+t8ScpP
apslh86BV9s/TMgkEC6EveH34uajIxov1hnOEflVe45IBvl3Dm23sD2+AKbY4hgZ7k+m9GPf3pco
hiT/SDsxEcGflOclQ+Hy4MbtQnD+17iwSYcky1OU8rOiB74dABTk4BkEZ9hBAe2gKC0VDh2ftD6/
DApZ5x1QfaopmCHVfOP0rNSqRszA51AM/RsKSbomv4NYP3x7FImsvuvvJOylC39pw1JzkvsB4B2c
FdNDLXzSq5l+nLjhxbD4LcKYNK+/MFU3X5ftNCl/PAuyVp0Bll/uWs9DrxcAKnjZ/58+20G2Ftvk
/NHFhsx2nSUcgkAMbC85j6nDBeMwzX1ntl/1dns1Rm8js2PDvIVwV1P76bMmRJ5wgKGtS7x27VDb
47e95y5Q1fqCCmm9e9WPZI/QP+9obOO08cqt5nzLjj1jugxqFlinnDYqyI79rjTzBfmTf03aDyF/
LcPR/uhHur9hgSkUmtyP9gBNkEZyu+TW7BotS6pWLjqrGepQNK/lX+cy9ETPtAy+JEgPj9TrsmIK
TyhU0P5//hCwY7Hbig0g0qwPFR54MYr/wX/fuIJOJaljeGS357MgiZlRFgcUrvAMgnVxOc/9yguB
oyMNMGQcVxBKr2wmyD+viNTTsxPHTDZAb1MO+RLEmQGCW4aCKWOQyvwIAxp3QkMuQjJgcsOLzERU
/g4BIrXdjUVJTYbCWtNttEBtm/CrgGXSQnFspL6rm8VasCZidX+m8OKal+QGmSLEQcRljQYbljQU
wQyTfVQBneJd2NAK5xuPB4LRN4s14GCx/UarDK61WX2RCE0DwDylvFz2+FsY7tQBmir9gXnskQ2c
zL1Pv8mZ6aVt7y8p7gCUfcMyM4HK9Xmgak5zTpYuY+CacUq475LSgd8DiAxi13ahRfNBaueWYqlA
FPR/Qg4lT3HkRlMBoc8I8RnJgeao01EKlwv7spgHBVwZBCrwvhrhMf+zwfp9/n6KEU4TdXTue+cx
pVV+GB8390G+yuIrvXaevutl5cfgKFsKy1bnVsiA7DtgkbjdRtZJYHSRnNWJ2PBV6B4QbDP7Afq4
MzyfXCU+OxPFXs8b8e6Js3aNjOIBHUQij4fPjymtqGeZFLlM8SXIhQPKRldM+z5f32erqmMGQO1W
AKlHLz7s4luDaVDLBPyVmqpa9DsHB82m4Q1SVmWSeujl9N+fIFAT+ug73Tl9/ZcSRwTHce1RODnO
LaXqC4rae3It9wU0OsQdrOYJ67xwaIRtkfYXJdxnJBqFBYOKCqq92wDbiEmTQGWAtdi36pJMiBUl
K+1FmoNsx/ssSgqnbt7o8l5TU9H+aEn5gKDcpJscRlgm9N7wU0hX/9pRWl0UsmhDePrLFZyZT02g
xr/QNXVEjyjYAtx3Sn4yyRV1iRAjTMeoBrbn8gk7rsuCtp2SDK+dLIjbZ3/sgu3TjeANLP1WpNKY
MQclB56SyGZDEgP3ODLgTQyqjY6EO5RvFuKnMZjDaKLAO0sgw3PkUjG5pPoARsscj01Cl260DHrF
qFY6Rx6F2DG9FPEh/vUTfT1tMjGLRZ9buW5M5WiqqEHoZGR4qDfElWmz67HKqAAAoB9YEekvbFwz
9AVGj5Kn+r2JogdwAUfGKkJi0eIHcUfA6lhLbq/YPy7eGpU/QtBdhA8qtkS1fekIMjij0eDfywKS
hIRNm8tFuNtARjCfWuN6cKNbWZAUj2EbCvelbjDPIg8sOOaw4gq0+eiOMuJ3bErsJ89EvmMqKViD
7tyD3mZOGPqexYjjUXQykh/+eEw+P3qhjUMiXkw7/P9PddzVdk5umV3jZoEIwp0rmvYxc7fowsCu
gHsTNwwNiCzlzDlzaUY/ir5PUocd7KAzZmiU5gVDvnnc3NXG2b/yLi2ZmE3qufsRywsO3QgnJ1TJ
UQjbJE+NnptQ9mqzioGQr6tGEJ/d/n27lWk5KOc8YVG6bJ/hSAh4S2z15lu6Fp/sbNaMG5j8s/WP
xlN7YETl+Fj2skYYqJ4Sr/IAAul1NLme1MuGk+zUr7vhoNuehr5JyIQ/7hAh8b4s8DjtcZ/2dPrC
A7/FH4RNAf0pSWR3uhRBjxesjXSo0J9uqiOAG9x5bQHX3mq1mOaGtlVoqoGJxrySeDap73zQL/Lk
7GjK6FQgwb16ihBvLwYIP8uqVPg0o7eRLuVOgcIPuf1TD+2e0NMvU5oSxGvnGr+nHWc/bx16FSqB
o8E9tXI9D94AIs4UJX1FUHw0tZ8vDoUhJFa1oRF+RYSpSuInEakR2dDgaLB1Dc+17n433BdTO/j6
jeBosgVQjgDusS0H8YiXn50Md7Z87XjYgalJnfmuy6SoVaCEyG14LHHfR+jHbO3hKoDbeMRaztzv
+3rAujKHq9q88bRfeQqLg8P68oltATpP9o11V/4pi3z3Qn7pOzkzQDxcMDaakSNG+1BHuesM02/A
+FLlwkoMLtFoyYdF62GcOT642NoxFrTkSXBMsmc1GyNRqYZV3Nx67FceTH6KvCp6uOR5Vng9TQxS
hUrP4NNZQdqOxMUiXPX9WEt6S9OhLgfU3n5kbJZbozjej6TqAMt0ffMQBoRPyEl0Pe5GQEM/OiAQ
433EuWUpAzicw+jlukxw5AFjdklJ8ve78NR3rHqdcj7RL++oBNNACEl1f1GN11G6iqMgm1Pfj5XE
bvC9O4xan8yBd6KxOphZZ8A95dyueUhVXT8qfv66N9v4tRCXpQEDBAslqyjyN+Pj98fsfC108yk5
DV67NseyqtER4/9U0LL/fVixiZKia/u4DKD4IMzjZr10z9h2uFyn52j4E1enIRUJ+cJBscbkhdwT
NGvj/xFI9/wh1yoJQCmXIpTsJx0Sx5fZKHlZ9SMkqwScgItA17VAR64CSmivoPegWeB1rM7ylSoM
VrD0Gqn3wq7LerpR6ahqW/qPLG/t7HZ6YBOgbgJks1oSCjyLDlunuzZsOFQQWzNCmr2bV8HOPibz
pweKsF7f4lKSl4p0Fv9hgAuV3irHt7l+X8qxGim7I44b9dB6tFfEBGzatMLiIPSdyQS4X53M2zOb
4INn3tJae7FQKU+x0vioXk0IUxIRheb5A3CknriMO7G7leYWms/RHK6zq3+YUkH0+ocz/iJ5McrO
GRhlXP8YPrQT3H3HIwKGOgdfS3WMrLE3O3e00D5xLWbTDo/I8f9XAyNdxYCc9IznHaZthZDYAHpM
/vrPitUuGrj849IJi8DaGd1wypHUsY2ivDEEtPE4ok/ka3a5j50kKXThXGGCm3vBzb5LvvOJMF7o
6JY36mlwZ3IMWE8reS2nUF5lEInKudDvcQuFJW4jFqumoO+PSocrlZZMn8AUiTl5tGqLVHDk3S3M
hGMnnmIqUAHsIE5y0X+l+x1tr516C6WkEzxUPPhcARv+Gjodq1xWIsy5xjpRiEm7TwUqzn0aGS2c
avnAGtWsfXjswaT4uZWO1fAuElYt/DHvo5GEL35wQFzD1WxX1Q+G8s2GaZjYpN80dMcV5ePW1sDT
c/SigfvtLkxOFgMaNrc14ByIAHv1tV6hO9TFaapAxCX/Efm4+M3t7vDF8WoKYPdh6Z1YfYhCamx7
9E2i/+2N6Nxptp15nSh0DxdoiH0n+ZJVZ3v+O05tyjuFoIJTiQO/ohnIGlN/qO+2/mlG5x7g96zp
UklquUkNVPV2Vjr7I1dH4OdriIGKrqmdpxzt1Briyeo74phySd/tfwR3qnW23JcQ6DzZyKPJ+G1V
xdNOyVgXXzoeS5E6Hz4oCKDrmbQLSEALEFrjVsijIQCUzQavUhLlga7OooawtMkQ/SVN48zxBK3i
QuSCusNjD2P+HiB0HXQeEQPId3LU37gV4uZGDf5DrxlM1P6Un6KoGegI4zhkMJezyzdSn47JHdoC
qu8wofpIRO+hCCoqqPzRfy7G9fTfUzFOqxatmAhWZd2Jr5uOvLG5NxE9Cnf6nVD1GomZZSHaTmGo
eABxOjEEZgSH5mUy2lyaP+7LjgVIWg9Apk4xyPWQZJcAplVMKu9ni/z1FRWbdF1kmC+EVsiQRmYE
GHvo/1vVYmt7VXl0hhEdN7zEhnu+4FocaPbbojqnHwURZ+AQUL+u5Fsm55Pa6YQ0fXsgJvGTfa2J
DZgxMALyOiyeYdvhJdwoGxWc1GnjQcRl128vsxh4zqjgt9oSCLubVyAVyriwlnNc0m0mlSk3hzhs
o1SOD1ZeYHB4PdJBv0R9uIP37keijI74m1I0CuRaUQeTZDX8VSNhyHlt8u50ZJzWpeBP6xmtahaP
TEW2W8T4o6KLwJZZ2rVS2Hd4jcklB7bbws7cMKppY9CCLMc+8iK8p81gDIiIMeC3e+A/oK/GGESs
KpgyAjDAQWQUMD02nqHDpEuXW8vNXCs5rpg5Nv9UcfNpGUt1oxlLrg+Y6hSgzdNK2sw01pvJp/yy
BHOYT5oES2jFLv0n4xQdjnotw/vb4mRtUk0Bxe91AWBgvRoFrSmI0QP3QAx6uppv6eooKZxOLCnd
6KTWxKasQua54RIYMeobLatYMloNtuUsAXjfTRP9xN812XnU8SjurjO5IdBTitTsARVeIxI1Zeqx
7Oro/0XB3vfOcOoP7Q7ty9J0EoptZwS/9Zwuva6SbV1iyC9wyzBxYPGTAsHkmrnwttePXpLTLuw7
wY/TuTx4N+tzhAydTkfuAnIV6jUKzaJvnTX+iFOpnb2Kq57voU74urLLeqk1ZfFwBZbT3s59d7x0
ySOMscOov34V2qzO+gDQ3xNyTwopP2mJnbVxjTrrX9RP7ZIxW88y9uW42D/WfBTbU8ySs0AJHg4C
5LnLlTzweL4X6GkKzMAyJ4UZzlDjG9y6/8n5LAKjF0oQPA1DkJeg70IJJGFS9P/wL0UgtGKk3PXl
O1sU5pQehqF/2Sx6OUv7ZiPqwmcw2fW0R4vlaOTX14KgWzNMMCWwwgnCJ6jlbv661u5kQ1lBD06o
ErJdUD3DxHq4KbmUPylAmqvmgVDj8eykfRV4XeAKWlmAdYrqiRysGtUpPELGtYIB2zungZMlHv4+
J9CA/7qYF6VIltGUscPhmSZ+DcUpGymr+gNW4ZAPO39b8KWiv/S8Q6XcphQIi/IhkYJZ149qfeaE
sqP4WjyfjFDH9uTiqE/v/12lhx6odOrPG4OHJrGyxEne6PFzgrCAtbVQbhCbc8fbOwmO7ErWN5WD
PF53E9a5IFS9mLnrqMds2LIKSUJ6pdrX4Lrp+od5BwYDU3YN93ZHcZ58EUHq/sjFXBOFMFRaTaEh
U1Fq6qCFVVEIYHpFoASxS+ordeMVlsW7wV5NCLhA7SRmjSVVZWCtATx4plrAJtxVdL6BAXsHQMc3
XmM/q4fmVVNq93Vj4HP8v0xOCB5PgEPTnWet38qOxdIMTppxhg8jcu+bCWLuwymevXKFje7XgRSW
oilEuZppWmjONquz4SDPzSYDFn/U6YqumVTrK5zEkB0RAlGSfxv9lM8OqDopUA2eqsRzQ3sVspKH
036PhEwtIfu7kpKgy35kzYFUy2oLZo/akVVlvEoGFTLKCIXAJP8Tymqq5uoUfm995ot1LYqJQZuQ
zY7Cwd8ldeEbmvQwd/+x7do75j1xlZSYWHnLZpwZzutHnT0nfEX3MBO/5XRkwq1BKNi7zfNU+HMC
Jol7/7bb1S35l1hPstPrDa8vVdO6PYMcA8FWLQvmP+SRqkamsUkdT+Koql9HNNeY4M8xzFXfY8yG
ZPdlolTIGHObCItgl1HGrDjTjRTDijbPxhV7keY+KzMYcSgR3e2GpL4z2c/1qakzegBxO86m5ock
/GSQaz/Foj1zMrD/5fGWuB//msIPkqsBiLsms8GYrB8uqbVhIbP8qifWIOOeE9H1m8YEnLZxKvjV
zrIIFXGgou1UPuWbieuxLxpJ5pjUUAmh2vsmBEPPfUdiz//JRRts53YX3kzU1tk/M4wkvi0YB31P
Z+JYrYfbW7rDn8Rp2jO+gz0L6YYQgPJ+6M4G1+Q25hgy/P9hkpfWZWuhp0Ok8WIIa6ZHm8p7RqMd
SmV6YQRqRa2lXxGvSxk9Dbk9G5d/3j2mbJJWZk1YAGuGcuOhXb7dLOYuhBlzCSh5ICEj7y5pvkk8
VVofhyPkR6xzYwiS9Jl7i4kVJkx6CDXYAkC4krd5fwly7PxRdFI9yZ2ar4q2OpKxX1EqVUXpmYVz
99WnBgWrSJR0IhmLrlBE0zW9eCzGhmcez7ajkj49Bkk/6VJwi0GeoqVOieWC1lElG5N02T0K8UD6
Sx1UnLOLtVQtdwDU1YzoF3k2noV6EP7P8tuxak9M8WpTw14sEQ5H0g6m8isySJBuTVwZgQPwSvLg
HEMPCubXln2Cl/V+mKkkG4B4mpZ9ot4HtQPbMrVP43PsghAHUnJflnKsqANNPQdqv4cm0QjNvYhc
E0zo1SCZwtSpVWiBsjIz+uSzswvkm2W1Np5C/yHYe2yJYJqPWiMzn8Fl73XG6+fXX68ZGv2i7Dqk
ehvV0ej9JbPB2DD9jcT9g2h1hlWVTer693NqbNsavg88TUoLAVLe3zeRkHUksxhirlnvR9xSmH3C
4neUcg404S1MK3eotaYZyXgDzsREUWMEBXn2MqEVZt5YOZQOSAyddpISSfJHd94Ye0hknLLrLMbG
gBIPrEcI8iO22jiIaD2n7ei8mGdxxXikvqCMgZ/h0XMFqXLyIQcvM+JcQAXdY0GFlrw/gxpfK3Xk
xveCsNHwh9bru9WANH7WEkUY0xdTdaqciwlR1Gbqkn0oAzwABV4kWD4m6EbFqA/ed/CALC4pXMhe
cVk2oWVM13sA5RSMc+MhUDeV3c4t/KQpaPXABNqkt5EAiKz3r7pXw+3Cz5/XWwz7yFHiWXrHnrcd
4WbiOKey+KnBTGAbb3XK/amNwp1peQwcsNK4XGSXpd0d45FEOc0J7AAEClKe0al49tyl0xc5Zbzt
PAhoWw6+8zG7uw5LlCpWULF5OyAxLcbGMIKj40gIDKftQlNcaxKmDi7ig4rN3QpJJc2lg+zC/0AU
ToLP0udvvhaHxTE1qrWLYohMUvyZOzDnLtIsDb/dE8zM8L0X+wxy8yqcAw3sjet2d7+IuyO9XZFB
vX+h9E7VGmcSg39To1fUuCFCyZutwEgSoy9v82XpIGHBsBRV+RvLvxhHFnOz+02VafYUgK9fSKZ+
vJMMDjPDUh8zycspoMzht4qkfRGCiFftOLp01oulsEbULQlR5G5nWvn/2wxlmkAWw1nxUXXPemz9
PjkcihvvhYb1AAC1k6O6QaoU5tPr1dRoYpvByTjjQ8epLPQRDjaWCRWENe/2qq07umplhq98pOlo
sTrL6Ttq63CssjFiOuBP+5ogIEFFhSmv4zUAx7jj5cr4VgXdLU4A24bhdKdl0RGlOG06zPV7z5eq
wwdbc9AK8c8GpFMj/OW8UaeslH52sDLyg7zg6/ynnvk88XbQvlWliFkMIlHFyK7NUVT2BOuq/P10
QyNTQtRXqTufxtX8G3UQfBFXPwqF6/VNgoAe5opDFEM21fGXuaqRhfl2OvbbN9gGypHPi9fySfyp
7m2vAGyDSSl7fT9ksjjLUdT9NxblzsUBrawV/l2Ay3/MorAV6nQ98XYey1iSIiaKehdEC0DhAMMV
NhaSbL/eyp4ko+n9f0HhCS9roOgu0GQ5NwOekuFyatoJ59XU3M1//hDP9kJXyEiwhIbjmAR/KZLc
hU7lhtOgjCFNW1S+foA0d3VLX5fv4fnLnlRVEKGIoYKDV2V5t6A7SLZNPRoNcnYVF4B59HVrx44/
Oez49ehYN6iZFqT8T1Y9E6ICPN978fujPkgL+960SwsfFke5xYAer1GkxpkqxdMpCXZAOeOjoIu4
6LyJBG5FwBrG1NcRbxQJ7+xOY40ftrxMEIQQ0NMiN2pfcoQSaSjJ7JHUsPxXePzZGCfDtUUppif4
RWeWW2USvWTKCqY623tDuVLX/I5gMfS3/nKcC9/4ogRhVHY+PKlBRVyIk1T6zmeOHJcQnmef3+F2
IMMePKAEy6sv71TiLQ91l4JSa+BIxIFa/Fc9DrVqBhCV47vavI2LcUgqvjtgyoeidkcqMtHrcUz1
BrcGTy3pg+RQoHnzJ/Z9kkKWtfANkeCePlfMh2ml2aW30PmOHXDdTfLgnCCbXVpd7PTvFTF4jGeh
0l184q4nBvw/v6OCXCpLl+jNodHKMYkr6vf81fne02AdwBovJDFEIwdUyq0M64xdV/0LEwgpB9GX
i+0nmiXaGdWesU/LG+IXv8+DbHi8PLXIYx3+8ar1YBytwXfFBQoKYGHqBJSej2AByaflw/EQGwMp
+Ukz1mJFAwka1dq/mqTv38BX33bhA2OY99uHY5Pi3SeH+1VxgdfMq9SvJYLu64mwXvCSaQFVptyb
mzJLzigHKSYWooHb0lOoECxHHSraNkhVERT5msfoYC8O9BFLOJRpvtmlMju+Huqoj+BqbCv74opJ
uun2r4WSmoEJrCDgjEEiUTbVtgqYzBUYtc3SxzLVHEGV5lAnJYEqyAdlNvr8NexfjyvJAI/VHbcc
hExp15kp602zY1vblCmsvCxydVdSmuYWfz2ueMGxsPkiu9xX8dquYueOsOufpjmUygYtKj+qwOel
LwtHSwyFsvIL3B1lVK0RTCxu7htkL+ksNAmN1Fh1qXJJH91Yb5nyvsB89MW0//bNfCSOi7lyCI2k
zBFua52UYk3RJhM2MeOOo3DwJBp7pHrNXDDscdsPW2d7b5DmbOuRwzK1yQUh+K6C5oYAmbh369QE
r4mdEWerXNtj5KGDMiEm7fzI4CrHQtQLHiVK+pMxJs3zrLwVcqUlP2itmPCpUEchhk8B153ZDHoV
a7yUmS32wwR+euyX0Oas4PQbEolGZbk3z4NQBlOZADtLtFFAMCXlGhixtSgiCyqQYbF/3sX0c9PL
KmLwAv16E7vfWlE3FcIjNiAsjeLsN1W9l3k4cYdhtBsexoEp5gfTZAPMhzTkgD0TNJyq80/0UKys
UyuKFl0q5t4IeSpRE5eZ2NWQHVon8JH1MQ0vIOdCnIvN0CgeTNrmnOjMZhCuUg2o/C/fUYAzcNSN
vN0tTZwrgpnJTLYknmFpD1cFhziWB/4SnEdcTFrWAsZMybDmPZJ6AUYUCDFkAQ7ELUoRw4d+ADJx
YG24+E9N1fRuGYkiT9SiGw2yuDGVif7vYLs/6wN/Et3BJSO/eiYziII2Og4BM3FKfGrns6D89kQ3
wXM67hHhAPy+Xr45BcYpQwt6FricaehZTmmxF84IjoGuPOT3O6BdxQCfajMfYT5meleAttUX3clW
m5qN6Y1kv5WCOJF+SoxCtJeaPMoVol6OnX29+4rCe0uXBUH6+5uWcyptcWySBeTAgmf2WDNaoLTa
OEc3ko4S9RbzqMP7sCEPoHBSVUHFkdvmtNXMf5utkX9omr6dmDYpW1WxTpYjSx7Y/PP1d6e0k+SL
cj72iJwYz67E2osO+qS3bfTm2VylrIMUKNgOUhqU9huyGtVzKPWC7SWlDPb5M1rmyczSHD39wB1X
sH1al2dwbgWMpqT7H8uOCYNLt63GsCcCJBhMlAnl8yOB9FjQRkb0fkJUB2P7ofKo+iMzVVf30MWC
c9G61H+VVME26m7Q4I6figSjUkxEWYBCsj17B0p8sBs7AjfxhgAXBg5VqG8LlGV2dSzk6/rDSAM5
WyKbSHjukZO+9sNlTJjcX30qjum+O2fGf0WCfp0IvCSP4s0dPYyIQTfUWOAFM+2It0I/KD0xW4EO
IDBdJYsjEdIxeTjjMFKNzlsEypTfLijbnYZ5VVPPgN7mXJ5GdLg7ZFQhfhOYFt/VEtZMNXBCKiW7
F6j0tEIIhW1F8xnfpSAcPI+bQNmVYK6MbPdv+9k+OlGGllHdR3PO8gpQjeG1/5vnSuN7InTS6TnD
ZS3wvPoGnDM6CrZpo7QSDvGOkVubVK3ZjPepF3FWRP4CdPHOQnP3BcS7T2nj27pmlzP0kJzM1ZPC
J8OypG3h/BdI2Ti8oaFWf9MJ3zg+DOkGS2Cku01i3f/a+Xd9MpMB0bO6CsRo/f1Zmv3KbvMGiwFd
gF17buIykg1kjKABSPwgrIDYVpp82niJBTxxWvhai0ucnrFEGD3Cua8Yk5v8/O1pWlyx2JR0fc2Z
ZGhvlRfJBIuY+DAd1G3Kfe/3q7Ro0EVPdRf+UelHR5wGHFJxssypf7DvADNSaqzDpAsR/RPTbKWc
smLYrwZ4cmC8Vf2uwcZB08GVXIY9lGqWyV+38bGg6+q67IRnOm0aCLvbpTI6TtU8AZd2UvPtME+z
BpkqeGUhPuPZxk+T71zzeHlUET5vG/XJba9Qrv1d1CaUw1ZI3URFYBbYlHE5Hvmt8jd+SYSTkSyv
vbnxVvynfHvRGqj6Ws5sWoQuDz996vGaSPOjsXr4pyU6JJ4GDtZc2hEpfADFI378FdupU1rA+Ith
Nqn0Ck06xB0o2tfyeKeZ/jHhlTvrkvN2U8Xo4WAIsu1V4DkNWYLlE2PtOl59PGArKAo/d8n4GC0G
rV1622H5MagrE1nKwIWoKnNxReNN9xR7K3SDR3FUF1JCcqd/KOmxyDY6vJKeIpAKBBBg0E7chqWA
+LoXn4MmsMmne91yEguijfG7XKVtrCb6npS4J/KkYQaQS2RcIUMy3yHm6sGI0QA/WSspsaRACYVQ
zSSPtoMxsoXcGVzx4LvT/BRZaAWUtCH3cGIhO3DwGiJS17afKJ37UzLhSpHxTgzdqxxqm0MjrdmS
YSIXcHViU8+B3utrJz+0H7BnbHVb+l7hANR0VnHH4QtUCmZ+P8pvRtV11xkVwPBZMbEalrV8Mmqg
tzaiJ0GK64ovc0CrBEJUh9Zx4LKEkzuDUllw8iP/ac6mtbyzAIGnbDlad5FbDBcLehOno9JOVyv2
YNpZGRVUKcfqC8rwbQ2yk6ajmkQX3BNvCP4mkx9H2z1jbgCWJkVb1SqZuCB8ZGSFNj8Eo4khZILZ
JZUrPOkdaZHQElwpxHAFcctgv3W64CDtEwxG9mhUfcnQb7fRgJM17mj5n9Yp/rufUgrZNzwUlt0F
mebc8ihEOeyKG0pixeG6QpTRglSVPjmoRlUA8hF4Q1YLKMkx47jlQJ+r7S6vpQXdH0dGjVH3T2py
gAaRJZ9L1Mp3TLxCWI4vZc2sJptV3si+sXM2rQ2nsLZDU+meXeh39KGKWPRbmWtw4olh2RNg9x9T
e+mFSm0WIHy1a87oZLvRRfxbqmYN19m3/A7Mh44ohoQGTpbSXWgOw/c/Jb/qww5ctnCu1Ga00uH0
9sqXEf+yUUcnrnzE73jP43k8EiyAVrBKxWi30Tulp6rLZl3SGt3Bmf9D0MtCa+wJnT3pMG1qAjfS
ejQ9GhNS3mrJRsU0o5sccY4zp+I8NMXa5NjIyiCtzt5fnuwKDdOzJklnKfzAgmjvZvBgB1NAz+gZ
N86TskcavULeKXHreEgdFkWtcEA7WCkXLWrTP9BMBCcsTRAEUBmpYxm8KKUEPV8g+QxOeKDXuLFG
4JleyoWrtUvEpGd+q84tkkwyn7YC0c0ae20Rxzn3NQbbfOcnxcHJyg7ev3T43U3Ir3Lg9RS6HbGF
6c/sUGi2NahBnOQIR9PIZU+rC+sBg1uVvJ6ZgikCmPmVhf9VdzDE5ytIStIDq7GD0KfpIdW6Ci0t
Ls3Qg1sA9+DA5vWi9QX2PUeRVxu5PapKaXhbtTQipmuIrGJyK2tizU6JA8O06Dr128RmsTGuc2QZ
+dIEtFYOCidIz1FqCxyw3aXtLimJoRwMNVB6d7uVTjuEp/iitK58tds2abeE7208kU0n3pfJjNiz
DS0uDw6dOP70ow2+JktuuRifb01Md22rok71dPsH2n7n8TNv1R+Zcn87LAAOCLF/MNJR1zKv3OEw
kzWEDlnDRub0Wk8jHN9moVvzMkgofKCNKt7xA/zj6zwl5UwAixLbcW4TzGb3+i9GjyqGL8rlBhxH
2eccYSMGTe0/xGCgvVk4K3akMzJTJhisFfqcfL4uKIj/z//4keAJIWxtrW/ZQs7ZS8fj23CcHyHN
MhONrEYqEwKPDBO601zCazSei+9MO7/rqSuSPHUUj9VKQ7md77D3z7YOB0uUM8ec/AH5V1orDJld
9cBnMTHKLTG2qFS/OLpi5fQ7q/OMxhwjWb5lgmqJt3ls7DFTCzBljL/rLmA8UAgGrnpZN2SrpeEN
g8L9ZLRtVPS0PdLMJhY+7rg4HJTEdSjQ6usYQao6v83KOWsMY5ZR+FWIcE13l7JitZs3frwHN5Zs
8a9ZNNJ20EMrlCIAPzmeBqWGPvn0S8xR3F2zCIvBFUFy16uGAlPNMLmJacViTdK6iz1CVGKqg36L
P8XnWBF43lvAxr04TQYbPqrhhuPiHQajtsDMnOdXQTbepKPJTDdpFwztBccXrX3EMaZ1xs34Xojr
BqrS8JhX4cRns7PXcETCI9CX3NQCvqOUtXuowD56b/K+1vxMhW86E5vOsLKBw4qVYDvGmU7lSUsu
qluJAN/NMM41gymNF/a9jvkJxCUmus/TqCOGwahMUBRRqAiitbalw3sJLmEtf5dXt+qJ6RkARrGe
/JFZwubDLo0M/wOi1zw6wBQqEATM33aDDIiazVFfu7TulLNz7p6ThwRzSNPQtPJfnU9DMosEUunc
RyEGIXJVQ/PT2i7kULJHpBvk4oHL/E3Y+xpQ2QM0/fGnU1JYt+HmS746+8YnIGRLGA5a3M2eeV0N
EZX5+Loq09J76IVKXiyzP7kn+tYr9dtEfRFvqO1lNZtNfKVAlfkyBMSxzFBL7wjdFn7hYXkl8/T0
OaIZfkPJ6s9fgNrGmCI5RRuFTXRD427zJrSsErYEc610KL+5FPag2qTzfhHB4UllsMrYAZCbMlCL
/ZRUyfsODhmKYJN6xg4Equ4lXp2NTHQpbAsFLx4efyoHIThDUSaij8lULklcb8SzEDMjRFbWgbxP
by6FArpWI4y0wM1JlAO3n3oRAhSL4QYJ6a5qJ0bw5Fx37Z8u8bt3y8vlCfM7vK99AqK0pDAuiW4y
r0hgANsDh+PCcxqMjgH4dXu8RpEiMYKsszzxiCTirnynlqtWl6FLe647K/V/coA5cYdvv1nH0zWq
1C1Pq3B9lUWJak8IIrD1boEaxUnV5kPQLr/FoBqOTIbqlG9qRMJvc0URdI6P4glZJPwTf/8ACm5L
ceuirCNNfVruToNK8XHTwH8j6zEBS7Pk9ua15+pI9uabHYt9tN57PN3cvGezDzG+djei5PaJ3xbp
iQ6n4IrP1+M3jfAURMful9ohh8P5yGrYAGjBYdOWrfSvPiHmeajRaPpMfgpyTd3W6AJORVj9ZOZD
s+Ux1OzSM72BMwG8xyicqLYNTgg66ya3+BtnotjMcMsVXj65RD6twW9nIzX6ZkP5jfEwqySvORmo
Sx3ATohA5FBrm59lOuVKCaIYKTAK7GBuCuTvAEOlHCJRbPeuwIJvSVzQFh4sn5C8N1JbQbVJYWsM
PJR5y7GJa0YANQBB3GxsLDT8+Q9HFhhnwQoyjVVGiq9GeW5EDgBIYtHLdOwtuSD9K/MqOP3M1KWp
AQPwdhygbgrB879t6QzvXh5xJFN1NFYwloa7oA3dBwLLnKO3Gh9EtTbBBa9OHX0LlKa2BRPINyf1
qQ0X0C7duOE1PP2K6sgxMwwe7dYdvmnTCPxM403rWxlW4fuboGrezzj6bmGPtkEnEi/x9RI4DxgZ
QoWs2TN1fzP1CQMzfyMb8D4r1cofRbOsAEYuY8VrcAaOBYvmupfR2Y90BFkovzNrK+KKjKdNrG0L
G1lZ2PjGOfzHLMjy5nDRV3rr+kmmq+SfeIuZpQbG+UFYG4iwpZDrByEu+rzQGAz4GndyfHQfZY0r
HIc+kOT8iH0aG2BKfSTHYN/CBQxoz5ZDjZXZZL/QXx3JGBRtH3B4GKA/c0ipDDN5el9fWwE7ADgQ
xcoTmPmSLT78kR01ZCrDTEsjTnS/BA09TfPlkk2gBmt1swsIdjXh6RaGBPkE0+WtlC3kxx7DPlEp
HSh6gAwRMsuG8c8dfefnzjiKbMPobbS0rxjJ8eoNkAcZQq2ru09nomw5Hb2UG1aYw5oAdLF8Xo7U
28xzB0egBcKaGgt0eot7qTDEMcvwBij1QeDZLelP+mxa7UhYmcRt3AC4A2IvgE5571uTkCUDmGqw
bZdgC+oCDwYUhjm5HV/pybTxHuAIBTCd2Wskxk5RZkFkwI8H+l7aSeccMMGQ5N5u/36v2ap1OOuv
fkMq6vsbQv2L6mXGNNM/KcYqiIK/0PN4iDTKIOEmNAep+owQe5qXtHQfmXqoVz7J/nNTiExsNTdu
eo0LQr5bt1Klkb11uQreZcoteznxc7TEGKUreGT02hWzv/00E2UOtV20eagQ5Zob9wjZn2+G9os1
9k7K0JBtew/A9paOjG+LOQPk0ZeqSQrtGZ+d1mGY7kUa3mFUntpL/iiqShrFufnX6nbH9jaW4lTU
T17L5YJakp4Q0vSFDp4AJUWwZ5SlkFMG6F1EBCgb0xPzBM+uhLoR0NaL7aWx/9eVNftgnovTNSEh
5uB/mQLrTrQ3+MOIGQqLDS6wObW7Bw8hEX/gWWPTp9uqBJe79ciydJIC77pu20rhZnCqhzl95bIE
E7C3N9BtHCfmv2HDgK5OBNH/xflQaV9dRTqKg8Z6fEAaxYGU2OuB5+oiTGGShyknlJjZ9VVR0ARM
bY4Di4FdG5VLv0CFhEcWqG28pFtD0NincqbN8O6z6ZY7FZZkHXmLSylsRbD7HsyJrrzDP+DxwXRA
ozf4Wr5d5Unwj4XioFwzE5hcmnljOzQfCGULeSfK7E6VHpDowu7n8AOtUeb7Ehs1HHDILGIyFNDq
IiB+o5S/Ar68EyeFv+EDcABXnBOwy1qojIIdycGK8Q04a2qhDhWkbpSNp1yDsdBBY1FoeUkKkc8q
HYHUYIsO9yv5y23R8MelXNLXdPl3ASdkDTn6Flz4EvS6GezwEXbldFWP8A14yifoq4v5mOfF49h0
cuvpWCF1hlDQ4P2gI6MGbs+E/JTljVKjLy4OosA7TjFnqh7ZbIMZPQL1lPSwls+g/2Gyrg6h0w2E
WjpVfVeVT4XBGvc59pZgtdq4+jD+moMfMpIVlTQ6RGwnQODhtSom0xtMazBqqlov/jrHDcWZHMgR
LATGInTGYzbOc/xLMKVGkCDE1yQ34u0sMlDUg6plS0pWOgScheZyc5Or+TmZIyruBQyaFAezKPM0
BNDNAbCs9+pbH3gP4huDsck+1xJlwF9xclu8flaLHEptvsI46hYTpaHKMCE6gZc2jdcavxBjcGcz
rq1tIpnbuYDb59LHSBiBeM5LDj6fqQS88Lw6vnfPvLWOoKShvpP3+8Vjwc7hFP3JGL+Hc1cfNdxU
KOv8ACua1XTIQZzV0Gd+9GsgYLXImORf/WH52YQNSGxWeCsg40n21KUIDmJTM9nxNC8aRM1FW30M
GjpX9dnAtiPxQNCbGk7gV1XPq6PM62szn/DcMpLoKjmGpdqnPe2vTtv8pIdL2aC188j60ceutcPT
lNDIBzR4s8iaqAkBsA+R+v20PyFy2nZgKuzNPI1dXIRfkbn/+8U/WUapsFVPa/g5oGdlpHPlyEgJ
hN7mPjJCnO0RuBcd5G04G/EsE/Jdx8Wq4scoi78/Z7EYxu3wnmtU9PpBZywNE3ohm5LfhjEBQku1
ITDF0cZgrOw5zHfsBE/LJx3wf0cfeeV2ZGzGWUj7nUApGu2c9QUYKp/EAzH38Lt9ZA7zV94NHwqx
QFDTdSafHxgYh2rfGorALED5LIj/W7NKl4NPUCxqIHuIfCafJJTdGhmSo5MYB1YDT0ZjVe/TLGLk
hK67mRt3NCGILYUceUgI6EEwp0Ag+67IG0KF5RK3kMzCrAgYxaJSS+89hr8W9CGByhXE75qJADL+
XMp/3Xzinz4hHfy237qtASaord/D1JM+hJ6E3FvJN5Pv5L7kxoZrFO3ONyqDnlcEVwbLlXfsaSOy
prhAIA5N7GPzFfD2Ha5lzsM6F0ylzfz+i+zuLE9bNW/eu19WN3zw65QmQ0vCZjIzR03oE8isTDin
MgxLTv6wkMBFTyXMa1Sj+X9do3aDlVRSvN1T1LyQY0l+Ora/ubvoHK1aCYjNVk4AzKvlgaHA0yO+
xj6F1GgQmvxvoXWyVrluFUcngQMCE7Wt9IUErODtnEf79IXQuFFIc5M71P7fkM/iwlaqe12KoiI7
2YyMuapBs6T3TtqacCVd1RQxc+QKrwmEStzDU1sQKVkEo0oGmzOqP6jsfepZwBksDgJ56AqMLle9
ya/2US1gYoC1zE/m/y5y3STiHTNqsl88P8HF+AmofqFTzXFUqpoK0VB5F7klR/GF2Q5s+/ZaBGHr
GZcjBFDwvhGaJSl3sqx8K0Ci3Kq/p2aFzKPZG9QpbIKEAHdqQUqYsNNSAB1hOg5uly8bJWBg0j0G
m1qYwZzkkRh/KM8aWcwBwCOA0F+mpTe+GID5BjyNKeQAq9gmBWwvo/9kUxubTRA8qnf3DJ4+ZdED
6IN2UiQyS6wE2FT5F2LPv0x0xZrtUEhjRkuHhl9VwfGb4yJHzwGLUVWG/OyQJ4vQPEEdmqPbxKD/
xgP0ggjBBpBtnK/5RqWAbDffOtSSztSnd9npOSgKv6fIdZ3rvXM0FL0RgKq0T2N2ow8ltzRuD+8j
uUDbhhvQ2ew/YM9IHbsFzSiOYkdrn7Gg/QaP7qKjHiepVvBjf2xHxUfFcODsvbUDR5VUeZ22Oeqm
cJHU+nVMtAX6+G3wxDRZRgzWyQtmt1cArIlpK+t1KJqPKV3uPnIrOO4er/xlTkhe6hHzJvK6bOtm
nz5bu1RvxcB5TfOSo2oAba81oo0Ned2NaQKUGN7cBS+Ed9mDxCIewFT+RzyYmAdl3y6q3qHN0ct4
+C/JBr471Lh4ANzcRmk6rtDn+cNMAM8huU4/SU6pSX09mhS0IhE+kOnVkb86Z+w9faflRFVLIYVj
sx2MxvxbkzrLwqG5+QloCykS7Pwuu8onADnkYO7qipEVVG5kUhC7nNaiL+nlZX1kx1ZpO2gr3ILV
a8aC10FFQ+diiNw3ES9r3QI7kkwz+mVKhe2hMcPFXGrljrbWWnihJRTe8VHRW2INCHiLO/z7pyIG
9osn7wY+aMjRhp/ReNeDBk1EQAz11TFiblmEPSaEiEvj3RnKHgG57cahRJ+adXwC84QI9nMQRS7e
lnRkCpb6+0stTF6pMu6Dj6NXfYd7nRphPPTLExLNOlfVh7DO0qT/8iCWIvudQlL6IyIqxafJXjho
58cxwFfMFzssUdQSbvA05mwma5Bm1UOZ3yqAp8f3NZs7i9dyte8QcAEmoPCj9BgObVqMka9rYy+3
l+EamFsgLd8h6NGMvOWKqI4llc8EwyY0CriS8qUrrgM+6TO3uq4mfDoPuAu4OiF1c4igH4awZQ/3
jxSEH1gK+29gfRpP5gbw7pRAk3Ef20Dcoi3y46VdZrYWXVG+PWq9UVC4+EEy+MJIRqJiSf+XkTV6
klpBzilO8F1aGGcBrO3l5r2wa3PWlaipA++Wbj0aMI8ooSGJ6/sx5PXKr1/CuqCrPR71Ay9vmcIV
TrtSDZTDuJ+pUbfLKp9cPJZ29uARX1nzUfi6B8kJ8JemLQMSoVih/+1lZzrck1lxijTWAysqWXGq
RG3N0ETiy7th96eeH6a8UJUe9mnWnM4GVPlIXNlU7QLLHMwrH4Jc6pi5MoPekTEaZ+qFx1AqNxqR
YY+PWrSJkcb2x5xXdFX9J8TUmms8nm70nxWITiGqN6xZcYcojH+GHqv/62d+vJOL53Lu/80TmJhp
awCVnfMtZ2d/WDnWwqIpZIkItqw+ti91IV4fJIT88Qb5lwnu4I1EqbM9lONcT7qAQF1MeKOT/Itg
9XlgvEcT9nVGyTKtVf/xR6v5naF67lScnlsjIiPZrvqsBa5xhmTKco42K3zxyH6G7C/3qzC5ga2m
TK5IcVZKQEk4xK06RcWDAzdY4j/Hh+HlOgbs9Efhf2nifu2Ps9qC8qqkS++KiN9V4hkXfNrvGP2E
3odFCJEsRcIOF+KCO5xNlJeVdccNio+35YqGR5iW2KGF6X7wnH6GdIqPllnNVc+J8MusrOVcfCvE
ZXmfSPk2eaPWb5DNNS+bnuKSP5Dbh5FwvloYN/cLFeVlBFnXZ2vhe425eK6OLWjnG2TMZygA58Yl
3qhs+73QaxpNnLvD+0C5+cfuxV/lMvLTz/2yvetVLNAnmwEMpPuevTkaEFfKYIm33ElLAEB8Tl2u
xLRPTocqPwjAU4yiX4GZV0OtgjUzSFS2+4QQXouU4WxxnH9JuFIYyktkmtM3LE4kqQ6nRWkhSICv
xdEl0t5oxpg4IrvN2nU2r8+hG+P/Eif2R9nh1qrUz1DubIcre9lCmQRiCdRpRUIYilN0MHmuAu/A
lCVq8v6AzS0VzSHqoFaaiWmTi9afovcH7NlHJoCNmIHAUPRAZE8rguYkQTuKlH3Z5vlxJ+S16oag
Q0jHALrimdSh3GTXRFOGW4EhYyP2CoKvI+J+17RJtpIu1Ojyif/ttFg2kDOVuiWqs8am4MdybL/o
EYJn2owYMT/jQ+W5iTsURWGpeSLj8+Jw3bF5SdT53G8rnBHJhfHyGIQDDguFpEVEuvcT27COUqPe
N/09QkAdZ9Pt4FBCQJ13Jc1Q2qVrrTY2AUQKduYFHV0PS06sylAQPqaA8Rz4xqyQmSY/QYAcOQV4
iVRelfVg4RBgoT9VTqwlpFJkKp1eaSqXEREa12D9V8VEqr9Iok8AThNQ6rySOBuqPr8kPf3mLQ2q
nFhsgD+oHKsiz7Rxp9uwbU3khmzgKqidX3zwpEPelYOfclQUWN9j3IzD2qXmPPaUdivN3ZdT/aft
cBGe5zH0/DXCZha3bcKIkmJBsxwdX1G7h4OMq1Im4Ppvy5jrTar8UArSs0NLWAKjM8zokjckva7B
p5UcXdLymAxpjeWVJsFWA2kSaVyNgNzM52Z1Qj69Q5fXuf8Bkhl7NUORq4XiJMDiD9/Uj8hyH97q
fXHIWv++WRlesiijsNJW3uABfX88MJo/6nnkIoEV1V9ZI4CbD3iwjlNa65CTcPi2fPa2VmMbxbGY
n96qN+Gximkde9tZArXR0xWeMTpDzwwISWSGUypghut6D4KysSLges9p+AMUIGnwGv2LaCVvPeYH
6PF9t6jJ+Yv+we9q6FTlA4OKjCB5y1WkjHPJ7inEJrEoPuCXadw4Nbn8xgT3bZCf0m/BpwXO5vYH
hR5KXxnrKo23dEA7k2+4Ke7BnA5beQlBePAOKSUTMCi4Ql4YkBJDYKykajdCsZl4uxRsZXikpaE6
W1EI8um8HWQhjorTuttxqW5KAmUjlFlkMK9nF/SNBx+FIOqLo40vObP2tqz2LzWY+0RWjIdgOAtX
oMUkFhauiJYpHrFo4RVR17SG+4+ubqVa9tFP4vC9DdIIeMyD4ibyAB6HuYN8z/r4dj2vkHJlz8vx
Q61tOO6re9oHymTuHdUlxBAsxtQLfa2s2oA9pKSwx/KZAnitHyoMHNo9k4sf6GBC2Wt4qYfMcz/C
+3vPXfCmo3E2neWGCKL5vWdj2zzySSeNQOiejCLZmy3MO+DuKzmaHeAFTZ+vjAzSiyWtr6PGjp6q
OTyqALzR/eMggo8xUApY/qEh85Zr4mzw8u2hWXYc242fG9o1qa6S8SxQuHZdoVprKsDqJh3lsGNq
bXd2l65+rP4r34kI8+jyC0pMoPq660nmYQp9midN9g6ucDTecXI8fLM1an8VfiO9GFxizmelB+as
ePfxscZeW/eSyowMmor8PuJW8KdG/0yYm5jCjMPhm143xg8BIqJ7klkDmxV3+4FLw7OMNXpiZp1Y
hWlkPngwTSRpaLXaZx1o3QlFe+14wSHWVlBzLv60BAIgbUNrspsCTb2+UeKi80J/4ijcSOSIVlqM
4NVHh7AqC+NgQj8nU/CcpvXvCVZAo8R4LG4a+RvHK/Yt/4//9TiMqIv+Uc0Hk3n7ezdb5QTB/vMf
yr+8uR0DgBot+PFq3j6ApH28+R/7Cahd96DJoiZobCoGsTdgd3IvNWHs40DToLrF43N1b3poWM4B
ocOFLXNUomrGIZ1QbV71iM7yV9pikf9HL5YbYSr2v4khq+YjAw/Aby1J5Dal0U2LGx0qoUDmrIYl
/vv4eB3U3pIQSJYjJ+Z1rsjFHbRnzGCEm6Va56QrTZ/Wb0iNbnQKbnJKq4Zz7DAU6q8l8guk9BAd
LKx8D6LC1ybr29YfdmF0HRxyFknN5OkIYs+KXsHoFK7E0w/PBJYVl3QGyPux08x5UIP8sgjoUzIx
agRO0GAugMh3WgJGpCu60NmkQ4WCAGQ5+jlnPkuyKsTiT97wiPTWVJ2ZiHg8wlInP65L4EcxFhVM
vc4X5+hxA6EEVHTYogEs90P0czLKltn3OKGrCZ+Kk2VpqVhUFOUJQZfsVZ6VFZisWxKJ4E5oWvdJ
9MwjDntACymm8Y82Nx486rXdpTvqUIwWLMkghsxxKsCelYWNZDnV1pzh6ssgcCOSeOXSqQVrvB2I
j1/RIofQ7V26isX2tVer7K/cOuQkOI1GrUQLw1IcCPufhG4q4Y1EeJoksDmzYPQt4+wChWSeQcq7
lyPdVLyP0gl3z/Gk+GZKJQAN+iWbN8TJrvZup3YRtV28lDsnVLSpzdsdK2/tdarOcrxspN9XxUvz
Aar5bCZlYGxOGQkemBh2hURVMIEKQVelei+UPFRCwdR85BtJS0aBTn83+ijlp1wjgnkLm6lO93Ol
CcpJpB/zalKpSG3i09PqGCzNgs/4Y7aVc4l3t8j81sLeuKHN3rGwFmmuLze+2ShnJOOLa/dd+sJ2
rGrshApRrlQdxW72iHn8Y0EyQ/6kHg4o2yFPQ0ylk2sAHrZnJPhKSoAc9VMLj9hkZs01GAtQM2ml
vwLPjQY+hSu/nPJGoO9thH8ac7VUjsjgyBi6zxkY9Q0NmfEAXDKROjEROgFT2qFMwkz7tRv2EcgB
D3lQ1L22nqDhbu28nwRQWXSqa+nHy6KHc8T8fNZstX6WiH3b7HMXtR7IdKNRZi0erRDGxhgQueRu
ktT7SqKvHzybslw9H31PEipO8Y7DVY8KQOe0gk4wgR3nq2D96Sg5DFtaZFVbn/dfiboAG064Z0yZ
rB8Y6Ktr3aPfqtXnivcgfCLN6Unkl8R/kXMkLg1LahBQAz+rcxp9wWplGhWsndAwn4AeD9hjLsut
p+7uei0VsiK0CtdkqP/ZFw8l406knSfQKeNL2gBEF8eqxu5/b52B7FHmIXwp/1Rzg46b3PNcCw9E
aJVpQzPxRT77MJWj43gzn0joUPqK0xMM56mISKyrCIT9lz5Vnri0ztfNvZWOaqVxMzASlRa1ZCdQ
XM2vZppcOb8QSLeOBm6BeGUL4Ldnv4oujNQK+duV6nL3QzTiXjN+fH/XSzm32tHqfaRA6IaMditf
kasfjJ7bVNwZauSsCmxJberowKdN8XaBl+1PMDCXisTe+NOcpNkhv5hc6h6FCle1kbcyhsRfRYk+
8ianpNCH1SJwY4MAzkupYUY5WNvMknRsapZzDFfQi5WtNM3FwZCsEeS7pB0dmwKdWBo4Dli9vp1F
7uvDPrK3ps/NVxUFG56gXfVJuxlM0TayYA57DfLpn3nyIxtj4TGw33ggF6u91mOUplYW7DSaQihG
6GdssA2NCAYWWj01eANc15u068qziyaEgSrxiPWzIY5ZPP4EZOtcvccHmcx2vHRqQfPD6lIP7cKZ
B9Z1iis8e7OaDfAMugUVu5FI4M1ROSxQ2V6YSVS74KE89T5u1aEyWYn8SBt/sjTLT8ksJv3Vv69n
jR+LiyyjqXCstXvJQL0ZYVZk5weqHTkU5XPeHVIfpDi90kbLxu/i37Ez4+vl81ujG6/cJXWmWSa2
iVNBRXiLCdcfq1LppWgnl5Ym+ZPbIbkm50oI5lTGD+RzV7iLB/hD+poRwN3r7kYFf+AzxB16YQUK
7fZOKIFG/qyJJsfTPWpnDv9HZzSJ0kCMHw87FdiRatJPZLOw8Y4Vu7n/9fmN3MU4hcc64Th6tEoY
8gvjdkL3QhCSvZmnPT+00T7RoJYPL1hpazaPOyLSyG49fbETW9/ZhB6nOUluqGka5z9BenLKHxi0
8fRFh4roKzGms9+lr3t0Q1/MW3UioroXINPnFrAFdVgroQjxVy7KgwaBdrOg4MFK2jawzEd9CtmP
q6CMBB4AEjrdRb8Q+6bqo6ub2/oiLHiCkKrxRNqGc0FcTsaoVnnPmZ5R3P+q9cbkwvhkldgNStqE
kRkO3OIwY6A5xBJOnSl6PNU2vHfAX+eLRWr7DMw1Grs7OFflZ80uqcWSjwls414qZcLauddDJB39
fditIxvgdupxLLSH5sDJyB6gDTh5Z5uitp3h0n6OpeHU/BzbDfWoJ2yOurm0HnZgDluUWHOeE5dB
UjyYY0cVe0fgeO0UbiB+3mWchFBhJk3iAE5JRsfGtPKm7eAwK00xujMn/NK4zfIKJRSxneYh/jma
1p50VNAoF0OXrnyXu6Yk0lcsNA4Jb7l1onE0YPMPZfUl8OBby3PCuHzJ2VS/oc7X9y7lsoanugqG
OaP4mJxZAtl5VUhD/G+n4O/iLwwtg9ODlNDd3Pyhphl9rFoy2vW3lnjxrBvNtfh+IFeV4OqejE4j
v/Ob5g+Mxe7b0AaoqklHe/uq6GkV/ZOuDUzdcs7tXqypJvKOt6UcgLF3AHZYPohyZrljCpNoLUIu
Di9aYO9efMv3rGQTApaIYIMwJQIQl1FfhhfxeMdfZBcxovVDXmSmnxpzyq4B6ZojcU+hgvJLwcwz
KVGLptQ6I+NP+ZmBRbkaNhulx01i6tcMzotVR5nP2enWTsKpO7qQCRgW69wSKfQCncz8d644FYJP
EjyhlWOxNwVvcQ6Vn1EULr/Vl93Y0oKnWRgs+W7pDlCSj+5Qf9Q9wVOY4Z0eI7sgYBHetdbYuY5R
gzKYmyR5pHi20NvC1d4kELM3T49Mina1QZ4djVjxoGwyWmmti2o216akypXTcIZ72H35OknT6IUt
pKjOUsQD3dy4SFzRDBDq5JTnVwDQzhe486qthpTs2Qvts3jD6OJzBmpO58vyIF95ZQ5m3NTEPLI9
kNNRUD5HRRdDNRW+mPD+jBUlzgdYyArTwNBEbpe9/LTtFSDHvQvQRyl3GSR9ZNoc40bFXY3jRjLA
iUSFXdBDYhq71J3JVS/waNNKgWWXyLuPhV7oEDi3NWgVtVeG7dfWUvuyvQuZRF6MusnD8lAzqiby
2PKLgT4SOZNZNXMMMRp2jRUkeGccKCPgA7LrM7Zn09upvfwAtbHC0ZfGPUNS+A8Krv67N3EjX9+O
wKFYe8mN+fvzsUwYxdU4luQ/HwoTlo4BO+ZLX9W4uBpYa1QOaCb0ob/1RlUORBAKVGbOnY/YdhZ2
tdo/v+11uefpwWj/rwBugUhNXqqkEE1dzqOVOBk6ME2lSSJVdoqhEobEgTaWUswM8KSPyu0vddMJ
+3WCqH5avydale5eA7vmmTekWTyaXR0CEFSKn/CbTI5VLWiUWkHVFMnist4OaVY385yOwXwK9FEh
C/VBwkiOlkLkpTmvB5O/lVvE7yDmKnUbJmuzDp2gYQcS0zb8ACyHs30fOA/m5fZaT9OR9UN0N/GJ
Ycd1QK5dlRQWTurpu65DsjnGfg7YkK8UjPCagGmYn7Hjr+029m0dwUJSjWYHHQ2RRyzYosQgFhho
xckz1U7lmX4LRe7KN47fEf3I5A0t2r30wJvDSWWLg/6NmNRnOP11P1vohFsXvhdvZsEp3kL4k2uN
1wR1ilrNIjEessiEly3KdWbvTb6JbNv2YT7wxksytk/Occsg4spMKDjk3mmD1kVuzxD6Bge0FtO6
LzcKe97khFd7KCiqiBT97UzKs/8tjNDFp05uNXuJjaFfEYpFlYAWkh15bFAE9sHM/nIWB0nTfBap
1PFtGoxwj2V7nUyDW6EFYqcohCx4M1oEgcDy5j/ckfYe6n65UNSflk1JpyvsJa4CgVuAJiEjuESZ
Yu0JnYlq5w2e//0GjFan4iqYiDTV00NKg43ocN/VNX+bRSnDzeddVXh1T8tFd1pooBqj+ndtShPk
+ln5K2U5+AsY43mCnLXt0+smS2uYD/aGA43ZyEHwjF51fVNMGLzDMM3iZLM1fmmxvIhCgI7SIWap
2+3UYUsJVpvD+pHyvQ0UPZi5kubV/EQQMglFktfl2Bu9Rf56Xlu06AAWieoloMbKq2IzObCwHCU6
bUb9HY0IE4RAXfq59f2rS9sYr9O8xbLl65TP4698n879Xsb8rcojuzS03vKCjJwkDy/t89gBTige
4NxdUnwV/sKYeu/S7741SHFHaSpOeegAk3yzUkxEeFJ9XdFhblOxFvsO04Uw81MDXW9GZtSCBo6l
8NqIBij1JesC+f2pLTTHI06lRkPiqXWYszI9Md1i78/L2DiatNBDKGB3+XPQAiOXR9zWvVVpW4qI
mkrA0ofpwtEwd/pkqUbR8fZakGi+hiyb38GOBI5eA2Q32j8Irf/jByH46G2BqmPs3aFvgT4jR/VH
mj8eyHgMh2/20/T5aqgC3lwEeFuWi/i0g6+VnuS2mVn8SIqBi76miNumDQttWGvyQKsesMwGLMHM
wXwOHobeuQfRe3IbuYJ2ZB19W1IOGmOTqrvxajvQh2APwHyjNEl2LjiW5Srf82Zfyyk65/2/keJ2
JBrgWJ5I+J7qH1sJtLNQcsquA3l/CLdJdpn738x1yf+/+Yr1pRLi1ouM5Uiew11N6x7yHVEsgr+U
KHsM3OqpNJi+vWCkUEmwUxKo9a3cQNrVEOmNsS3hmVjUnbcL5Dqhn6KXBOr4J3Q4HZHr77/BLOB3
6YQTTmxA/NuRUdGjKZt7GRRtZyfzfz9N8nL1YUvuj1Z006Ne0Ks744KsnioXVHgc+Fygo7OouK8a
e8+HVB9+fEXVPpp2iAxdAVn+5vRPQwYh5WbkJEqfWGWGvs4KrOFPxwWbgentwZnAdl/n7Z7SQGbE
LJuM8j/YzPLK1M2t8IF2g2ZFwUH+gaOLwNAGc6o2nIAJdxm7Yki3UvRMVeYvSgwPnxauZ8v73RkS
9iW5UJkGwWkNXBrSOcUrcot67sVVN3la6BXgzQNGadZV0vqdaeanX7mGYziRFKEgIZQBNieYQckl
eY8aZooBHTz+rS1wGKu+ya7q6um25t1EOszlGdlbYoObnjIXg7oidaKk87uuVJPMQiJIcBL1HjQ/
RnVnooRdZ+wtU5F3UNAb0HjmEu+CSkEn+JDK2q23zytBChSXkR7hhwB6tMeRK8Vdo6GKBz1QERVt
RNz6lsAMV2Ff7gkjHYjVsR1kk0YwsiilLOA9aCYBlSTXXvUvm2IJlUJOSkIxJ6pplhGqZWTibRbz
4EoO8EQ5Z82lJmhqiSuuK1Br3biK7bN4izXbQYA6DE8K1np8+qMaluygXWKaH68mfQWpsE2lb3jI
c6tHOO9KsxKrd0DFxpTHRDte35Xio31MsmVwE+K8xrKvB4WCEA0WVp/jeKv6F6wJIy2UA0BlgDCq
ZBrhBrvYEKR5neT5t/LpRIABstSYpUFQS9+XftVwlXmxkmmEsnK90Nssb/Z3TaiWpsJlfdUxY1LJ
Io7D/fiXnXX4jx8OST2KXMNGMyfSx5yUl0/dQU+Md2ILvXCY6Gm+vvZf3Qts8+WCLKYLclcWTNzx
8biqQ0jdrMk0s7C7qgNdRL5Az81xY+2EMybAwEMP3Ht7fGi/x8Cps+lYvmNmS0KjT9IJHUDicIaa
SqAZhb21Qw9Pj2UCZEqmcF/j8fZQyXnTCNMZd9X+ry+dL3mgnPTdAmL8BxfeBs0pFxLQfofk8TUo
PEkhRavxtOURKrqC/1rug3nyqZ9CuMf+nb8T4FFR5Ky1CACzfThdsQGRjF+lxOIIqdfwmZdqbSgz
KsdTpa6bcSgatSMziya4vEIQPxIpgEunj81aG4jntMae/00MITO32/pkzKD8GOr1ZcuX/cWf2eJZ
QqvfjUU/4PLXfRCCpCo+Ue4AE+k3C0hTykVSp144e4o7jagjQOSycciqJ4mX7jwsvA/jMyiDzs2F
bYZjCb5YA28rJn0yAnasEb9I41J4WjgDysoiaktZtrlUgu5RoTpylhqLIVf+qpQwpImEMUZPn9H7
zhbONKtJRHcUoMoiXX5z4ZUHKFsiC4YEsWNzhq/zdPpJqhKzMMFC79SysVZdlOLS94HlWOsEwKO2
j4DbgaQK7R4egHQbF3Xbw4leitqzE54UI5/0KlydUIyxbhhxBqTOssOwXhF7pMpb5NbVOcMqh87z
pgSTC5KNsKSjkAwESGixgG76oulKzFqZfGoKVUtZNaaMp8l9N2EzDcoxq7A+tbI04p4ATjuF2RW7
wAvAO1Kf+gS1dFzLiK5cx0yfdZSrPtCaKFVIxXcEjQuiIhfS1/z3SBqqEYQaeUYN4zGOUgF7rMzD
68c2nQkB6sMTvOelpH1leRCefRa12XwTcjeAONX6AQY4J7NJDKzSowc/ArTNhnAqmm5PMAYgptX1
kohZSyD6AJJtaMIBcLcRXFk6gpRs4CNukl1PkWTxwX/rP6QZvNGSRIfmoiRXe71q8RTLgS/MpcHK
UynU3XKa7/Q09xX/2J9Rwq6EBtkqPdHD1IVp0zGR2uUfPBWZfnkub3BYMN+WejsNHKVU2UeVnuP8
Q2XSMYG6m8pHXXurHX7XU20q6cdQjkBR+DcPEE6qNJY01nOcsarwghiX88KBrP5RrIu92YRxTqT6
Aiw1AEFwmo5SP8ne6n4njrbCHmLKDmXjh01PZGaxPHamMDm9r9s4XaGEPUfRoOSMgAVv1y8Gw5Sv
wswGJ7Owemd4vomIjY3ZZxBrxoJ7WRx9dgkW5B4CNPGw3VEyyHDcDl7ih86p+t4SOTyLj+jSRYM9
cR99ppUUQtakt4byZSSav4hmARPrAL2cerZVRpmOlZELY6rENvyiikpSTjI0A6CzkReZhewNqUne
SBqoMX+UisJo+hJ/jPBzuuC9j3hSQL263qXjgAC5DxAxD5zVtgqQKXr5BlYTSfqn8h5CKfE2aECh
Os1qEJaL8IxkJAKu1OOsjce6DPEvNAAC/TB4IgDiJPI3tpGbNeliXujjuuTdPmnIbkUXggHgCfbP
+pLulkQX657tlQIK92j+2+KHvybs91V5rmJMa9vactN0q9Fp05bwQ5J/DzeY3cNyTVFMplVoWvjv
7SPdIUcO07ii9JG6f6XEIlOCXNGKt5+yNfMpCPDaYHdLL2FZGBHYUqBqVMcPxt6RO1NE3HlD3vEM
6qt9kgK0mUL1BckU7oSVzeRVNCFpW/GRUj6p5OkXpFGM2lt6wNXor5Bdo1ycn7NiIOcXK3PRGecU
h3Qp7cHVOEmE54yjZql9rIWjuXpFexQNBw0/DQUFCVt3Oi7ukbJG428nN7Bc7YQSSdsy5HezmcCi
Iyg42EXZAbnLtZHisrboDR74isLJMFlZ/fPlRzI3vbGWAOn9KjENiXv0Fqgn4DxpjxT4PPmk1h5t
mvLJu8X3UIw02qm+1FQ4d4qUyJvt1a6qt38EKGyLUNRGYhcPyLuTeezvA5S5itd7Az4qibUme3Qr
O2vEwLvO+pn7qxhpSvcn4F5WG/EVHsqKJhlAaVeDoVNaEyaS5y7LivxF7QspQhu3rCEeZkjX+TUh
7azwJEezm26h017EUo/x/j/W6G5akiH62gCP4pYB6oW53VmahrbFN2LfZMEqH900/nZ9v6zdxcFD
rKGZToYyxTRl0kvYbrwMF69c8Q9w7gWm2n4xFHjSAI9hy10WDN0EfTJu2WdskGw2mKCAnX53pjT+
G6HhGvxSI064b+Wi+hluNkVBnQGvXKAmUOJkCTyImGLWjkPBwm02aw2IXlNU+vahfMEjGNPQckSt
ZGHxRpYsFL4jLyohzgIccP/FBFMFM1nWO5MunLDZjZPgiWxg/u40iBEh0VT0m5qfduPZ9xHabHnC
UQYf/TGiX7lIw28WFAWIafMQfPxnf0DURyigRbaW/Q46XSHH+pDg231jrSg7hXAsfWKPV6WKWQPF
/1piwMn3ThkVal46NmFn+SQCG/g9L/du32ydgUIFho8B0uFj08xKFOBuFqSYU1IyC95v9GCuNvXS
11Nj6Hw5G8MX+wTlNrgtbRd8WvxY3fNSU+fXnYHoSVogluLTRaB/AVJXwiVWMRhDqusG1c16iEjD
Bnmdhd1RvZcecf44s2uyj3whgFTO30ZeILk8ZX+2WE+BS7JDIWZawd+2lPLum/7VmA/3juOIlBVf
7R9dsuQZmT/csRNaISrJcqCXpb/Ni2AgEnyElt8PqC/ranVlMIf0O6PthN3mYZwXr2+CZg5WN8Gl
w3M3Hu6l6wORjkmGaZfgypzSm9+df6p1EeGeSSVLKnd2dY4cAXGAc47huznAmvUJUJsGSBy8/lYH
ZofD8iw7G3kQK276Zeg/mRpMekjJ0gwxVDfdu2tUY2Sqd4coHvTUEZ/LgspasucAa7lY4MUHC5a0
GJNSJ6QzserNlg02cRGgMuIuOufsokPz+ptukQi3f2zJRrw+8DOB6imolL1ui5LqOP6ip+87iCk+
YzXSO9SCy/1KtlVM77XQDFPfeThQfsX4InLQk0fJTnl/4uEN3WQV3NXLH8wyPnda4p6PssDLbzBh
dzOCNNNee5S8ddvFf5JfJo5pf4q5EaH6J27luZR5p6ARqcOHpNvT1zhYuFk0S6en/UTeMENO+A76
vk0RRpO7x0eUK+5lwKJ6Tf54k7g75ajYDMfLShigBsxA+TEw3JThHpiaoRcXb30/JvXcj0QuPajj
hCInflRrF8aJxkeEHLhESNo7hLgiBFOEVrBUYTLljxqGsV8qjCP8qF0FOt5kv9YSRab/52mMG8ad
eW5V/ylt35kGJD/0Qd3cS0W8lwDG0rKRxMDcPAyWtiYY6Ifb/v6oRn6fivkfHNNQNbb9csDrHQVr
4VnU2niucz9RI7tEgkFUhlc9EMYEOWk/zVEUiQufFfQvB04gk/wqsLIjJfSN8nSfg2pOFqMWKv17
fWsRJZ27LCFrUsBqkBxLgnpEg6ydy4VFkmvcO7F8IQ/p2jjnq1U9pre54a2qQ1l1M+3h+ylMj3sl
HOnvhmyP4D/VEs88hb9rzRhnM3NaT9VQTWxQNCUd3dL/cV33WxH4OUd8RAZTw3/m/+S42yBp8hAa
mwLS1Igm6OUETG+5qF1PZh7qvLnQexEctvXrU+ZY2xOBUR07/R+lYUDgfFHiQcO70m5bP7xIQsqw
Q7HxIh8pUC8S0mTYrYf4NNsyPclcgDuIacjVPHn77rGMguY4QJdtMRAXaiNTgiKmmlpzjiT3/Wrq
5dzN0324959uE2y1QEscqIAXcOIzgFbJl3MKJM+qazcg3SfGJRJ+Q2EeNoND6hnMjoKDqgS4KmRd
lOHq51jCYlltwhT/I9TlCMxpdnsezG5AFuSxTFZs7ixkqNwj1wiYtltEaMzYKsEnOy1cBRc4KeWy
i8nS7eS1jAnMiZqafxo2w9AUdKueicUa2LNpUKa+DnVbs9SHU7sMHE3VbZQcHBkEtlK/EQqImEh0
Kk3Bl6joNJSpEYYRGntMn6Ti9zj+qKM4bOsMJKac4c/neGox17mqY8HIb9fUcAA5VBzqogX7H4gU
4JB/Fd+VtwcUxtxcp1fDFzbLsYpdiVpqg5It2u72FcLn56MOx5xb5WXzLWWRtMv9dFNkY8GSMq9V
r8YV7qEtKAduQcRopX9dk9/lw1/4HsRYOnraOWZjz2j+zvzMUA1UlqVjN207uIislE6da3lrkpV0
rz9aSMK8Swf6uQzu9vMAN9MmS+sfQ1dqF3C+TufmS3JrZDYjfk4tFIkEgEhfkmG2p3LeZa01uKla
FbfVLdT+KHbPlfKR1UaMRBkXSDyzy/BkdWYH6J69CSCmSp/nPeK6YFudqr6xewXk6kBOytlf1ibv
Vj2ecyc6lmnoMcUn4OdTDEcxUPvIC+Fu73FIS42Re4erEiYa9aqKmnH0bhq5vfcx0yRlp3Ysxvud
pIgg2RrXZLhaN4wvGwBfCsri+x5FhhrYUuZtyQ1qZXrSnNwjSeA+SZ7vz1hxfdealjBydEpU9T2+
Awzh5YHg/1y17ia5rvxvUAuU2tbmKCU3cEUUHvJ5pUG4lDDfXj6UVLx1KnUGfgRqj/oPuWHiDyOo
PVjPaK0KtyqTbv1ZicSVTuWYVbOmKS0Y7uvDir/3quBBr7zCt2XTAR/x22GPuVXqGYxktTSatArb
FNe0AFswrVtDZd9lbxo3JN5TZgwHGxBEaAPvYqjbfffxqUMWWHqXoAnIsehLfwE4CFGVdky0pMOt
1b9yGu85SPVifeQGjLbmB/4TK4Thm8usgYhA2DBkmMWFGXizaoOXo3nuTYNX0B92UaYcX7Qa+WHj
Y82RmVp7CK+AT6onCXUfC4YLbcfa7XfPDfXnixwfJzNNyz18wi5xoJCuPe79BvHtQfCdH7djFhQp
eMvSBdJm6xDZMdezOJ2UqjIxPjEi9hdElQVpScOyBxi+PDpu0SoTEVT9/aCB0H6rm4Rf1S5Z3rjw
KTkfiCl/5gObJXLjPFgLsg9cvF8747wLE8WVSHs2Vl3Yfq0meXYiBFrXBOXAY3XTbOyHA1mLs4S6
EWNOu6dqo4XZ8vHs2u0eWB/iyCCabRpsLPkPLJ+6aTeZWAzV0Hs8f7AfeREIgDN4tSpjJxatof9D
Q7eRCv7l3dwryc+l8Pli/Xj822oh7olzMTlVCUllD5c6YZr/nD3WQ4S8nts+dhV41Qu6/ucYHYlR
TjvNfh+0NWS5OosEkV8YQ6KjlCTjGjVMYcCzfX6FFA87Ap0z94ZBLyP85EjKsM5/gxAdR1VNW5jd
On0jy0jhHJLsh2Uhu/Kpk1REmlFFheh1e3iousu5V2iaT3citBBV/0237av+El7MQqD8/K+3V536
WlgW2WkUmcG8YMUiLtrsrB6gqJMpikMFJ7SzUqSxytMUeiz65Y2vi8KcmN4GE0o2OG5AaOSSbXJf
NnlOBgQNoe4FeDpJx+psjH4KF0TEVeSj4Ayjl9uN5mBWOuY2JnRhXUDyL5W27evpLgr153s95lu0
y2LZht8MQFL2jUxB/eBxvKUVW97ywVzCApR+IJQlsNhx40hOZeq+mRwPN3fNMxc0c1uUT/1Z9WLy
L5sd/vC/Hwm43tzQ3g05SVcsuq0r+ELB3+FmngN3Cr3D+oqBjMPvElUJxWUjhV81CC9EAkDQD2LU
t5+7a/VwcF+Iw4i9l67Sa0kQU37v1+UA4CLfu0i2Zc8tXIiDkpTwYdIVUAmWlfWIZN09WO9KpxSy
F4keIh9dm4PcCTZtB+qUY1Gd/qdp1IRqOAH0T9SWED/3ZjD5gJSKxDgRnRAPeFDNQIqHrDpNrr6D
eNJe94U5RR4RBW/FmJHfWxEizOlq66F84WA2p87PB5NegkF9GwhD8PYF2e3PELquUSBveVC/ovK2
gjsh8Apo3abk/nHEOIoCMb0LmWGlDYraE27hS8wwmlXaOxe/rnFZTI5HY9Mrippiuv6vfU9wqzoi
5r1FmmWk+N/K8uJR03/Tv7xbnZm4UyDfF3gmIJatL/D6MCEkq3qizTxUzKDK/B87OebqR5HaUbPe
ojX5Um6e7ieF/5paoP78SMxbxD1FOuUEoXM2Db5zzhfM0zMt3iaMgZZXO21NXm7YqiO8NSfZznmc
WDe++Bz0T8UGKpI82SFBBCeiyyQB37g3Nny9hSsTOeF6Dc9FSL0PjtQkBWZItGxFD+dA8sV0GDhH
q+Rm8wqVuicy29976oV35FCogeSvLl2H2e8r2cWN72r/ymBOTg1zLPVZm9oU49PE3WfI0BLmoN1V
9v7A1Sktod/ICKjBJYu4HqWocOdUW8q1FwHwzsTMQXi+T0M4Bd6mns0YEORvbo+xlWh7lp9MDd7j
Kp6QJ3GOUCGgRmBAswOYLbsx+2Qy37gLRHNTJz0BnOQ79kPe1FeqwZ8jfwkWUoG9HyYCm3Q5cl5x
sPGhfJvljUNKQVON8lYXfHdw/6NOFzDyscnyLB5mrOItn336ifaFzS3mp2ezi9hdCIVGaPAEbylA
I7pSAkQTePbvKVOhfKl/m2pHtnaDSPd+ua1fguJ3fsnq+mq2VvJeOCyLv/RWwl1R9bjet/KgEIKq
QVcG05cTG/NcZJbBHR8caSanH6CrkuMkfr4Sb2iOLlWhr8SjaDafRoAZmTq65x06CFr3lNDh/fG+
FTfSIBgW2hih7Jae5ckBGG7VITvoPh7U+2/r5xgVBrxlCjvq+IFh4iSCl3f3D4X/qpVrWPsxj1E8
JpmSkZN2vEdP9vezyNH9ya8KhChyMSXGSurZsbsSAis3/pp31lxx/thxCCn92PvLvqHxAiXosX/+
r3BqAWMI6hoFf62dlxB2Lnbjah+IhKUB2ltEBZcKFECqQeYTt0AiXdAHxszBJyk0m8YB9uc20T64
yH/5j2Z3BqrndSNukhQykjqEcrvw8SfP3dwlVqO5u1faw8G82+hLZXOtWs8HiIJ7Ar8nbwyLHADH
1rlrFZtRHUdGQZ64besJvjsAXzW7NJqu5nuvh+rv8CaEs+P3ZaGQttg0OwwuxNLugHZjOSh1njtc
DiRuwNNM72owss9lJYVM8ODVjbnowSmv0oxVMxD1OjlcpbD+oFVSLG+m4gZaSUwYV7u8VKmCYYnr
+VZx4f0PrMhKqWtBLe81mDXpqBwxD2B43BZmcgzcZNGJsBALi4Ywjhw3OcD8rr3VDoO0HbPupkN4
H+tunOAv1RQGBEA1wdUdUDMrPHkSiZYGxE1wo5cl3kkq0dqjW45Yhqh+d1toue5sK5rmBF2eguz8
NnfT19QnMF/+JzU1Wc6u1NBrEwXV8j6ZRZdNitB6aFFV3pSNa6pOKeIdizrxc1+pgJBKSZy5/pk7
1z467oDx6RrZzNAglysyHpnWOA4knNqBJmzNf0M6wjh83OVHHW5cAbrlGwlZUxrBbbfmemNbB3Au
rwQ0zXJQWfeQ1cB6uW9ItrTTdNegVwttXwxbts77Vt+bUmMduijLLJ+mhf/Oa/WLygXBAax6xis1
1krB8Xcwhu/hEtfQZ7iNrTcUpsRzW6jiSxaQRnBB/8CuaomhES1QPLtrqXwdisGJYQ6WUTpiJOt+
1Rpk7LGR9thKYGktc/qcBgCd6xXXxavGBs8aL6Fpkvs2DFWEymWdjDFOQ/lyg47lD7I5Ibz4JwbD
upv1RbAix3HUc9Vk/Hr/xscyn/6HELRd6ICaVn266qokqdKLsEKomQeZvqrvPCYcCDQ8+cApb/Io
kecXlhu0ddSL/b28Gj2rCuVjoBcd5ZHt/jKqGbw+mdIUrZP4LJrLRyjkLpuVz1ptZXN+WRD4tU8k
vymghaSL7PW768RCbgcRGG1/VjGijLKNQMtNPPKsS4/FWvIA9uZg75S7JgwOLhGdrntQXVus/38b
U38iTEv6Xf8xC4d6eSV2ehgCh9/8OBCierhzdsCw7GnlW2/1mm661lYRYXOiNsqXbammUXTe2F4p
W7dpQ/WhDewrCA/UHFfWvKO3yirM8Xun2Kz5/YT0NdZN+GRRRGgHCOix/qVpqYfSXrqLILc22MJP
3zBWkVHaqal+lXUPzChvXGoKbSMAoaU3fHZ5MOgIFgcXQJMEbBNUrIpMg1+FJlef72lti+2Vcm3O
B/r5+l9QTtotvhi9/G6cPNtAqOxJyqqZvgdDZwzV/GevMZOVqKfauikYVY7ub+XtT9Tcd3oArMt8
pF7l94VUsb23IsqZBd3L4a84DT+ycO4HWRvIUJtdw4Ow54us03GKT7DSDhUeZ/HuXVRTDKqXPYkt
tWFxMMvU+1YrJ71QjcYoCT4ZvxnDN6F1topM1WU3DQD2us0kxWD9VPY2Lv8xwfEwwVVqs2wwjoFs
xZc2cBx/wEvIqR0otupcUBUhFhVcc3uM5F6x21mx6VQLc/BpcxPtntd8MaCCoKbfKah6p+tmdJuj
/2KT3Qikf1/Gw5hz5x2Ksj8sv+U/x1OjVqp4ZV0BNlBI7Szob8sLI93mJIF6SJ/2gseyF1qK5pO9
eSnRhZWDmLtzqlFVFYIRBZY1M/I/BwfQuARZxLwzp7b1S81N5mqQo0crb+5DCrwuTKpOKkABC2gA
w6vOdI57ryCXSHxBytTQmJKAiTxtfcZxgStRPmbBguKnotWIFKBlKKppb8NM9QJt8VtErqgoDihq
mcyU/ytbcqIG9oiovSFExwX06+axsbwKLcNsofO115bj1FU4JxTv3xEb79UIcohHUr8guaHraEZc
Mz2hGrZLzMWMFBzOucZbP4nDkqfpwyhHFbPdpArFhAYGQRwylUZ0Qi4RaTD7WYhnnaZgf9L9n9mK
aftmMWS/JIkc+dp9FkU5W1O1YezmMAiAefld3SUe6PeQgphoblD4CUjjg9RwbDpy3FCh61jNawbi
5dS5Ag6OyJSIFxtuhVS030RNFbTqEBYpe3cujbvyDaboxQZ24nVUYjtSaEBWFH29W5y/NJ3T0y21
N3UOZfrhOf17B93dzHhIIssSiLWRgzgYHHDSo+rWuhalHHfNxLk2nvnjbsgKFbt2kERrJm47o2G4
Y5mlNgFLfc9LVUh9EFtXa8qBSQCLco2AaInQdNu9gqFpj6xpNRmU79pf320fLLrenfRpRiQT9/LN
E1Y89zCnVe5vLAmSkJpXrR89q/+e5UnUq1vXwv5QKgZOL7WqM4OKGfqcGkJDU/MLZsUxoeb+a0/9
dfa8ssVvBNnoD0oioE10Tg2Dj26q+xLTXCJ+9nwZmSlIbjhwwvQ46zyzGgCukzQ4o7CY654vMPIR
GjIQPd8cpkQ7Xu4iyHSEVpnMaxqmOFPdRMoMvzYk4Z+huL2+SY7UQgNVxtSfmSlbfDGDa0hjjeyd
tqrGNyv9jDiM1W2UBDvOnDCcTXePBwLkGH1zhVSc5gcdh2cLOMHuLq7/8SwPOigfdDIfQZi2LESQ
4pxgyp6+m09EKnMRnq0eFHw3GGJc5AeTbdBQC1aKeBQ+8tKGrZ7FIHEhIsLxD3ZXaNZ2P9q6X5za
eJ3TjJPnF7Vv0chNaFqRuwkE2TQ0GvLFn1qBDnvXf80VtnkLx+rwf/BOZuaxk5ixl17FIKdzjptB
8sfQIgKPs2mBFipVNOOBALqPwx76dsWrCN0AtwBNjRrJdTuZBTf0WbvWSC5/BbpbossbbYUECvZo
uz54SgXSvSdmMcGgA2jPNwi1pxCkXnuoSI8XsJOzhF8cAU3vcEVekVijBS0EY+RgOTedjKz3yzdP
OssMAuDCm9vI+5QWSrPu6ctT4ugsAbpe98fNRpyLT/mT4vpkZWu+0j6AS/+UuSiZVh/ofuqIXnOy
y6u7Xp1d1VHg9YLRTWcIJeKpI9H+SFHKNcRJ7YRgk8TcbSsHCXfiIlwb8KxNoYFolKm0bjLLF3PQ
5LUyODPRKO05ni8+oyOBrlTcRnTAQqqIpREeaQkeSYUS2Iu1fLOhORmJ8HfuHGbsRHHF9VY/7IjL
0CFAPqAOeE4NVcMu/mNNzQ1WWlcFNDZKKZSb7dLbvSDcDXMnLinULi5Ec2KF2DHYEr531eH4W9Rz
cfQaLLUGOVIZHYn0R9dYBERwQS86OiLzIQtT705DvGknnnZps41/E1WgL7zkhMj+CHH+4IUfx5OT
tTUP/Z4PpUR7rcPjR53FODi3cm++PLPXI4oX5MqcChrDPwKMFnaeryn2+vc9Whovarix8NxWn4SY
viJFtUf5nf639N+D3kIvOZNZDapQefOyg+Qy9bntRGW25ofEqR9yXlWbmwbO6B51qy9MUgcZci7f
6mbgxUvUbprTzo+ujHV9Fq8TiBGAqxPBfRJNlRs97S44ZJCTxU2eJtGgVg3MGL6MR0ogxZ/PycPd
KqsJLsZxVrCXaU+0N1tRxCS+NQMaNxONI1OKfo3Uxqtn+hq0zM6o0fIDKxsM7VWVDVKptFgLNN/7
9+PzyRHQDHt6yHB3qSs7S0+O21XURRwiy5upso1afJhUMKv2cBNcrOdBTVfTFi8oMkbawuXwPQpr
OCPR3MP9RM6xQByZ2gYJw8NpYqa0onBW+D4TtWTZDQvczP6jrWf9D0bS5ZO6NKgDMdgY/AuP1zM6
K2qUFYvwfJIU+4ktTOGAqfxzZGvLetOCDQRWaRmujj43xuNXLYezo9PVD3n0ftDMgxU3Yh8JJBKB
UJfj7zrcsqxlEWsOAufHzf8zM1AGbc2LvmEgEKrrkV8GKvA7UZ2zDSJhi5stwZxgln46veUmq82u
FIfvXmxhmAdYjN8tXQMPWtwWxYjIZ/ZMd2dZemWRvzCKeAuIZs3mgJuvYmSEAcQxQLvHOxGN66UM
ObOlCYOrT+DuYhh2zSLH8Oh60jvW831LG/CNrboTa3yrLYRzdBarqnBiYY+tX6kcefKnPKdBjZVo
xTEYSOoA/nyQq3wY2+wWMk+e/OwVfmk9Pm/QKtXbSvsHQCVJvfq6Qa2lQr2zG0J9Re9UuDimRcxJ
bWgOmkOQXVSjQmoGHZ5os3pJpb6FzCICPwWnn+CeuB4vFcWuQzpgBu2oaXOv8l7yZ6ymi8Tebcg4
cU7QoCbHqUFabt/pKSSARNwGU4/dQIfEq25gNbKKXEp83xfRYxTf1g++MeAxavmR4yl473FPpeZU
cfbiK4yOKnFBmocJ9QErpxltEhAzgmg7tWG93hWtTeu6/QUCrHhxwaodWZ5ek0ho+v0Qli0IHC78
Z6autM2vDbv+rrhqcRDxvxqzaUA99MKZnp/F/jENbUoBmS/TtUPMu+ygUpsqyJ/QguJTOOuMSbZT
qX1R1X/RjFcfN9ywt0jSafoZR/cV/gL3wfmd0eHli+duqh4sSJxVAo2OzxaF5gXyfylwHy9g16TR
B6c+gLd3QExaeoMxkUx3+4T6UdjvLlLUBHmzpyhBjWzQCeDa+OQeEAfJLxmrH7W592jQw+r08x0e
CZdr+DpdusWJJ/3XUka89kr5Q0bTiCypD1DIX3xm1WA3L+Dla9abzRyWbfplgi035CkZBiNN5naJ
MlkXOnMblhK7vrB5TeuLmUBv2h04jW7qr/UbAmJGX0zH0xKyux7kHCBQWQhzbiiXpLA5POimOmKr
eAhacsMj1SozKwC+mIKZ9s8l9HaPbW2iEsjio7dRq9wL2oHIBQVD/hq3vvsxXVjKvnPzIF9t6f2Y
twauKcHMXjkEkbkzBj3cY1pz0M3oCa5aWXYhPDv+2jZVwbR2rPqECF+9JN+4Xx4oF+Fj+08hiWs6
YHeZZH6F2d9lqu4eHsQKx82Ck8cH8tNuE9hSdt8KgDSMfjVPyf/emULlDg7MglgEGn2jOeR5+Uob
XgQdxe4vm1ZKmdtxsGnQN7e2TJa5tPJVM5efuuUu6WUDqPPE5/4V2JFidVI6+J69V/+uYpnybUTO
xdVftyem1isqtp3kB1tSKgxdgujZPZbV9uU8/TmPYhuU+nQUJ9mHPEfcWN7XlyFOjI3dvvXUWVed
quxurTR3pXe0BfZ1MMSaObpjNFYs3wUvh8GMvpK4pDqDCh9jRfVLJ2s+YK/JpBuWbLBjOgrwawRg
Bu3tdmvqXeredQHcUzuNdeuwIu/srCyPxC+4feXS/0gnGCnAqekIySI7qxOKbZTNiqCbK0a7gwLs
k+7PWwK0plG+rIrB4Ej3eg7q31Paf2pmbTwYEvEC/V9+ABqVZFCpIRfK3ot9M4fM9uaxbfN0peiL
+xxIiwXix/8TheDM1+K5k9KshM7U7rjXVAvb3vlxSuYCghWiTNPYmE75T+E6q9PesKWGyOEikxie
tRH/pADx5176ZyYiIF6vTN3ZCHYMEstCIjvaHPe4OvsDIUZEG5YRXrMwkUla0oWisoJ4WkrgYmiw
4iXhcn3CsGgISPFLK9zt1Dxr+Cl3GEHDydJAP/sViEN7GmVTr1PX+3cpeBRp0IqkeE3LwMe8jxE5
igF6zhW/Ymz9KZzm3PS8OnWRD0NFyfJVa09J4/6x1jHd5oEZ3N2wB/blKERyS60hmVhu/xilyoyu
UPicG/b5f1Q2bFthI/wLooL+4fsqnCgW8YCM622M1Qr1f1xnwBeuZGTylXgqXeLLdIsVOM+tfTC0
TCkV1JIGZOVmCN5Ces1Z3qOxIp5ZjOzZD1Fig2k0MXrrs6KK607DXmYfeywTmMhUcoaao4IL3+47
MwZbdfRX3LdlVqeM7SmtckpqKUNBNDbOut1GqMrr1s4Og+lNJBDJ7guO24dT4PWT5G7qA2DytTib
Syp1CKbnyKtrCTvehUYyCBcqzG0QYCA+YhcqjW7/e0QihOVn9bOFFyCcLmrCeCXc9wGZrBM9qWk5
ymDXDXIE3jG3SzxqZlsVnPyMrSb+obLROpW7JKB3cCQI7Ou9Uhnysl8D6o2Bd8efgVwffhESFg59
MkC5kmK4yPA73f25u1dqZRlcCE1f/KnwueHQ2UPi1JaOyBPLU8LnwONnImy199YQMBHLOGY9BHrT
9ZaTYacgR2NVwN/xvm1gr7Hfl1q8fOojnQZfW808ehXXhdklfXRDU+hPPr0y3CoQTE64NpSX9f5h
9KD2G3os+URtVeqedP/r4krGsza09rMSXM2/ZBOA1L7mPFFkPjKHLiuVfzADiDaqFkOo6QFbpiqP
mpL5vjPJP/QUTxoJAiMsUr6hJ1xVeZpUfAXgzc/lVhfcssVu7LixwC6KdaKZOkioyCgX7NWpuT+U
Fn8cPrV9FdSCdWFXbzh3vXCsO/k9/6XKDnLd3iM3xdLyFTxX0U/03YS+/HZm1KQ+y4tyJodX2Uv0
TIvS4/HXGmmVhNca6JkG98aCP11RZRIGUWLJsNU2XlGK+p9IOjUyfuDUKm9B+wxYjx5OJoiK4iEp
Ep9v+OiNU4pq/0yFtjklaQnJDw5MKh2dU5KurtaXNmF0Pgl3kxE0h65LxR0OvyOQYPi7zWA4LsbB
ZzFCu4OmxVckAwaIoNNrLoRRqzPmebAwyw5D3ZsZN3A4va1GQolNvaw5CgqkFbhr+n9cVAvX8x9/
7hnh7aUsmzZ/cQmFlcYAyFgKmRDcZquuVxFJJ0SAfySJ7VhmCgUrrYfHATV7UGvNXQbAWv2ipmny
PZ74FPpFSEuwcBxMR79asN4H8bUhKZnZ0nqO9DGS8mt3UCmVLNcyv9hU8wTEk+X3FM/SzkCbFt01
RGdF+px30kjIAEd9UhTTz9BxlwkrmVvLeNyMmwbMxMIGw8hymvnW6IFpc0jsfnv5mYM+heDo52dx
vfv9g2NYzLWv/ikox8mY3YCTS7DWVRAm1HRwHv3PA9zaWiuEh3ThAJJMkcEbUj/APYXaVdtEALHC
iwcSr1JZAOWGnxHeEdgrmCmFDpXCNiG2zT2vaR9v4lZF05JC9+oBGwKMl3rDL/LSJH5AKPBBur0+
3I+EjiT1ESAfdAo2XFQe9Uq4rpu7kh5oWTvhm3vYPd4W5973V98WH1TRKBvLKloti5L20Z/rIGmc
S+UdJ/ozaTnwCTP8GTDRdhk8CtjT/z9JUf3BOLUrJ+pTfJ0AiDyCyvYfeIw+LTearCM84q+/U7i1
9PoTDI8ax7Gb+Isz3EX3v8JV2rlz34zTaK7wanOyFfyn/5i5Un8jnSfanTQsvNA2dtzINKRcA2FS
KehLtJoAI08il3ziodZLeNoWjVdygoweslgwzVOyvJSkazpBE6iArHkUdT6I+WZTr+MDiNV/1sQH
yJ0BfgeGP9aDWsft9qr6QlFLMFmhjvR3DP6d2VmuZldBQ7DPY/GuAnim1MBu2hiyVoHeRAOlDHBM
2+mxcxOLuq3Ubh7pfUPeAeG/f9IAJWz+JLcYlQ/ujcINHrlgum+UbN+83zF3oJHN4+IKRVhkc2UA
LQ8nx1GzGIOhleTYA9rrrqq3PCEskZSmegQRHxqtenxlCVQIIK+5HpgrLPajVddyktmeVPHOUbdE
KL7wbb1PJQNr1xiMeifTjI0c0UEvMg9rLVTzmFlOlqSd9941Yy1/u6iSvP4pMLeLAchKpfkvQKUU
jY5JG3z/MekcjrJVMutH6MdgEiCZ9m7rIidawvttJ01b0b5ZEqT39Q8eByIMRauaU7da8MQFF2Gr
sFY0FqrsAqFYK4+SsWSCKbqCQ0EmZtBTCq4nxrl3hZNBGv8uiDUS8wn2831cbMAQdJGbjPX5CML6
IitW0RPuZfTA3FszjDpNSXlPmB574y5pEC+I+gYgMjWktzYulK+QqqlCc5nwUnrShOz6vl2Sk4i0
q7vNjbgdQkxRyHK6DgErjZ5BLHu+EQdlaVqbw8Mg3dbc9BgJhIRRUUrPIPSRuXdwYgbeNMDwjS0+
+hb8hleeVSd9pQHNXxooZE70VqTSCw3Mp0a4t1wtYZIzY9l5xWTKc/rBNXnCt3/rPgtCsGUNuGDd
yjBBIvpgCb79zU3Bv/AjkYKZBoucvk8BnRUW3jnNIH2TMZgQiiqP1R7TbLUlRt3z/eSxsmmKGhY5
JOgn5Ozt4Lwy0Lc2ackOSIUbu2ZDRnOtzaS3/Kpf2PGW0ufDYTzUVr7K0ffeF4Icx2i+4z/s0ufr
tyY5Dp/XAGeWBt7rz/03Gdxllq3Jq0nu84K1+ax42/i95yf8eKLrsUyp4gplGWsAzmQtyJsxbS0d
gDUoGjiq5AX0fGY5tGI6U81BkSuOecDLKX5PrRBJSQ6qsOq+IksYUPpocwuAlPmrcYechqQeQcyO
GHgY04P8hrz9n9sDz16is3TeX/utfloRp61gR/vyirxpUtgOp5VALbBR2VnGzqC//D33Sw1ZGy+j
HuMReulvuQ8Rjen7G4Wjc00KJd0CShUP+f3sHqyQpMhaxbdY7ZC96aB1h8I497DzxydphlxBsmsk
pyYWqVkjxN8q4xExTif8Q9aMUgWZByGoXEvvxFhHfBNqD7K0MYWmMxQkcdHKOhIE5qFlRYRgjeuQ
pViPCLggEfle9KCkNZQLPhAoc3tsJkHB5k9Q7LB3W9EttUA4gabH2xt0Ubfy28WYMLGTMCsgpsrj
0DgehJZaVDwFwx3IvK4OAM5iHeRqyjLTDnwmBGw+rQR4sNE/LBY4sU4y7suC9Jx44i5VohUsXxNJ
A1XQoKD6cuQfVhphBd6PEEA3M/BEMZHp/2kKAgORBlNrSBlNhKE+o5/XMHC5mQu8nLNeAm5uHfWw
xtGQJABCqjKbQD27KwcT5etWZDW52qqqjGxRgNbSRe70cVB2gDJQFcMk2vMMPjNtrpBFfeSx6C73
w3mXMCkx0n24Ol66dx9FYGJEvJc85U4Mgliuwanh69AdUWd4MM2Fhd5YUrNeyCOxibbNXdHJU8xo
hti/RoXS2O9BaiO1XyRWz3WhZ7tCrqr7ryIGTRP6K4tJvSQ3lKOARr8gW2Ci978XUiZQ5FXyvYbC
bxfwB/DnTzSqT323iW29dWOS4969NDCHzhhj1MuGK36CJwcAnihuA0uhxMHo2iAEua3jsQphxbhH
xyL8bANtvWduLZiJGq6PcYxgpuI7nTiGF8c8puQ2pCmsuarBhgyOrGFSh8pU98QUbZIW8K7dos9X
ksmqKPNRx5T+nUa6ON5GOBIAyp9UIC4rfgm5Md5UolviM0JaeGWPe0ByhE8vJ/pwY64qnzfB9ei3
LJwJXK12gw6BVJj7u+hzAVfkjEBnqvOgXNUaSNoKACitikyPjWu+JFOKHP0ytplKOyoJ35Le77v0
2yaCdsooMXyMGqEnw6s6dvdASGQAhXzMDKU3VPtanxgbnfPGo6yGDdFkcQ7eTpsQBfprmh5Ry9MA
YSb0eGfpKiAAgamoACJC4VE5HaXTaevX/aUbH0esArwWC9kpV4f+EKFXdpIQv353hOVR0KQjgdub
JK0lml3eHmO3MBi1XS0I62PQNefkCI4HuOfMhBO7IA1NkBZ4cP/htmdyyI4VIKABqVJLThmlxxeU
lF0gToNDpz1kRRx4EGtOnqtWA6MGiTIAbik6NF8QlowYxfUGKdl4L+9TMag7jjh0Zoo0/QqR8i5M
Q0KOx1xLrWBqpMRwo491oPOqs2Jb9/9vpFKR/+wdWSPVjzfi+3+G7aJOVHiw6j5PfDP0s41V1jIV
ZxWtxH2ZVPRcDnfCLvJvg0ITa1kNt4OWggzqh5yQZfrEh/UzAUSWYlLe52XbvLI2oFSXjWrCQfLg
V7PI5j11CIououE9CsR4p7y8c3qyaQCaX2F/NBF8FwtJ7XCiaBCtMuxC9mSKwIqD8iWrT6AFtdSn
RmyFibSgNE0MJzokQMwDHmubtsP6WJ2HiATo4SIo0OmD294Db0zG0PWx3aZLk0FadnDI8xHqBEDY
W4/t47vbOM1APji/colV05vhzrgXmkAzBcYcDefnB0/eVOf4x2QXizVLKNmgg0hab225pr98Ved2
Bo2jloLG4GNz4ncPKNNybg82H1FBGSWBrkmxhSoZEAFARJVAe8yA8bdBPNDEwPNcaItOjc1nq8i8
lNXMoSDpG4WDvK+Ba+ZE/EUpreHqNJebwcbJQgZ8JxvJ3D8jxVR7YktsEvy5oppSad9h6hmp856w
HY7VzJctsbMASPZYGnuIlQgiel+kl1rty68uAqFWRPSANaxfSIvFHI1shYwjrN6mj5FuPQhTQgaF
5mjfzA8thkiWS5HKb8JDTg41/XFD2psVR0mVx6uVD85BceDw86nhX3uhx2WmgPPfHiTexHntEFwG
xqmE2UsVbOKHLofuyr+L7wdbWgl+FhMjVPZYc3jo2vUZLIuj7HFT0QmzZR8RYpMbsn8Uic1AVBYO
YoxeGO7XI+jgWeUcK77oXxRgq9P5h5SXCkmRUdTM0DTuHxjzHag43a8Th2vLyvfyOCxug4MnI4mQ
jesBPzEuRchnqsAEIVpKOdMkzC6xlgwjhY8sncf5nFsn1UEy6LNmu+bKeWFS2XwX3Ag6TKpOwFSo
F3OoN4G4Q0K0WnV0NmM57nvqqs0ZFwoHbHkBZqsAfNMylbQ6+6p0aapYj30cWPRYDQBq6ZA3JqC+
s+6afbXmxDnDRDiwk7fgFVF+4ylHZx6n1DQ0o+JLneK7FlM/CNwIVLJcfdygLBF0zHbeHxBjmN6/
uxfaY2fJyfv1LOqMaD9JRJi+9B7ursa7G+6ochKVHgaCpGF7Islwdq981kLnc5vozBJGASPqALIK
0EG0b4PY4bQkzagiV9bmqjmEK5M2RZP06PNgLhyBxUxfbOvglTkusMMtleiU58ApjWsntlbFUVwN
7E3SijkremE5vuclOx/K2Nk3ob6P3fFFftr8t5Lzdn6NYIz3DsveP/iG+rk2hc1bTdCerwPdgnFg
tfRmDdffls0ILz655BnQdJlda1Bf8vfjECzdirzfDc5l1pFWzHL0mfnYFv6Nhct45P44k+JteHj7
NhJru/z+RXLjMdkuQPC+A29tmITqH3D9BHZCAQMX0OYJfNp+zZhR2Matte5TlW/Q5TzyQ8ZUbIdg
u83aYud+KIviJHRe/ZQYr/RYGU+a7Fo8qXIY7TP8kfXcuIjPYAAb2Jhi4IRVwb6j6eBOvgJzPZjk
LrRJc+WPTHrAUF6ge8ajqInQ2OHvgHuV4esjqBlaN7IawhOhxpZwyPef4Ua4TxMfGjcnd+psgbwB
qbhSZBIWi/A3W5I8ftNhd/wxY3fY2TVF4Cy2N1l1x5PTAIO5JRF1TorS4vxYibtaPSi7SfZGvpSm
8rDYW0HrrEy2DKC9lbcaYZDigUmmds+HMlw6Q3WA/UqHibZ/13SfXealEHmptWV7lgBFGUvVEiN9
lp1Ie5nNoqKZU51KxP7yyvr9lMSI/vp3l6ZcYyzhi+aqjC6jCmWrsRvPxNyF+9cmch2W/JuSdylU
6Ua2y0mbR44Z9u0Pp53f+RRaA6qe179w72yTRjoIk4OKJdbjPvgqCjpCSJySnh7Tk54TvkLdGrJQ
ywwxKe1XakoLNBx0ugK2GsO+zbC1+yIq9SXCxBCPnTfYw8/S1I0yRpkuSaOvZqMqniucWzzVi2RS
zxnW7fRoT7tvhVZDJIFfxXsw+YP3Yc93iOZTTES5WlzWBFW8AHVk2dE4jD2cNOaa0hgbcwgiXDpU
OqFwxiUaVoweikWVIwh3KwbsHuFmZT3Yie4TavICbiIO9wXhYqQz115y3p0NHp4NIvKcCvk6zfNR
9lytvJgreRiVFc+e2sqAHR3AiPNzEMRYg/DyuG4zBSVzc7S/lGtI6heVb/8ViISgKJt8lx2Z+/xV
phEQdnQkvlc5vWv4LTJlL+8thI9olzblRYfseECG4MCSYqZ4RVJzIB0WrtMgslhhrXnFAeGWfMfA
mHsZTuSmXAXLFI09F0qdUOOJU9gXN0jITcJtkI2G7urXkDxP6XL1YyC6QIG1KQmbOBfROS/jnBjS
W5MVVmhzJCW+3ZfZmExu4GqEQCL5lcxgqd4fRo14nTkFny8Mz2DqpMu3p3VZTFtDIiW2qKao4eHc
baSXiHGlEe4Egy5WJPP1x5AMfoDv8wH0O0ZQCtIAo1DWdCFbRMwyae8cMKi5fpwCpGNoTJKbS/5j
+37tkq1VNjYJkTumQIBQ2XntY6xIchw2TsPOdrL0/SYNDHeANumx2ge28h/PvRI9FMIHveN887mq
DfZqEORhGiqpU7Xkws2swaUXdTb6Wd6l/s3JOSQR3KzHJ/YzVsFftjn+1E92bA8nmX7+gLfELE4f
kJlLtOta2ChVNJMz5c13LEuOOh+z2MsSUTQ1L7M77jypgfFSfofiKLhrABjcV7h6C6aAR2sWVB3H
M0TTmFF2BrHMdJKlIFrGlOyezsddnBdociTlUm3Aey043e/oNGxgmxMvexCSDeNY23MgbNfqj0Qw
FUuBZXsR7+A9D/omw0rTxDbcQO1D+EQ/p6iCiKJ/2OhSLdZxKkeJspY40YtC49E2hpphxCNYlF5w
HUSae5Qove8yNSeO21l3e0bZBzTOTHAv78vVUBhl3TSjQAPVJtU/7vLlWkDHnH5v4FYwxLg615G4
oLVCebUVU1zG6uZYw6w8fFX7/YGFDehQKO/EihfiZtn/dw58OEomYNvbVjTr3R0i5mu66e0kHOgY
mNRwHlaUIdmdnLOJoiOrRVk+HNu3GrXUT6eK4emuMruGuWtQshNkG+NWHkZbX3vONhzhY4A7veQu
xsaD1OgphD8q7oho7F8sqPt3NbbKU8aLS0RvYseu8I2rbWccLtDL3mIl2jM3iOVce4hCmqfmVHk4
1Z7o9IdBqbvVd7MQOFF7hqkkGpi+ID1FbnEFjktQ30i6hjUi04vyfUOlUJIZ92VKb/wB8Ue6Q1oH
hr/23cWbLwOgoHlAmAgzaMOOFWiN2nbhlS+gtrTPB1IaQJck0QPN/CcMRRaaPjsfc6CxJZW5D5FB
U2SL3Zhi1yvdJZhhoF7Hf+y9HxLpGNTIzqldLqEKjWVhfsT8ZYy9C+bnFeiwg860p2r7rFnfRU1i
1lDlsw0N0yTaaVuGdJNsMclzZYbYIx9VqEWGgGtWOj8FKc4VZdwE8aqcLSiAOJhWmI2wFbEbdji5
9HJEkKrOJ2PACnllrC7m7IRCjO+np2wuzI7Av8dGjuSJuIAUp9bUumpMB6YGddzZ8RbAXv4p3dSP
1/b1ORuGiRjUi0dnUh4K81w0NepcK7KPHPpO2mNUm5kjEGQcNr7Kbk751YHi4IkgSddTh0zFztsg
ZFtPyes6nrhGc7lE0p4cB8pY2SpJBAiFjcQKK0ALly2qV+hxvSk5QDXfNgMvdYHvUqHIxFuKFsmF
TydkBNvCKOFGZQ5jkKtJLjghbdmcOZnlqHguxrv+KcDTQF08/z3Yyrou21HnrIDpnKLmlas0SYIW
LjoWoSrIpcwZsxAiv77E8itzUoyGP5gNs7YkjKeFUAU8w21fpD/yjrc2fKiubsM9J18q5dANYqZF
GxSiGdk8F2pt5kGj/IrjBTsog0irrfkLNeYbKw3tn62j5kRPr0jMJDc+24BzAjKA+xEH/OVr4ZfU
/MdXsaxV3Bwb0MsGu7eT9sc9hYidJsHDFQbr0x24w3IVUGCcM/SiZFcRHgvHJK/Dszc2tpZmLkdz
VWFgLW1H3US9fO1HRxxXW/eOy2eLluNcda+Lw+qvs9XyA3ebTh0gMFHKw6+Nu+hi+ewj6FBDd/10
8h/0fdtk9ofDXKebwg7yISthaq6/Mnc6qRfxg+ZpzPCrbIlxvOkbcDFGYdQjHO5s3Tq2OfWi4fpY
fOVcRNvIB2YiA9V8VKGCBnND37PIrxz3HE/gkuZvvF1npODFrVg55+G6p1oSYZfFQws88q+IDiTO
grhoxxQsLAGL1/B0j29UWx5wvckIb3BC+HQJP14/IMuk92G9VxOSUKsQjO4qOoCRXcdQ9lZgaJC4
I8+W8mRR8HciLc5F7T3hGx72AfhStcUPrCYkl8DEUTynjoC+nxcyRjxd3wCX7obqi8ocs8cB7NcY
wKkVcY3p+kWpJ/+Qs1GzgU+2gSd/l3Gm61IAxYtd9t+qMXy8V9+JDVh+51UEDwqz8tu3Rq7QjrDo
nk7tAhLeIu1Y9xTYMsYaVezv1co3sSbUJ8QOZbIPQjqxxYvBZitHK6Hpo3M6Up28wUedR68UD1PJ
WYmDCQkiN7ZXNrr4PIg26IBtn/WvOwiH9bgLvgLadpQdr5RUZBir1Gr6bPcic5nHdzWmwyLFxhIY
x7MnWT9NYrQ0HGEIHSeIrwqNYcvsHoBvQhhMh27JqsZ1ouJkOF04HIuuZvYmwyOAzs/CoEYIgd1S
gCn2WysZnFqm5smeOdq0+HoxCb1jHkaKhr5nyuN/gZPX2DC0IhlAOrutGrO+F/CieB4gtcz60K7Q
OUDs082HyPhp6KT2y9tICWd8vu2N6Frrn4iYwFG21Epbj2dt8DX2QT4dx1mUwPrsDVNfr/UlPKmb
Io3Kv8FuzDc7tGKCvrq8pbV2XJZs4uMhn4n9oOLwkilT0OdDFDVDD67SLviFg/Wsbj71KaqjyGY1
tbJ9Ep+QQUS0Dt138kDxnwyqLZ9VOkGls5UDQuftpOU6TXNMH1z7Hb1Q1CD57Y7ECqnFe1qGHRp0
NdOEGNC0BdqMI3kkSMzJ2qsk9Q+0LtHMgNg5FcGHF6r8zpxOUBj8+a2yeXX3uX50Owl4E9vjVGRs
sH8sT57vTei4owUo+3Xaf3NHj0YtAKst4Mnf4XqmJRDVo4xcr/a3VMk44FgISJBfGYfXffn3P7cs
djMoj1fG3L2SASnRmpzo/mMayUb32rZ35QFs02vfO7OZU7m1Et0J0y7EMizX3nrFjyCBa9t/lShz
OOlgyxYQQ1Hu2hvSEHEr+zJCRXPq47aXSp91WdfybbCtl1qpixOwaU2KRdE6MwEO8kPAgw3SHkUZ
I1Yux662kDvBMHLOjsv1YIlccX9UujGlKsnyppXHDySG6wVcOXrML73sZAwsvFPhWacrJagShDYI
KNMLaH4RRTomV2elxu02tx02z0B+1SF+OC+hPGaGqv9WytCPX8Kvn9ghFHXtFYlQBxp+7ZIVBaOX
7NszmY13je3bCd06U6uSZeLR2FTRx9FqVOGTdajnxqO3pMoJ/IhsKWTMczIODHb3vSEPQeLiL8Zw
O4lrKtlEdLS5uhqxFfBYZohyVHHzSHYqd8/LHJF1qxlCKsShvdZPqFtMN9HqqYkjWB92I9UPUvoW
jWv0+UA9LOQXQUaOXmewnGzdVkerCZc1h1btfkpKS8gGzoFPxEWNVGbXYFWRfHVOHKH0kc96DSjT
XXNAF/angz4fwidoLk/b+Udtnkh4lji6txqhIBxEF1iL7yEoTyVfZ6nFqMZ0jkmO+DR4iL5f6fAd
3p1pefySePQJqZ0JHNAq7Nf5e4rDjowTtQ1kgZsFrGdpcgD0182WaZenFUJePn+7t8E5XWhpisNj
DKoX+LjIXD2QV1zUs1EpytkSpQX/24eozBQWVE1avLVRFkQBHd7Awe7Q7SJVlfT2KlPQ6ryIooxC
AyUkKoMfNleGcU4LUHw1BjATp0xzTZJcwddaHJyudOv+5KC7cKEwGtrLw05XfSIfXBK0P+jdpee2
8K2x5Ep3RWz5s7EABYPdBISswLEjgIGvmQ92mRZWspVHFfWrUFIIPhk+8NtOUtpbTT87DOSKHbmk
x4clrgmn/gii4zy5OlvKkS8PtzdN8ycHBGY13RuENdu/RbAmFNF8oUF+1pZEbWS4pHt0sgTSdSuN
ZlTCXItHWWWoOyvoY9tz45vO76+0iOUDxAotvXYCifmidoSF/SUxMqge6YIX3pKlmNCp0n1zPR4+
aSbOb8IT3tOLAbsQFgXzsLG/VwKG3JwJ/ps0c60AToQ0GKh/0cavw9mXw+VKN/cqvvC4MBwHYTSH
n3+6P71xMSo2gfCfHWSUBuSHw87P7ULCYjVewH2U8v/gA9OzRthOGWJsoD1fLlxn/Li6arjbmXsp
nb43TBxhkGhurdxag20VXveaoMM6HW7X7SmR50BVIusonwK1L7ZPKUa0dV8Y/a1632DFRyJl9ZSB
b3Iev8QOO7yuSTt7nKWv1cWWjSS0SnbijQJadnO3Fjvc8aGAddDVosqgC32aoHJgQlRTjHA+IjGk
q5MdHBiLbIPp4rmpMg6LBpjbkVut8pxFb19aRDkC9DdGx+4mQf6HZSWwuqdS0/ojj/EbGraB1krP
Vm3WtnFF36zoFkRS36E8/wo/IdYDoYDc4XM4TlqhFRDqOq0YyS2Rxvo3J2OypuHfcdwJbubP+zT3
IhFPBxpGY3ksDXn0eK4LNZRZ5IdWkp7+RS+zpr2p0e8f2S9qgaeBHAf+2yjA0wuUj5i1Hk6BZwJt
vb8AFhnTy4oTy8wOrHHbUOpV1cXWpDw50RoSKXqM9qexdjdaAEWHrF+kTyvXGIx7hYKTjkym7z5c
A5byGzEltnFKjA09Rpzo8kFxtgoDtU/O8OSRu1HP29zfGUnuQaD2IqYT7X3MzuTOgBhfE10U3xyJ
sVjxdIK4WuoHtNXRmBAyNGvWYpCu3PCewmTh9hk8GQ5Za6CZD6g+oQm53MBZZbbHLX6U2Fjoatxq
5TSzW92Fgt5KeQgCxEiEZvipqqFS5CKqL3JdwUCmYInlpBpF7hGwbCyjI9AGQfa6tfKQOv4xElQQ
5lWDz5dimORd4qyxfBiZQZcVnFlgq4se50FnaWaRre+KO/IHzdJiGWJLSkEYOKJHWJSq9xK8gB7D
zdH9khMXZPQscTq7fk5XCSXkvDV0fpu2pZ0l4Y4ClWgMD1JMw6FrquxKUOO8/NV4lq+4jUffRi1o
mHx0t9ujPG/fDnGLfvyIUl/4InbIpYrb6EHhkWMb+eG61BL8bOc2drp1l6jwp71ti6wbCG4Hpi5z
WyEY6ARXey/bfU6brKGBlAIjSmhGGb+QfVaPSLiNE3cfWKC3zDpJryRasQe/FVRVEkhOyMf6mM6P
aQVMnskMhQ0YQXkbaqpjVIylpjHYYxGDOEPGAkbwR1xe7vPIcWbNSzs7HuYg+3OMosgQsQdP1eIQ
Mx2hh9hrmpqAYF0M0F42HzX/JnBFN+giw+kAok0yfGW4NLXdtx6H2WYUpgzqLDS+el0mfXEy5mlu
9dLDriN1MLjjmKt1td/Y8oWjFG4PmMrkYMiknPEB8CatfvXhcqyihXBMKlaHzT/Ea5g+OcKK6klM
gxp7sAb2PssvaPni1ABJU9xYXiA0cavQjF2J1hAZ+vcLnh7j4YOj4CR37a8N5wn/eDE1gNrVzATj
zvPV8dcH3QGyM1mo927bMAWXwxF5Sf7b5yDBGusYkxXRNnO7M7ou/VE7bEH8QhAGvHSwSGcWkbng
xxrxqD/UGZXVT4t66CQxHWpD8rbLJJLSBzYnyq9LNZN23U8F9kmFVpqtmHCnMPXe5xSa9BrYoxnI
s/CLdthtVzfdP7omrZb6l4XnrrBardPSxbDmMHeHRiyZ13Mex8BUPJMV1VvMvar65HAvVdSQstqj
qov2Kun4snyIb19EwkW5u9dVBTCLD5yx7qN7XMZoj5NOrdTqaRebP2hPFhF7hPIX66Vd/ajYY+eH
iWoQUQaRUnTzBnaH1qq9E7eOQOOObl/ZVQ40osgmk259HH0ajq9/SZZNuv080oPzSpB5ajs9lgdL
ErXCWHURZP5F8h2ElyuNXBn6Es1quws8G626gDkBko+21UNt0i4aiPo/gEVOAC7iN7Omgkmd01pU
BEkMk1uNmOekgqIIoMRBF/al3JkftPXYeyDM33Q/3rDyOIa9cpYSx3igXwR/XVnRg7f1mF0ERoNo
zUa/OeejEtHCywa0ng+plZlEWndsOJJT8BqaZrJellZf/fX2MqEo2JnHF3E6ayWST+ox+rMpidde
l2FUEDMvXLAzxgsS+NQUVjljNQBhjH6rfGS9lvOK2aHszn/CIpr9K4peNKPAcCvLbT/dGLpf5u0p
fcOgdWZufk9HWEL0kkNYGfMtVRrIGuDM6uodNSxHX5zA6SjR6cu5nTvVy9WMGNC+tZoj0BPEoDUe
7B12rNQfnYuTOXuJRcpMTlQh9fm3F4r1SFrWIGiwukT4TWxnnejNpwyUxhadbuMBc13oto3J8ccW
M4l/Y2ZQwRmcucFPf0k6B9jG82rr19eX8SaDc/dppI+u0zWTNEDIFA5wd3xPzc1agOL/N6B7sVug
E9tg1VRc3HFXRtI/pQmAtVNMyUgSqHnS5nc0dXJiLXmcTWIU6pauU5vxQv///pgZYU8hwFvwGqH4
GpvUwHAg1HqyhMTUIGOVBFG6DH12S9OPsh/gMBZ8a9BGs0gz0fJAe77VxuQy86bDnIv/8zkp9v3f
c9WjfLrXSMFExUn0aEsHZ2S3qrabPA9kw/O2EurcRyRfWnx52vCmAGHatm51iQ+tQnt1QmJM5qNJ
IKfjUu+XV336g0fP7hRU+U3TN8BZcFWc9b0/avKLjlfOCsaDf+7/6SaGWhviMud0+ShW63Xts3hj
V5xSNPA2koh9egwacyOi/GNY/FgQnSb/6nWaaGvGEqDm8kSqZpXLQJQebhmDm7xsMvAABZNVtAdD
SbbTE0befDCK4SjNZYPx2W1EWYl0zSc0OA5uXaDYPQXg2RqIEXq3Ux/DYZlZg+RwSkzC6sw+Swlf
ureBpdZplzfPWpVaoEW3HcOmt4/aGh9UsAQ8tN39NXwlMzLMP947h3ezCq9aC2TDvSVbGqXc0h9D
L6eYP7xfWeTlSv57rj9UD9Igby1zKqHFICbYcKtUt2YA/sX65r5bsxKCyZbmZEWj7cTk3yZz27pZ
/vmtrFOKDEwNJOmyuDEqNyoxclR+urEJJjm4+5QvgSbOXRCPK2A+dkBymnk6TuaQqG/CfQbIVB62
rDk9Y83pcGpvsVwFOJy8MRIAS94cV3VyibJxrlGCR6XwPDLBweUrsrYDC/WT4g6kImaRoZxLGcXa
J8OkGfof+heNON+Ovhfo1eannn2Bydfxq3n3q1N8y18cWJ/pLEQrxsqYLyy3qjoOtSmXws0Gdlm8
q2NR2R1M/U4mFZbGdIMa9D2gmxAtmPOEnfRupT5gS7cfStstMN+awRLrUuAggEcZyoNsqVWkpGWa
WMheeCeVjQJPPGsUn6YXHDK6lghsBQfPcO3IZU1wgIwAJN/BkWCv9HHSQuyzpLBBtpF3na1XY1tW
qxr6DQs3Q6j6yUdxSG0h0Y2ENaX/vj6Huy6KKU+zMEpsojMvFGK8020/4pVzSha7gDhghyYlDmks
M5HWOKNCwYlSKSCrV7n3XEFBPSePtQsvb3WZmLSkdtWAZnZNUNuIgMgXGWakDcliSvaoP9do8VOn
XZzL7JZzkmXhVe9LvPi8mAiIYO/f8l75VHFSMkQsJvKRw8PDhIv4517SCz50l4yi34qGBXt1W3vA
fr+kCeABFKJ6EYCE2BgiyqbQhLCTCH8VYFwGdtUjmr0cqn8E/9C0EwZsR/AISVJ7Qd9lNRIJ1nN+
dTL/OPjfcZxxu2w2Lem2wxFebwcL4keTuVUMvSscUMOVJmVRKJMjF3s7ym1/gzmgk5uKQzBf3iIE
4WMFkVsrnymjGWWkvdui3veYZxFvnnQSnbXmJlVQGLJ0dsTHYvA9TfDmEO9b2uANWaeHCENvMZ5X
eZMGP/tYl7bQ5Xq9jO7qFtwOlulDr3zc6Z1E0dcYPAXDmWFDvW3b58RwEvQg2THS4YL2+jNlISOF
czKNrsnMediLgOs8cG1iGyArmARuyUHPx0ONn5e4N9ojud+oLPL2AXg/GLsnCPutvsErXL9+DF3A
Q4TyURMY+KermkdEuAZoMkXsIRrFYhgfrT226QEAOzbafWzvBqAW/2jHGo+tdCNDkU7isEPtWZkw
7KNcwx1u2IeiS2giuP3Kv5ANYhthL1G0e95yWKKSmdGeCY3GQ6FWDZt90kH5LKhldFKcThyEHQTt
ex2fCxSBbSp+TMSUpfekmv0nCdtTDIO432hLGw4IPl0vlgT9j9DaXFnwbNIT/EpA1KUu74XzZSX1
aRaNbfpRmH96QrfS7FAvFYvvlnjztPns0IEXRvxXpZDxJkoVcU8nfAlh24tm8PgdXYdRifO7K03d
NxmTEeitTvqBTTzE64YoKKNqbHapMgqlFPUunh+mLJV7MYz06UA10ecjYA8cXBLVfUp02wI4nlZE
bSs05bYdqjqJY87PKPPnNW/VUrtVN697U6rJfORjrdtHCocX/OXsdl5wvl94X5jJktPpzG81NuZO
60BDW+ze/PaH6ZKc39zNvgOF+uykhqK3/A9s991kP++cS7qZyllwo4jIDpErlMCdMrwi6Nqdt09H
MAs4euuKT5abCq/dRLioMBq7xyOBMdagbmKmmsTY8m6PSFYkOHaD8WSNzzvNhoOhwhl+K7Yo+lKQ
w5GQF1QwybB7kHgAZ8oXAh4ig1qRsIhABm/6CcrkCRGfSxwrUtLYG2E6JGTBLLOTqnfkOqj539Iy
LWdQjkaxjOuifhuQseZjvAlTYa7J/2LFdmmphWwxUxMzg+NR5meyA8d++qwc3Sv6tLzVQ1r31gQP
i1frCJI8NRnp5ze2n2/MJpg2GgCqwVhmvXBf8vMn6zEXMpdqxq+O4OqFvn/eNdljZckyivrQPvmJ
Jr+Untb/lEoyZn1WrniLIYMX2jrXjuoJH3wgtq3/NjTV1wusaMBg8tdkc/eGiuDUKkw8fTCfToAs
TxLs9/urKrBjn9JNMd4PHhek+djlr3DS4nFW7hAmrytOqlENRZmHgdQj7ozxYl5VVCoBKRxfgEah
H35NKlICS7TXVt3tqzmu7NJgsnrNnORo0XYmUuWYN+1ThtZnDU/JF78J9SJqhpumCXlpId4sW/We
mcfsj9V6NbtjKQMy81XTyt2CCQyrvndflWG8DSS1jktDHI85GIRlXtaGXeYZMGxgxcd2AhAnRak3
Pw8qbByZ1KKlp7++UhL7WcjGohqMgrIfU35OmfE1aK1wZdo5bowVw+SQVuB/Iad7rw3vxPjXS6s8
QTsYKpq5D3g5yqZOFgBkkkK20pW48GqWw5GnWOf5jMD3Aa+ygYwNerJ9ARjoZ3S/a4X6/elY+ccs
m/kcxLjWFd3gWBiC62Zi/Oy4/+TjsRW2JzWxUd2fW6Jeiqn7RtrSryDVWeCGSabjbmXdO4OMrU0a
UjvOZO72VBhiD0TcOHUYEwv+IHyhKU4fJt8X+xVpPwOYseW/S5MeeFIzpVRW5b2aaOalrKh9OTZM
/sxYQb9h79wgr5GddiPyX7VrZR10ViWx9EN3/XyGDEqPcFJtkEMKvUe2qD47ahK0rpTk8n4IGfrS
nouS1QN9E8TSTLjz1+wWZPKmOPMKCqjNvPS1gahZ8rSxwxqJOtO3eEaerx5Zk2r6lgJf37Kl4ijl
EeLe+oPrUvAQ/CO504vJ2vdoXbI+Rj+ZoSbI0OllG386i3EUTatOQrMGoI2vqgyMZnyRc5ZG36V0
ouuZ//WNrEMSD89mhbrTjjzvEAwZbtw1WKC3gxlHtLgh2rY4vNxt5UEuKFus+OFyzkMo7+ilmlD+
Qr55I4eIsjdhVoUEKibZ54Dyb154AjRC6RHVapaEc8U+N1jnZvZCTAApTT9cJ7LjIiWoPOqUnAZI
oQOJ3lDwwIuYguxFd5tyKR/jCOyRuMAtLmHJjGctQ4DmxQiTQKl/GhyLQMNFkE6sywWGr+j3YrZJ
x+lanxnDhPFzA+wMLBmzoJaVP2EBREN2gOr1w0wkIoJFHQuRxrWiLHBFexlVlc4yjmTK0/4TbsPg
Nlort5XhfPwmLCPgas2pIXHjg2fpYS12IZhu1byJ0Vb6G4k3aAIY3qkEjuYYLzz8BmtVSGvJSLzR
80/sDhr2jfXnHXedWT5PDM9R0W7BvwdRkWtaYp8cqptgEB2WLpBIEc0eXWFTM2wkXl3qNJltGWJz
OzbfGosm7obKyeqeGZpslhVqKrhyVFZCVeN9Psec+OH5YWNmsjk/TcCSIetVh6sabOO06rF3Ug/X
6twZp7YWuaJA9lf+8ciWXGQW/8AhNkveB8v2wKXQL4QyasPnXUscIZfc9K4WfEcLK1hXdF/AUS5h
KODNrWkaE9eNb1Fk5r0iFSTV9lOFZhOs/NNSph/+Pkm3mhJ1bIocVquTuCWeTOHlr7jnQ9CrNwWH
v+V9NJ37PUDuUl5QyZZJLxh7S/SEqM66fsdGqjREsEPU27EPfscn5OucUhNfS2Rj9ofkYw6Pmk3j
P0B1OwHDWMe3ZoPxsKsNZuCZxTLsFVWzdxDhEFUt19cf+vd/hmu+o/cXKC0pgYInpY0Aqxxd1u8s
C2DA++5A5uGTBGBtmBdtF9+Zx/rOyer3FuZPpfwyEcb2rwmlZ9fZQ5IbcfwiTHvl6ukNJcAPx2vQ
ETQvFgAtm83OBnX2jW/71Cyg+5csO2bOlKmv9wJcUpzCLOwWEzflimNsqufHfiQE2FUHtBQKUlnv
7aHslSR+XRyIh+tJO+Zablbrzg1nAtIKbaFs5lCY9vGalWwwBGHGnYwjbMOcEiGvJW6QrNIYsXc4
YPST2JUzE7HqmvNWPuKSiMpkiNWQa3l8iDlErBExdFjaP+pPtLJRk/meoE5bK6Klb6BKHgXwSi3P
u87IRlB19/dRgHVXwUNz/SHvRD/SLOzPNmOm/yExBn1aOqNxhBnzGEJhfp6ByP9hal+F17yUksRd
toYmRhaBZBVsfgvIQ8JrhixT+92K+x17tA3NzWfGUJF2UNUI1FyMCOw4p1cRkc6BdnhBe429xeoi
jkz2QO5K6l0NQtTofl+B0u/fO0j66zTsXv6UHAcFskx3uEFgxj82WfgvneM7sj0mu6dDvrsVSWUO
u5AIYMT/kFWLT7N6TzmlQIOTUkPu/M5zyuNA0kICr1C6UfMMo/ch+PBdBIp+QmQKEBVRH6EPp84R
gYILf0ISouCi+YjeDWr61375yFnCfkAz63VANk6CYvMj2mw41TWVs7aZkxtz8Q9CBsDWU3Hnqin8
SYxijyXW6NuVgr6P8nH+WYZkgsl7zUaZ2Psjj+t+7SbWLVrPZ0NLkOcmLNoeNO58l3BZ6Y/sLch9
jq+tyG53ZDovZq4+neEIGWN76m+MQLVrKT99NV6EImzptEYctkhQN/n54MpQcaj3cp2sy0jCRyZ9
chSVTVUdi7lXY0FklwypqhvsBkx4QKmP1xqhSUMkE8kK5Uu4A6aE7X6R6txqJOHu6+ERNDzhdwLK
1l6gGYNwLvumkIhxRCFuYHb2dwkYTsJE/0kw4vd0QMRd+n3S8iX3ciIYvnml0owCr6Xuq/RpG1v/
enmCDw2xNEPaZ1Aps1m/RY9IzNLNV4+5HamTzIk1IbmcOz/SC5c7waLiyNJi30IAv4hTwhAxoL9n
yOHm4AbSQRAT+SyPDVgqtgTk5JUk1cCXTaprpOhPBjnvQHJ/EnomMFRpE7yQKdhwy4YD3APAHCBC
/po754omTfxCLr771D5iNIx1wrvz+cQ1rqj9YA111JA+GSl5p8Jlsr8i7iIWSh3TOgCypU3exXZS
AWYQpanV+PiihH7EvLmvPN0Eq8fbv9Nw9MFIXXg/B2FbWng67ceL/1RS3ouCmkCALfRPdpr6GKX3
J8x/vuMInzYqsBFizrn/XaOSD/S/VHV4i5KyeLkvs0Q2imRD0gqu+F/rDPeZbJX2/z2IZj7YAVge
O0mkLwhIe6R5SuFgLGcl/wbJY5Vztf2ELu1FOXbKgKAW0zm1MvIN7vNoAsqut1gKy/4ghv4Mci/k
N0tvSqt8LbUMdbLmf8y2Wdw+8oRrRdqfSTI2DenfGgDwh3eVRZ/HlK+sgRBpX5HmnxosyyL/vxjO
SpW4A2TTISY0RXnpplgpGwwJhVPxELPL6wyOS32aU6JDsteZLPJSftk6TOS64yTKWadjIc8c9RVd
r5xNpXRW20gXRd8uR3kMOQhe29/yP9UPXxhgL2lAbhr7ijJExNmhGMYpW8FCgAiEvFfnWV3J+yvg
Okrn7iEs8p5amoVUdsrYDIucHQdV1mjnJmykqklW4XP2AiTJsvtG9Jjf4UpiNZB4UAYSeFaMok1a
SsaV2rjq+zxi3+H/sOUA4WyCZdendiDRfCnHYsQ21GGVAqUVTYNWJOinIinjJ28ROQJI236Rwdt1
8llymSeDob2EfQi63yYYY2hzHIgO7IxerHZgofAWTmCS1Qm23QcjhSVDhasiKPOTlo7WXVzRk4jL
r7Vph/tiOQsLsl6GfQxmwADCkAVg6x3FjphO+uKGB9UEQms4/UwlUFGEYBPNlnlDK/sW+nIqCBkU
2jBo1mzeQ0qV3pQQatqERgh+ydjRrNlLGpo/FmZYFxeCjRdP3+iisCSbAozvRIYobCYYiA0IDBlw
RbNSCBeQ/i+0ONoMwAynY4+jLCukOQfW08SuQSR/IAg7Lu4FRr8F4vUz6ovzwH4Oo7s4MhDAjq7Z
tM1BzDdns2JFc0J6ciFJxLjw/96y5CmvTnzFzhdEorjBtgSx8KRS6U5LYrb+sECKzvZLKSrD/l4V
rJEQwDfIeO8G5HvPoZHO/9Jm+MRFqyOAsrLbhW+ieD7GbUpXoy3Pfhfs0/+rNfFGN9dHilS3swB9
v1gs3ELb46KXCVn4yT0vw+op0XBoJcWjYwCDgNx4xLZeNgwg9ANr1dBxW9gMhAk/Udbqaao1TtTw
Kl+B8I+fBy+5CGSXIeH3K6aBQB1MnYqDUdNcVxB7t/fRiuM14BCq0WM8Ifp/IekSF2T/Yna5kD2w
6Aib4LEsL4jzqBrOOMqLlZWBGy3xud4xO1L5sRwYA6jVR+uzewd7rjqwGdIU2NbCQJthwEi2uvPr
wQINgLpo2pEksHeyfgEWMzxdA5hvKpr3rmGnB0qZD6sKDMjvDWs1j2WAFQTOUcqUpbm9jO82tny+
bP/wutFgRO5nuCUMFLJwu5d8Q5Iqusn3fp3uJXJ2mrXiZlbRBNyiaVYIL5dUR6MtoDjjpqjzx9Es
dV3UIbgD7xqES68tfEVN/JlHZpR2m1uHUgRUXrJdoZ2uSK84/7T5xWvfopy4u+9Qorh60ICNXo9Y
Gj4u2My//naaidHoxBV/poJ8iRRMT0m7jclGiNfjweHiLukJxehcm1MqZSLEoUCK85EL+aSAcMnk
2BqGwLpT/QwI2cZ7TF0UsTy3SFE5NTJ/8KRGS1QmoFQUwHfQTi7uIW2cwYWWdFgATPzwvet9BLbv
okFaLjzX5P6AWtL3kABYtkfkjb0NfM0F4DXKNI/IsIMU3bg3mDiJYO3AMapu6AOHjidWClG865vd
1G1Hwu12/OW0wS/ie82M1uT+l53PRHNlD3LOT66pu+Z/5qr9RFlOPeHeO68bK0iv7SeT6BY84eP5
/wEJRwqhmheY4v+669XL/efY0iFS7jBLlM07L46AdugJTH9c77q13wg55vuzRFQXf8QCgOOYAzDb
yhU9D696+ec7fcoZdAzvLzMlmJJv48GQuys4Hzjg5tB3N8YJMLweV2dgfzLFvJi0T0kT+FCFUfDU
nf3dHWxAb9jFX2YyWdi6DVn94rO3FYmqFk/gItDFEe/SvTbyJQDokRQyJrDzHRoD6liNSjkxcqfe
IKunroDwTLnvPcKFDBk3sWBKP6yP7LqQm9MokU9wNCvJ10g5sY+9Qt8XKYIlh3Dsa06JMu20ow4/
VXd4v4F6MFx/kIvYkByt92IiIX27ZAwe3g6pd6ktl9s/i1U/sQm+bnU2GtdI28ZLo+kM33T70PJc
fEYOjQdqy78vsBe9DAqjKm9X3+WNjGcQ6hwtQX3j8LF48lFISuidyiqK9Icam7hPqVv1KpWueWrn
1G9yUHEPirR9YRhAJAyGv4zSQdquMYwvRJcGx0Jj6R7i1P8vpDDyuWdNPN9UaqLdUG4JA2gtnT8L
Tp08xMiZLRaMUh7PBcsh7qmJsGOgojtbgwz3HEb/NzlJsmSftUrWurnPAig3mYinlNBpSqTzkQov
HDFOFKZC1ntrGPA9ngDhFP+OCfmO+zimmP7dLlv/TUXNsqHQeYlUmgcY17O5SXnlzjtdBgYii5oI
9kiMnxY1g6XK+V65Q/pvLi7eDLj9VrfT+74QHVgbbT5UBcZSTZjX/dlCOAnVcDC+aIjBulyVrP3c
t8dxDeuW1xZA25dbIkL+z/UEbkD5ibV+fH6CMETUlu7n5aQoIwooCRbR8SuXg4ASoP7K01yKN9lx
QW09CGfdC+QqqtaP+SJx9wPVCvGFF/mJzKoNrigMzmAYK2PVQT6bHqIBODkjfV/d2ZDvsPnFqz+7
OPzvDvuejN6OoeZR3nXqkjHaIubZLVfLb2kaCscb/kQuEr6zUcuRbZesKw1KCBvXnGIoo0cAdrfa
CVljOjS+TWM72Xul+kIUEqTIGWojUl9m9JfscLLJUHrAfRlUn4w46CGCkgB/gfDVCkWzY/OuKvNP
JA3r+KT7LnwDIriTmL/z+cUWNG9KBeJ05gJ1qhyBmMwA7IZ8I5/RLSBT4nsq/JB6xUQVIhBfHg2u
vATZTQUFrIDXHE4qZdWLWP6blvsdkG08/oZ8k+Y+cSYZR7D/wou6+3mEccaQtqKsuNVUZJqE8Buk
IvMPYTvwdBfWULxuEyXBJAmAAWsgQBY8mG3lESWprxahIm/f+3wk1E8y2rRxo3XRyZGCtFZvU91u
hKpH0seuTaWAI4kKkakd4f09QFZPu1HUOjGNajAPD3ZyE/HzN1JNKN5JB2ougWHVQx3MccsUld5H
KP5wxcoGYKDO6LRp9NFESKNhVmZyx+78ZXvL6k916jhJyuj2i426L9MmroF94HxFy/IHA7HXwcyo
8l9Y4PzamNESuVQFgYl/K6VRUA50VKvef39rU7pGwLEbPpuRLopP8iOYGFAvqcQ6/fH5drSQffRR
JWEtJ9Efl5wrii6kceheZGdlaArIwbkSUrdtFybRq/Nn2Zcy0bKffsE9mCzTx7XMHgyjFTan8hM+
IRaBVhWpq8F4fNZkQjeR4uxHVXcYSsqnes+yD4K/GuPurl8D/u0K9acGPTBm2qseCkePMYE2myXX
WYXOcyEdv984f0aDIe5EyG9dsFonlVtoz4+vOxeOFoexw0mZ1OdBT1FVGS2RyINDrZOnE4HlNY3h
fSz745wsH6JF1kKbXxt1/oPNk+3iva4Ul2yyEFGcyinFKjo5jRMD0C8v/eStt5QVj07bUk7EGYKn
/p8wNnOdnHU+4rAkfXYYZMcghLXu6RxHCOWVg+zsJGffiRC1EabgYNqf/QI8C8l5ou7jrIiUXzrF
zNnX8Wo2VDpvkH5/jnfp0xrFB9warUuvlrWzoQ3qdVykTHc5kJ4GZR98rGJ5Byol5ZZIZvOMT+UV
CFrvsA3oLo1lSvHjGUFdmiiJPgbWtTls5DXTMjWHWJFTv9QrcpDVAOKwzV63ep7fc1bsrLmgctGB
3bT/h1nT7y7qN/MqKRlf968JNl0ezO8xjuKMqKgLA99n6QPFuT+u1BzDdzQeKp7OFcZMQ+kjqAN5
PYTiLXEtIx1JeosvHnnKhQ5bxbLEckBx45oNDorqDh7U4paNWLI8uoCFwAGjl296nwntZa4SayMi
m/Y/ys+Z6xOlctKSMjD6Yl2aeCrh3CJTNGQhdDh8wNc01pIjS67iS/S0SEKTQsdA13OCpJgb/APU
KI8zTzk/q7vDNZKnwveLwZKvm4sKjoPwwBo4NReTvH2QpJUMOEdJ1vQcOVe0ywegqkjUAvtPUAr8
TToK3m+ZghHj9crbd2oG+Eof8b0/rzTJ2bQZsbnoriDT3x1rul/XB/hzaldkqE+F78/rtWSeclWu
bmMfTUke8sQPTYXeN3TQ6A/gWvD7mn9EwhSaw+P+97o1bsz+v3G5Dakq9itznAG4Fh9U4eH+B/Yv
inKlo8yZV1xM6W7Z9f5bx7PbeElW8OadoeYQDNbbKpZrlOKb3wFFDDrpoFAbAlAf0vFareyJ0H9w
H2XYN/3qcwQgApocQq3PiBhhn7pvoB4mcV7Z5YqqAxzKuXh9I5sXzj3KK1CVAPDSBMDekRglfp1E
T5HQkj4B2tHlXckAza5RN3fnPTw/87lBGUxGsDwK4ReYYwEIHvyAqeZficVS1JIC/9jVDAolWLpk
usFMa0zueZGvWk0hZdLhM9w2wZqVNqCxgP7wLXxdLXaOff6QwxIoSqW8BTNRBslNopenmaGluT7I
BAsFwvLOj5cjXDtL+Vla9XKq5l3q9nuZMdtEIk0g6jnCSIGmWUgJc4dUzQqV2hzZ0lYyJHHoZX5I
+Xv8o8e6ADrDuN3rAltVPqaGLipUsUQvh4WZ+2cSIE1Wg7uKyiQwVRwCXvA9YjM6mHvbHa9COErY
pG0jUhTasXljtuTkZMKqeyfvd8Yu8oWruSoAyEG2NACH7jmMuMgR6vI702pmgWvisjq3Cd4VQaYd
bKyIxIin4LLkInuTQ6at3JfvPyvpQ4ToFq70fI+iG/ZGRC1/KHO8xDgSz4Bg+CDstnOQ1qjO9naD
LR8n1hoVbks3J6iNkDPzC0bG1Upyk7WDnJ3XDjf3FO7XvKjmiX+h2FICyRrES08pHP30Q9M/kcXD
QFTxd7f+I0OxJekrPS/fMr95bx+XjlqvawAZ0ZTWyVIX7GVu2EpPBwFpaXryqb0CCSFN/g0jJ4Q9
zxmpI5QCpq1S1hNAVVBXZ9cLoZi+IhgfQhGEmiMNI1Aof0ypNGTjG0k1vNDvH9XENzPnBJgeRGye
qzM3kI7N5++QWAJ+FKWPuBhWlpxXKMvtRQus42RlPZ7Au2F0L7rfZ7NE7hc62JUBpqlxZCDq2Hso
BoG0NvZbujkjsdAyn0cmLH9yXiqgYtwwqghVSnttWk+Yarujz3bdZlAmSPoTBeJAAIsP9bg8Zsdc
D62TFL0zHMuBiXVJDwxy0piSklrbrR9NVJwkt9Pm9Ry/AlXmFzeWz1Q9dVccKGGzrG9GcPcD16zJ
75CeAUUUPQ6AQK5OUc6pNNq3iG+EQrE36Cy+Q3mz6Hcq+BlW0N8/M8L4qULNWKlZj0UwxXSYoeMY
tyacBar8MhSvgAqY2wAuXblTzIq0dHSsEUjbBjDtS98bB9HIKfzFbYe+AxDthi4e5Yt5ry4QvTB0
pw3m/11DrOTQ6CPNYpnYc9OfNJeaHfvEggN95PdDIeGis91HaQKOITKOOi/rd6n/eDy8BMn+wH7k
cI3iYUtK53+ZSI+R9kSF3U3+6bM5Rlpt/QgfaywiLZ3GAPllwUMxqPC7C1zxSkW3vRAhx+2Dlk7o
Db/T7MqgVTYPoXAg3vVrvZ0UzoX76E8YDdMdoUz0pjG1aYkSHui+qg+qSoSdmrh4OpgnWICeUmKY
bQ9GCpiRnTUG3KK/f/QUJlDPT1De53Dx5QhYPwa+rz/QC+wNjkk81USpXEHiGBZckuxJ7pzpBKyE
1VVeIHjpER9cKCP+lj5C2OLHIlRgHF3ypKgt8O08RAjjBjIJfqfyDDacZQ5pnCCvWjlCeKsWr69Y
HZSwKjQUOIOMcChNnaD/Oq/XFKlhNpVCNMug7U05Y+Z2+Tp5Icv477bPmkmJ13NoqEUEi75Zumnv
fgTK4NoPjNyRs0lNHOl+Kgaq43Q8bFAw1hsSd0QeEIMvv5p2xfmbqvsuYgDbLLE7ja2Dxan6XiL8
VuVE+p6U9gEU8Q1klR4MqjrNce7RL/Px5hVHPf7+DeUhwugDGiYP/NXObcctObZisVCBC1DO7rU+
lXJfmFjRGDh0Cgf5g5T2pF3o2sdCe0WqO2BLhAYskQyWLTG274oTaIZyQ6qawJiwbnTicZyWYn1K
QDzqRaJHXQ30k556dWIVX8VTjxDXHHIlvjpIgk1TZmeaCrf5glPxVAm4OFI8dtJJqkzOZEMIOSXu
HqG/3k6RZoB3Ar1bO4nZ5nKbyBtrzU9LkrfxsGruj/iqcTvb6XzyaAopQvjJZRTO9lSzSgWvB3Zo
y31Gu2HT6ubNhgrKABDUBJF5Qx2fgSr4EBFrLkJk/52+/lw6j3QLmb9d1Cqem8lvwOMRcdZ4rwpP
U37FD7GJvAcucnMj/EXkfkTGp+MRKIo9h+hw8XSQV1oM+pjzcesAwciKSHHQty/rhDhIqsl0HKqI
5+Y7fqlwhGk3DWJs2d6e++V4zGj+xPJCsTtVGACLfaiLPLmGn32S4EB+nV7kWfObdiaYDvPvXwhM
V+dZHTWkDhQ2hB2Y+wDS7lk3vJec9iI8ZK5PaHpYdkdrLys9RFMzFbBKPT2vkRa9GDvAxNLgopNW
UhRLsS/emVgTPZrdQt0VYPfXiw9J6mF8dG8VKIlWVerRRjgaWkXLu+eimf1MAhw5E5ZXgotT+150
ntqRsC1M8pSpsGdr15BFqsUKHdTCZIy7ZnRI4mXs7YAnLT2Ww5AA1BFJ2qUzQ+um209+WPNWHQxy
j0if9OsGMWEdnIajfU8u6EbL0BnrbOgnzP/eSz1xf67rU0WuEsfgD0yIpmbsA1fl9sLbrxhQOvH5
6rtjwVfn9Naqp5zBn5qvV/fDeq4p0Ma9iVrtS8lseIgnsL50eqYxWA7AJ/TvISBWAwPkexCGIVsA
q5WTzfeo2qDzUOPFoaerjmn0Tg6peUjIIoK7RU2IHUXyxpSJvwr1LvpXkUq+N5SrR9DfzceRm7VE
eACqdNpEV2FhhRiKcBs7mViYqH4MyV+6QNywUn3EJm+O8V5T8187YhxJRwmkz7KmbQVEbOWrpMI1
coybvQ7ChMVRdjRdGO3NqVB8KokYXwns6nOQ+tvdHWRa2dh0bik0cxEV9HlsPXoM2gts1arSYjmr
AIuYjYmnf/d4mmB9CUv+Ki32kqXhzj+UR4ZuiapbS9KVzwQuNOi3wKbHG2fimefsfdVAZdCvW2P1
2EaztzV37/yTwGAIIrEONZQawUQR8PkxclVa1qKV2r/QDc8LKw/hFFv7l3MVpG/VQFd0lra++z2M
pJarCy+3Jgq5xC2q07ySvipZLzm625bdRPdJYlvZ71UtDjcqIW+SFZPQdkRiI3VtWWfAgyhZwDiN
/19w6zkLw6Jhnfim5LZK25z2ihIfRlCPwQXkrES2Ze62t2YX5NuSTr7tkHeVKWwxhmhUbHxSXedk
V6luldm18AYLz3Xl29sjso27ydfB6QwqHypMaDEjGRpXv+FEnlR3t+QbxhQdMAhhFHxkiMQ4+MHQ
+8MuzcnuKUC9vAqL0eFvfaN4dcwOYIdyUTPB2BxR/qw0oXPdAmdZe0N2pzkpDQx2pxhHLuySdp1i
bPXkm2+6uCJfAfwYID+R+1v11y9LmfrGN2/svFpu4qJQ+x2znRiIm5kTSles+lz1MVwJcp3a7bhW
ns9Iza+mPTYDgOEusgtbmIGFuKGFEde6mwrPQ+l0Hf7inUqJZEhND4RFUpyNloSA0lywQqlKmguM
PH84faYSQj/eKfGnG2nI0KTmT9+4R2KsgusuxyQzW544T/8KCD/X3AE56aAek6TLk9BWRi2L6oDD
901q51K9LU66nl77LrGBWdsYE4CH7FCbbbCyihaia522kHvf7YbOTELBfSk13KHVYmcgQvC7byfL
Rx17OU7/Yhr4z/Nr3AWgs25iDAkBEqvHXXZxAObNMlCAd//5oMDVRy/MczoqQPRGBKvFOZbhGR2x
v/sCq7rUUr4sgCMBTnJ6QXqHI5y3hXM6ySV61xZbxotKX2kERypRKXU6gwgZULrTAPBUzvJF+1Ko
MGJQN4rv9Xpjtli6S70SXca48CGozJBnMGqLVyknj54oItKEvXeXRuNXkb+SI+6CPrkrcqxOA5jU
QYiM6G/qriZRQeWirwPXjBf2KEQiwrHMrCfqkDVWNn2yNdixum9d8mmpgwFiQ+KkNMsh5FBSxmZJ
qe1oDMysLSYeBK0oQvO9TywnmeoVdd8sMKMUibyaS7m4FJ/IiVDtDr9W0KB4eBxR2BRH4vXOTCCG
r8CiPX9783RY0fWYH5Wtnz0n3Suo6nCyGLn5yC43Bkp+U2yeXBYW0l7lfqsbvS6bnu5L1Cdsz/Sf
M9CBlwBzysX6l6OlgC8slUJlz4af7IHzTNheZeB/ikA1HYnm2k0yqS0Pua+BfLM5ki5BzzIszjz4
6P7FSP8ah12kPOyIygMkGVcTzHnjpg9LK+fxvCEzZHZDnN+h2K0Cab6zcIO/TcCXj3jqyMI37zOy
p7gE/QW1C7pXPNWA4W/lDgAsM3rlRdxCN4ky2ztGfO6izlI585Vj2p0ioZefZEe9d/nAcJjuUPq7
I+67TuaollH8P+dddd7oje+zOK/qHE4SRPoza7Uy2sOfOTjoYeHT7gFsXlgy8O0/qRoRGJYSNQsF
wc28VhcvfOHWkHq+9+00MmDq3FO154R3KzYAzZ9yJXJipJ7A+LUz4md+Ub2CQ5z/8GCXcX03piNF
oTFACwquNaRHQdeukTPOqzcb9+Lql9btvPw4cscUnwoGHwcwiZT1SdcMMnv1i8IKXnMyueidetRh
ItPZMypcVeQFXjY2NI423hKfUNjUOhrRo/9RkWf2LTlIVLwI5akGuDyucHAaO355kNxEfWi/HQoD
YdlFxYGAArg5kLPzUudSwp0Xkv2WmGG+L0mBuYE1X1bg9n7U0OU9Q+XXqfrifmmij6c/G6XteuR+
ysiZL3EdMG5p/B/8s1Xv7WpfFpfPsEgkY+O+jU1HDe4pKM9s7ToJFAzI75jSx99QEgubK/iu2Ooa
CW6BtiUURZ19ooCaX0m+IEwcfQ3T3g9GTmz/rWwk4K/5NXVwaIX9Q/RfFCHSSzujak4C+i6dxzmV
rUFRtrawq/eOhgvBe8FYruFxgkji3VdFh5cwirKsRlJTw+Qvmypf6sGFAq+RoP5Uounf82kc+f/a
Dzwn4ZKtHZPv+5SBaXGiuuuagMUz/0rz2fuIGdpq5sdVWoLuM9R8DwcwG3nTuaFsoKpLbpCbfp+c
DQT+wvRavd0GwRDU0LciV1UkecazggGPHwFCmvWNQRJiZRMBT94eREQK8uAMxRu4f9+X7WTZapJo
nAeVoXGC/SnGbwRSpkbmD7xV2DOOfdo6FvgGdUWEDf4pjZYM99WoBmGwqe/Lw+wslZ6ckbYef7cf
uJHzTG47LkTqfrZN3c/wDEfB0ixht4uR5urRjSm41+Kx9C7/CdOnm3p412CJEWNivcaB0Fc5qvSA
z5aR8NC/UmNpG55obuZBPzmBkG7VehvUNLjW69x3/5JmI4BKKVerCjhwPabDVVXXQDcFTY5RvNH2
yJXo0iJymPhz0oYpQSrMDr1nPkJuCk3mvORH3NkvcnfT4KKc8RjmXYcqInZKIXnm4FBBcByBSP1G
z7yox+IhRPJbg5/OTuk+d4dReRbrytB5U8bKmDZXlEppbhBs0Tw8jRpgT5WN/tNc5KOIuPM21Eav
bst5NCVyMXCecjEMCdSdC40D6fIlLFrGWN5L4sjetZ68K+lGXWe0f+T6DFYPQ0bCbO81nVWrbT19
cJhFGSehKauK5gw04OcWL4NhcoPCu2V5dv3AeiSK0hv3LzN93gV9w2UOolLkDTyqjinpLrMEMQ9l
juFVHelSFBRysdT8eW73a8lMeo2AG4n1mLaGmudN+mPIfBcvtJlF96EgR+hOGMVCiLsov1hEDkJa
tbfcwTlnjexjA0QAsqNlw+yPFYjN/oDeFMIRRD+/W28EYVdFcUlPQ5+vrtSF7UEC6QKeXaVH3HZ9
cyY1oYyW0p437w/PfBmv/lZMvwAI0UCD600t0Ct+y2wNsCPImw7S7fQkZ8cLnWfYfaujANq9L53k
M2Yk36rQNxlhC1cMyIiCaKPsgFiyEDqmGLU54CgCM71WzPZXYFEeypnvAygBlgMpqBbfmhdCXsGj
pTOA6lHr01nc3r7kbt+zapyYHymIWw0Ub+yLmqMfk8xnuhYTxRj2g9tRBxdlHr/k2ZTu1cpOnJK6
Dmt/uYbMXaQnsyGSN/v38/tbOeul/iwA4R/R2RyXBaLzogsbFmDDKDYDIq4Wa/NHTQkIgemJ+0ke
IxN6rSaHVtGINJbsXOOIkTEtuZJ0yyLA9Bqo2l0QQDnosbrc2CGiBIMQ6Hn02NmPK0zeAYGoKtfu
/dBeNxGis2m9qMxS5rk84SRjf+5glTEnOvhxYsxNTam4vdX7AtYExUSOOxHj6xVqn1KKqQlzVDJY
GL5zKt7BXFnJX30/5AbgMrXcDni26KvmSrY7Szp0lXTBOWyiKiBIOG9PDOFX4fhaqmRYo5/x1zz0
huKFuQGWaUJIAHQxn3i8RInRMIo1djaOHP9KtbePrKXY2j5ZlJbBlhsPHi7QaIQ3Cg6jVbDV3aNh
1CHIXqnBoOSQK6qKXzbTYMY/p7y6pwrF/wIwduLA8n7Vlv05B+HVAgkl2k9OsTvFi5lBqhqiKB73
tEOeUa49ypl5Ohb5Skkqjez+Lj0+juSpB5H1KWqXrzECe2GbNQCO4oquyM9H3N/2AnPXsI0vxxwM
SCCCjUk2iFdJsdEjfK5UCH5Ngr98R/iBAH9eCIYnUcKSqTkThEvyR4L6MXDz8l/wFdBp2HKfUcJ2
Mz4RUtcxrkj7v/BlY9SVgXuVWGp9pMyuhZdKkgllzi1pp2WtOnxcBo1ECP2R+u9H5PYTwAwraVty
yUSIRQGXA8gQTi/YsCFu/D80hzwxpfQcWNwrAuHyMEpgk4kXOPjQNg06z+hgBAQswxy9QQ3tlKa1
T119+xiGKtkVwbc2E7cHfhRiuu6U1AVlX9EDY3RTvYg8sSMg8dTwXyjGxrUNkmkFVTlqtbD62WsF
i/7t4NZ8hBzixT7AOdfC4smUUWK2Pp4wQuloaqC3tW+sMvBmJ86jwJ5kfqmuo/kuQWJuac/If1Oi
lcppv92HlCFTfrtlzccdPaolOb9rpcjKtnuP6KBYYWRN16vNev9/YTaRNgwIMphqHcpjXfJZ+o81
XjZoFRkhCr2/vz2veZ/ikhHrdZe/t19PcMPZqFvz/mkbwaHezd5fz2IySEsC5h01vH34v9yMHA/u
ELZCdkjs9LL+iHmvQvQHjBSbWsj/p+mNlbn0ivovcvKgxuR1BJS/H1e5kHXlYesLbdvwvx2EVZW0
926ZRCFpUdTJ+5y2N2RzYPifzSQLlbBzeUByUeqVfn/nZ2YRkoMIRfJUBDjM6oYvAv6NLMoXaFPl
TGYdNQOQjZL2fbAODyOTiQxAZqzfsMFm1Epk2GEmQ78UkgRir7ZdPPNeBnz1lhSv6upgw9tSTZcd
9uXGBaN3WYwaWekCQt4/46mVhTH43Wm166iKUZCo0A6iw32BklnsdThTtAqYzQBdzVvV/AZ9Dno5
f1d8TO1QnmSz2cdGj66g/xmU7Jxer01vUuvIfkyVwMlaDvRle6ThV8wkXJ0qBln53XKsDd2LQe4O
yeI7+lzYre2ZCUh1ET868pqrZtoMGV2CEphhWm9nvpT/a6VIKJQAHPc48qRdziCUDAyi76jNNbTi
IDv5U61ViCLSag2JLVEfdrFtgtLTplsIhJSMs/AXgpCnd6cfVxiR0QgM8gjy+tAaJDYIfFw/z4JD
NSPHjfZzDx3qMfyuODIQsUAnj+zoCbpOWssoI9E38wygSFVanAfGWR6l1YtgPKNtPsS2E4I5xMze
nIj0FAFPEmRjAZZG86eHg74KDd1jEGeqf8boeNEIJi10IOBtbyQRe8c8cyBf6FAeNm9Zpj8SHNRD
KULKajXE/YL9HZ2N6zWXLnx1I9NkWC+HdEBUKVYbl2lBcRi3+/odyNchecQyqLtImxdtEp9/Fgf1
CQgcH1XnzWzzObikGCbH/bxxf5fH+bcb/Rsqi5T0NGuk36arhdT6SDJRL3vUkIbBDHJ1uj1+ShZU
56DfZ9yq8smeeK7/hp99hClSf8qKPH6BqJ0daCHDBaAKr6gEFeFcMJBapc8b8cFb1GQjxyM5SADA
Q+5G05OisLqwHhXfDo5Ij8uJI6sM8MFJK0M5C2mm0fbwvxhf5GEjoQobzM51zc8TUj8zG1kv313k
kJhZ6w3FcDHBuvSILwwT8dGJjXZ7gNjBZ5ZDdQ5yA5oTgjwxWkaYVK0Aux5+wIYVRLhttxHgLpxu
NlNnVOjARoQMhbeDrBL0MGHoSJO5457B9x8ltTubhVNw/Phl8MDo+25KggGQM3ermzOx5wpUeHNt
NDCX0kh/POYmWO+4G0EiyZzECovQ7Iec6xXdr258xgeSFxEEwmJFVWHQuKApgrcuF/zOht0LwDBG
MvLe2ukuKsw/iaJveVJPbqLdnNF3MjU4+f4NZP9oFsJoDa3+yWkDC92ffWfHcT8rhVcth3OIOXsp
Z5jd0kSiFVrUVv43IZhD8ly6DtacL01tHE//2od5u6gOo0vfuzoTIcEjRORlfe/0989CEoJIRn2R
vS64BlxUDM5LU3O92G9H8ocUm7scxaYSNFzoJXxdo+ibXnM8+W14KqGhDAc1syKX/31aYsLL3KWb
V6CJVhbOay7TOG96x7Fg08N+Ajf+Jh2US5D0MjxnamXNdf54eMS4AOVWKLCP4nClTvn92JBDEk8p
zfMbDKWmJIvNa+IeeuY+BGfURHaphznfn61y3RaYGmtIGZH4ymiFqxfadXHJV7TrNtL3CNzmuk+/
/Bykhgu8Xle3cGy/FkSI/uWQwSrHGDb1rRCaniLV1gfC0rjiA23v7ZYBp9LvpE6ECZOWh1NCpWjH
8jCaKNXoL67kD/fk0cv2MRnv8E5paoFklChNxOidA7+/KYqEbN5JF0ySTTqTKO8r75ghfWkrUMwD
zJg05fFSROvVud7sLl1LMkIKxbqcQcbEXmzBZ/nubUuUD5l4Z2pTlglDOqOcPzjqC9ZkrR8d1xtv
TCA58aQs5hM3erRz3zBShHQRAxe1w1dNh6MPm3kKMm9SBV+/A21lX2eFxNI+DTZ5uknAVpqv0T2I
OlgOdY2QDMPLMKehIYc7CoFR+sSfhFZzoGpseOlnhwqGLMgtRh9ULBqdWGuvLmSuhNfN/dEI7oZ8
DLU8MC2Xn/PBrheWSmx+P7K8Fs5PRhAYUPVSEBfE3nyW+ceFERLMFTL01ijNH8Dp9Jz+7dAnvi0m
1hhwipDtV+jaYUg1GaVDdUDisFRj7Q2NiVWvcXKA8kjWveoURxzHZ2RBWtqwhcEqLTO6NA9aTePa
TaL9/dqnecu3gdHRhO5u3h4JwNNGd1J0LxxV4hGTsukqVfPdy7Hiz2r5H3TTAVAHlklVo4HEcnty
NpLcflcl0lyu1gnYvsji6ZBSQTGlEtJ0fI+z0y5SssIh+/uRcX40E6diDa1UZUyL5RMHm+pm1LIK
7hoDqzYp0uzCmymgHOZXagNeUtpSJ8LvVxVAFNipG3i/LR4kiFUgKhhTssSUDi+sMGh8W6EI2tJa
AExvmTEpTkTfpwiHRk9NyAT9jfYMh19EQYKvVLj96LEEsVkrJf3BaLnIQ8C25xZKn+uMSbmjko00
OQk9q8qFwC2iLmc+VA37eqvnCCbwSjQx6FG4QOIEzTm9e1Hnw4AkfZRWaG8sgE2cYo/eQsAqfLod
bA/eOtWArMiF95vZxW+CLof7a37bwXOVEt0VlUlWonudPTJtMdy4+fWDj12uTGXxIUVLIAbzSkPw
zJu2SRiPDdRs2NdirUJO0u1AshXvWNJRtFsfxcOlNLUcxKW8c//7hxAvqbyRRpOhEvqrvgTPIkdp
JMbVKA0WQ9fLmBZEgAJsVyJXrLctnwzjZ+N+iXq+0JY5jFkFGdczMjzO0TjMB9UdubaBjYZXEFQI
4Uw0jB0DE8Q+rjn7HPJJkuiIp5WphoMKIWknlS6hkaNO6A2WTODE34xtvCFOGn4i54wAIUikUQVH
qhVFPLFTL16+UVLjxbuJTGBuUOtXpcgOYgg6vNa//bPesOsz2AbJF4QhZufC789LqrXHn73L61Bu
fbL04PipHImVngEXvCERgdjytpcK/xb7HKgwtdYvZHuoAur9eTMAGlJETnt6egKUXPEmky23dkqA
Z5BwnsKybcqdGlhJrtSlSy4c8BquK/eAXPN90FbYsAyIvIQjonzTPXrzxiys4rMldPusWjYjDfpn
OOCdrde3xGHQCh5AyxgXPB9YfhfmpRNDQxd+CWaGTTANiEyLfN/MsXgMP1mnwDrVGtZH34v/Rlz7
8BgsFLOnZnFyQ173ThwvWByM0yNWB21NcLh+w328LPWAX1jLUfA1FMLZGGQJO6xOl5Scvw2P6vaw
2uSuVla+x2w4vMrlScRG9v2y8vHH61uPqIY6SjiAZUNx5sjmGe2Umu0Zcnp46ZATGgdGHzSHxHl7
cOh8IEHILFZJ5mipTnSd9rrEujy2pXLLokyEOb8IwyrpmoFWvS3+p9Oj+SG5xvICwzw5gcJaMs3+
OpnyAqYYRp7uq0OEXhTIWY+BfSWCRWPFSIT2WAOtpdu6i+gtg2Q2R647PR2bgIWGvv+bi+fad/7c
b2duGW4Tci1Nh2zsK3dGeYsD1gmdTEjvBUUSiBSzOA6PwhXeNRWE5cDzAg2oOuij+xO++AnmonP4
mjPg82qFHWSOoahmtHu7tBer3JcG57T99LvCvMd8GTZORg3tzAqZr7ADcXm+VrqpB/GnlGMd51x7
fEmht8yLqMfRCtp7kYcS7hWpGKzw5GWj6kxXLxPD89YK5gyDBImgWE49i5g59E7jTKMMrCQ5DVQO
Lkh46fO6tgDgGV59SuYxltDBWjx5qo2DSxEl1HObNYVCN3HMOBmgzQUdR9GEQeyB8T5/gYPJuMEa
VvTHHM1gbwHORGpfkQaHudPhA275fAD5N1Lt9QTBLTeyzf8nUeuxssPGeD1bB1i2UIkJ6WYH7cvK
gjkpWLBlygvxVTsp9x25R2FnUBZ0XpNroW0xThDtG13AQ3J8CD6TYwpcDpGPFYOZMcnYdRIRlppa
a+dSobyv8ewpaEXFhQtVNr8ushgcwCwzG+cj+x7xzD7Y9vWbguAJefaSZ9U6a5gbG/CnqL17vVCj
LUdEdlJCqPFNpyXzS8LtNk2qqHhlhGTRhlbrSBW/qWhIOyXlYjB01pOaAbDW8yIBznO/uHU0Y6yt
UvzPtztT4Js29Lse5XeoYgi/IjdSO7BVWkhqPOOOWUucl/6B1Wo89Ub5hXrTh11pxc0REvQBbAyI
6Ic1uKKR69zm2iknLROD9Jkdk8xDlkLx6tt5hGiUtvgF51STdcsaR9jK6heABQwRsW4NToLShura
t9uM/g6VgFIlY7SvqtJ8+xa3kVuPR9+DTfxWnhb3kvm22Mn2+mHzvLI6AUqOHP68xCgDxqbKjLho
DVHnDNS3wquobfg7dIO/7TlyTvpRIiFO9gYxc7pMTEK/0Ck9wtencVTvGKwBfrAdLoOnhqHzhLxr
mV4ylD4Ue/ThBYIs4U+fE3nDb2FlJfXo1wzh5iph76fZGvQtg/XEu/Ccku0vryYVlgeZV927er1z
O6NlAdEKUCdymK1cDG8QihuALbRA6AGJx1qKXN4NJSy2GR8iTJ7NwZw5ZSICU43cN9VUEW92QrGN
i02JE3O07/iPL8+T6Ell7qDKQc3juhdi/gTqMaoD5mhtEibzHKBjkgDWZNYwV9oS2KoQX8L4rtZR
f6EKtkHW5d97DZwkuZo+1+BHiDfcOGQhw7C2MRJIknheTMzCRZISIFLs4PbfDYU3T1sYCQrBdLDS
2nL7aEuuGR5WLPtgzI/LP+oIDuGP6axFDnuVnt7+PgoAW60e7uLe3psKqVOXYcuIU0DqBZJicpQW
472U6YsOf+m7C7SAi9taxMawf8DYb+D5U1PVD+krfMFF3CN4EvPjdQ+UqruVEDbUP2rVfDmrJSAm
bylwfgWfyhgBASAOEYyZRe1fxjsutFyK1cAJIsbJX/OWEA1o47jNgWuaKw1jvcc9iQS9YDs4ZDbe
wWvvTXsn8gYF02gMMGZDrxbFpLeZkqe3fPaCOWZMeDy7n2ZA64Txu+wvlQMDrgcIfififP1SgZ7j
OdVKesTkE9dTK945r3CjJBT9zQsF4uVXuzuKsZFLtDzSGH9pKvewjUuVV1Qx7KSnVL3iKdU1Vgw0
xkJqdrTGEMkYyfEYj/rr5M6Wae5bYewwc9VnMVhY1vMbltE//2zpx+7WA2RUd7FcnFjvuD2FTUV2
tzXl9+xfNHpW7QlsFJmu4MyvSIKtBeHO5Ncro7O0BjxA0WvNHl+TodDkZeeQbz0W/SZTwJSFNtgA
8CQ88TQ19WqiIPQGAcIxc6OSLtUvYVpB3H1YqSGbZXAQdQnsraQJ72gcpXBDl8uuDKgaV6AWBmXr
KBgOpK7IxTbnGgoCP/6bH7QNuaK1+kxS3g6aXFCpQ3CuEl8lKCuJ5g9JEEiQryUVyr2h5TEmZNNE
PAHambkFjnZkKRm5Fx14q5VEGc62/NLv62BSIJciQDdFq+ZFmam1Df0GUi8XNdCRoZOYL/b6jymF
OEvTIAfI8fKbq8EQF0e4xiaaLhjz2rbP9uRINPnd3OCIqLLcpHstpIMZmCyVAAacIKBbHNlPRAj5
dZXi8m0OjQYtq6uJxFktIfipegTrJ7/zy6Zp/kqRiVzFxpldrA+3GxfzgbnSfESWWjO1h6yE6xAT
Q8xV5kZyb+Ba+Rv957EAK/uW9z0K48LwioA1YnCu5I3Xxhk3inqEV1Xm0Q0Fkowl2ScZSYzc/yny
fcddFfG0A/CCqPElq9s24t8Dz7ZRO7ec4J6eZFpHkawKw1betUWLPMOSTh2eK0ILsdZkL/+rUQNi
chJO2mzf8fBtCY7SkLziEEL3AqHVxzb6VXgecS2bwsD8ivFwRqPqNxeRD+TTyjmttRGABN/uKtpD
ojroyD1THLn/4ozOsTH1Ljzrp0CYl23YAFfZXFQF0Q3EsLWwsYfiJ+aSOyCoMiRDlNzQ9Qk5NFos
H67H6cDYiH5OC8F9JlEqEPK1p+GssISjtMMkDCjjoDum2wOv5QqVmnok9omCiWJC7Py6q74UPBz7
H6ih1ohQ9s2K2Lhnvk9mp+Z+zFiy/+D8/IqYn5uWOY33aWi8+bVG7npMhtSoH4x7PC7/f9dTrP8B
EpiMk9Qz1LQDDMSYdjTEV/LQFG/84OF/Wo5S3SHu9jgRHe7o8gmmBdiiuGDDKQZ3ceM7z2lhPUHw
v8gY1NzQWP1ruqZsvUtx8fPXzx+oFlk1BOIXpn2boRFZ7FbeU/CYWkrLYHTVfZvvi6p3LhzUhVi3
dx6C3o3UvnmxUh7Mu6rqREm3epXiGdC/WnYztJnUnLRQ4C6DtZhXji7QcDDMACNG3lgLyaLGpVG2
dRSSbdbipsdp5XnoyGgcGRyxAeyUYFqsjNc13BIJgnbfLbX9zS1PFmGKTSQ6hfsJFNVrJThWODlZ
2zos0GL0zQWsMl8XNu1HG3wm5fHJj/iC7VgCxB5spBX9S6FR30y1nWMjZDNkaLWYT9KUTA6y2ubE
6LaM/gUORXX6DVIgc/v4V0/j6cwMm/0YACNMa2aYCk87fSQ7z0ePSDtvYdSMly4/46k8YoZzUSTZ
f4pNyfNFnLj2Jxe0Ky/HOvqh3FKjjLAPqORQ8p0aHeYYFWxHGX3Ua6m0E8mI0QiZ5N/jIG7ysgWp
Al/XPOCy+gkLHtVVn0esIXBxsa3NVxB4BDHWLvShpT2tDrgzWj5GJs+mp7/05uOpmWv3NwzhKmn4
GLYIme4GQhomac0nvRpOVhM3GlAxZCQcyrhQ27zSiIhRruumb6XKG4S/ZdCAsAA5/f9HbpTUhRIR
ujgKL4t5MMpads3Ddcztw8aUC7RiCg6GpYRAq3tCxmtLPhqB5xajqbezH7i5TeRYfOXNCAkSVtDF
yLRq6FhPi7BGNS22hK0QIleiXg8bN3DAU2DMI/f58oZPdoTewyAr7egkAP6l/i5DNSVFiRWHnip/
J8dk6TK4IFFXOnDLyCYLHkrzPrJv1EzUk/A/WRAqjHVQ7iKtM7/CdZ+SFp1hS5MSFI4de8bhLJdA
9fCdQY2K4RU4mAYq9qBj69VAQZd6nkB0p+KEUIDfRp2gxO/mITPQs3K3sSWIc/cn/W2EiQ6iSUXz
HhCaNug8ki0YDFMERR4aUa8WA6GGkVTP7Olf0I79nnGkuYXtwbBIUOiBlqTc7EdAYaCDEsaO/rFL
xPkeGAi3XQ6t9B1mENXx0lYXjQdKvZuRBeOvn+BLucChwYmUyi6QwBY5mSjea/Ec+ChVz5LX7sH+
2FXR9qIvqric2eQ4iRr75dtgpBoqZ8ZwoJ0VSwXvgDs3Unf53424tBXMTvQPVz7QD63n1t5pt7Jj
QcmM8JL8xk5Rypa9cVOazAfEq2cvjvR5Uzi3FDQfayv4IGvlDjevY5MCYjVT10rUlNBXbQAw63kh
g8lS96pBbtU/psZBVfIydIQL2wFC4L5+EcND8oFyy+1fiN5iTaftFgcMW1c7V/klQ4ADsLJoQmlK
xT0qBLT7zFr/VCVqI1y5GQnVL5a6k3JG2yfLHdbFAtJcGBeTPXDgw/RM48s9NhbLmTpelKZriVkY
l2mLHOqAiUuy4fe9rzvm3d/2sFeC4+moTKQ2bxm+DTeWHt9gUzvt38QoOorUBLm3VraJJ0GVGUIa
TTzmdukodjyQZAtLl1C/vyBn/4lRUfTeRpy7+FeUXUrZK3ynPZeAe4Tnp7pj9szD9CwQrDSL+8u/
4/UsEZmL/74L8V1Wxsivlm7qe0QIHoqbI9KL24QxnkALz5duY9UrKZNcb8BT6P/PzYqpMPhbzO3g
7tox+tQiySyWYjXq60ohU3RtxMOw2DnYtw3s0VJ/elYM/uJbGJrMZh6yeNkK2GL4bcJPyV41XCUK
log4nrKFhypaPAhPoGcxO66iw9ga3qJldQBc2ROgxVakoVCuWYtiK1yfLxEZlXrUXa4zbn3veIMk
P3/l0vIPY/eMxOoDAE2mtltNfYEb7+iz6P53veFZiFOuD9ygdFPqJsPVmZ0Iz0EtZuIH6o2ppuDS
4D/PBWjNjmvio0FwgWWZhd0OyLmJekE2BhooqeOQFm9rp+60SbUgK7orOltppkZjH5Fa0bQeMbC0
nHCnWkBqQ5v/f5IwOUvy+iWD7DiqrS4o+7gBNHFGpbAETZ9bMtLDWyemx8ZMtIiugfPNuLfxJqB1
GQL3l7cjw/l9XvCWE4ePVDCpl1+AITFc3gF0nPehtSK4GAcS+omu41LoQ/c1y4IwozYm0SkM5OSG
7F0bWPMSVHqm6l1DPpEm2ezuVXdX3DB/oEh6qpiy8Rv8LEVxtqS+tkNF3C3XGD6JoPiqVobGl53+
XsNemCv53J4Jw17k282JHlSVs59qj4e+XxK+YDGqGNpavb/CyQlDrLsHginzL99ew8iL3d/yZHOQ
r44ithIDCjXlu/9lPToi8hkMbPku+8F+Jv9cYIo1/5XnnSjRXUYY3SWrqg7TTa4Q6Xiaj3mlF/Dw
kqFYEbJQ1JRR4imUYgycbod674yXjuJP4VHRuOF5yG5YxRF5r2Y+1kzc1vkSAHn/4qzGI2DG5r/j
oqc7k8UOK62hIRyJKnLNfvcZNbUwkOmvaTerreDF++B0IiaOBnXKqIYobzW8cTOlGWcJC2iCuhJq
QQNdFUcj5RBK2o0qicxQilGIS3gC8EMh/HOog77AAIEOrS2v0zmnzi0kg+Fv7eVlzvASV5ZtXTm4
woCUiyx/WAPQ0yIeQU1yVahIsA4DCv2EusHnEZ4mUDphvHrp7+r46c/idNnk/I+KjLV2E2dglikv
nHInpPHvpGIDoslQgANbOB8k5cnfBU6Q/PKCX/3XKRv45zQf19cMILJOPrHzcq2YYXdRt83yWa9l
3yDXwg0eYoep3jJNr/58WKEdEcfUUUvKUeXOOXfmF92OqeeBSl5ysThTT9yz4iEQXx7NvAGs++qU
Jaa35OVdxL0P1LPht/TWVw8MJa/Bfip7oyYa2CE6TU/ihcTjjVEqXjT64ZRsKiyeX/yGyxQD6HUo
5fnBMSGlvyY8ye+XC8eOIJOhs4fHs5ee0hKrdcVBbcAXHt9XoFdYdxDdpJQgJhJ/CZ2V4VDaCgHi
4hgVlW9v40xRsQ4yqRjai0tub1KlV4oP+TTqtYCJRklj79F2KX5KV6NBoJIkofRV3Gxfj9FTBrQK
jTSeEI/9DSQdv9aWQy+V2WZr2yUzzX1Bxb7zKXhFOJPU0sC3rU1bLWeTg34BfyiSB0pEKUCpFypU
+qgMMBOxEqEju7Lh284BvN4p1QVG6BuaBDNS4wdxramVGZgmNnB1ocJKVjTVulFo/KBUKc45IAOi
wIOJULzgdIVq0UTZJE3viEhoT94Udy5MLAuAVW0tIQpKj5m2pPLsqKHYw7qafd41qVpBU+302CU4
FsfI+IN9ov1gvN0LQjVTFYyPwfvQzrfW9kAmE+6zXoOmjFzb2nkNpbTF9b+2NF7hEiYFhC3/g+oA
YrkVKiNU4zUPTyDHEg2YEA0jdl0tscP1TKlD1PRjYKw5NY5O04rHtnLSxJuuv0onACR6fJhRvfm7
7T8/5JiNpVsBagVyOtmRWqwqFHb8Ap7PUA6ekg0WgQ9CCeL5fVgO/kR585Uj22d7fw0VIrjskGTD
h4IhrqBebbQ0ZIu5abmOytbrsTdHl+7crmNxxH6EHpZGnVLf/7BtLMM+Zyt/hxDRSrnoHNIw52TG
GTJ/ylCuTItrNvxPigVtdd/zLTkkOPA6YHY7JJ4ofTiiD6/I1yqDCyQutr5apjxdc4AXyeRt1bOC
6Tla9mw54xo5HMdYsjDsZ0xhInQKtIKqd9IssP6ucQ/RgcJYeGcZ7LbIkomxUhks8dp+e4htCYdv
u8Pw8AjRmpZsbU1wm8b6BKiPVBkFJA3mxlTIFwjeaujBCeAqaUbXQEf8uk2RDQPUCTWyTbgR1lvo
NqwvwKBJuROn7XO7a4NuwG2txn3xl5zSw6IIhv75qczHGUZFDOOM05x++en5Zksdh7H6OssnmH9p
WxIRuHoyAG8m5kyT2XvERkzIjoqHtHUFsk/VNfCfjuurpT9NjoVCjhUAW796u4mnuPNH+b2UvKKT
H10PSsjw7WtAFYGZvn6KBLyaZ4X+nsVAYORGOKhBfWMJ8sfNe/jUv6R2XgqZRyTkp/pt5qjKaLNc
Soin98eu6x2R+wzvwylf26Pcl8Sj8buRlqMbl5XK3RQWWnRR5DMCDhcUU0aIjX2lXIuw05f3JBMt
b0iOEKiav+TsTi7nstRH3w+L/8QgvJ1evsVGyZ6Rj52hXksVoehLZb9SwbqILGoIM8/YfqY+tocU
23Nz5Itt/rycyjEHObYo0N71GgkSquxcQioVBquRbK2hKmDX1ZtIlw4kbcYGGexsOQoFX7aPhQI9
LKu5JgGjC0BSzwC6Kcob27IYSrwfUYrIrS4nn8VoOIRGdbwXBndb/6AlWtY0uk29BI3JQL6mqjhy
VYceCk9/WyiMwMMzAe6lrPgzGW+k01d9Q/Jd/NcXvlbL1Hv9rEolT4QK4uw3FWnzOYzQZTkk4U6X
D2aCS14/7ZioaewebumY49Y8UskY4H+bY+HTncA7ndKmNsJn48XwSxvElDHIYQf/A2vPtMNOIXBP
6VsME0aS4emdVrwJXf12/LrUvSxri2P1s06mIoCuyXLDUtwURig0DnLsHU1GdyI74v2Khi8bH+Mw
KxOwuxzPhBgUZyrbJ2QkSwXE+OtbXARnME4SDiJCRi4L6wm6X8z3o4EIRr7RnjwdlWd+oSn5JkcE
HLq0USrdJO8pby34GPDMMVIEHARQsyjGOaorIaYx7Qd/jsVRwehjTTs/Zs12J3BqscY4aMj6eG82
dkYDQER43DLywsLtj/XjZa6BTJdq5sgrlrbr1PnXGoogzmUdvIG0hHvqQOTM+pn2xivRN+Uc7Nvs
3OBXXF3aoIfIi23ZCMezllN3IUxsDggyyTryTU4IROy+83LoYMED60yN6xiGK21XzInKdzpf+f90
tXlhRxO6bCySkaB9GHBH14IwhzVyca0tTg44IfpvHzsaGU6w3Vz+WYT4aL3/q7Vz6Pnw7b9a0jVb
o5aSS3OcZhYESm5pw7gXKzQZnQAnZrbROQcnGKd+R3rxlAi+Ys2gpkK3fkeDudKX9WNcUR5zRR9i
Zl50YQGj6bod99jEttW843mvk4zNVldVfR0QnR6slvPtn8Jq4fPDMJrd8OF+nNgTo7lJOLOi69sh
ATd1D75t4LiEgHgFZTq738WI25Q6spdyPx29WxSDBAo5NHB1T0oCsnzwRCwTSlzvuy21WgO8tYor
yaEPMjXJ2eZQBJdjq4AXdP3YluA4tw4XpKlfMbpl94Yk2vC79t6vxTqeXzRsCi+gEJ5y0MAkjuvC
Mvcs1ZRaQM/KQ9VjKfLQlMgen68GXC3J4Fd++F1I848/SaZPQ3UtTSnFcx4ebEe6h4Hk8bvLzX0D
BzbRfPGoqVWcLfYniPoeD0MUMduOkZZs0AfkjXF4/Ybvs7sB0+kxdm1cegH7Oz8ETO6c6kVBaww/
Lk87Xw+88Mq/Wd4guVoCKYCHg+ssPGBBNAAvbW9h48og4vRrWTiF8ww8dkedOZmGmeMVzZb5rl7W
dZu/ORPcaItNOhFMBz9vcMH5nKy85WAvzhaZIZKecfBn/QHYaP7O6+kcptglyynj3CAD8yoSJ27e
CPb/NemGbbOj1zP2JNzfvpAA/Va40Tl3874vPw4OubCYjIRw0+LcvFthnsJoPf4THSyKv3oeyMEv
z0R3eRKngvgjO3sM0g+M20hk35Cc4/BPMmfBVgyttKsKiS6Gkrfkyu33FvqQlNuIKqQtU0YgtmF4
gm5EfECCokfrY88yBC5VRZSiFNqEFq1nzWVX63p3Htgz+B4sX9Wlwrh3uhj9ILai638gAaCsSwHW
YdjoJBWpYkQ8Jy+g+qjSf6UjTCf9EiYJTWveiN9wzdwUR+SYrk1sAeSQUCnfyDQ1i9JycIXX8JEL
oRaM+Drkk0igxLfcTsppk2SWlQq1RbVzyU0n2Gl1JNhQN2HRizzYnji5Eca8siEVwCqgudXhnPW7
30qN9TN9Wn6G6HRenA+uLu5MAJWE5tjYulRHHf71QpJRvnj4i5iyjMsAg6oJcvKy1KvI9MnmHbKi
FbGyYRmpsq9pK2hsd8SnqgTvKd2w48IMdSjciRLfivPZJrbGAVbuqiTZzDcEqytODoAD5HlOc+Js
2JbZu+AoP/QLSNdm+ufCUbXyohZjTsAvISU7RCmMAikDMtwJTT80DBEtECm5gUBl8Q4de6iP1KS8
vEDKXuZ0v66UNyd1L6EepnhcNUXwo+lh2IHtG0m2uDUHpHvQR6kepwQeJJ5xxyNIF0RqJRZfUO1u
F7Iide1j8erPAf7eFHzvYTV6gXKT9rFGYhD2UbN48eIRjzIDRVaEKvuZChDce+Xq7X3an583Ym4J
IdKco/pSMgH6xlmj0qXdqNLzUxsD/xk4o33ZQPcPPVdPNp9nETziAu2+XFrF79+MgiIWyb0/gp0J
40PAMufQDbBTt+83RX52sE0in3fAWuZMl3zHXHeP+2DJIqWeJxwesXlqwozR6jpUtz+AfAPNcYr0
YkBjdTBa7dXXviRR0ypUY6RgDkIoTpjx84+QGUJSsEZR3LX9BbTl6khISRggJdcCF557dFvFM8DU
eoMBD8mpzVurYmfZ1QWy8AEEdhhXF8lMY4qCFIXoXklDa8BDLqkq7TNBeNEdi08YJQocZWYr0Xat
/vk0lmoPamC3qdQ6pgjjsS6+rYJAGYnmRlpH8chC6xrdUKiUQFtMArEqpeyRoHCJ6wgvPQmy6e4a
yI/s5BrQOTqFuM0opmJV/uErnXmYPTkct+ZklaLZqlaFdHKkY5r3hCZ4lzsvIhWmb7Z+XrgQI6hL
lBUW6iuHtZEraus4v/ucCbWgqu0+6n27lpU8cdPmSDFxxPVoLaMqPaNASVKFIx8xbW5e961YKgxc
ZdghxPKRXzC9b0qt7/hpzM3ul5SRjCnlCokIqsx2ea/rT5eHGGEuZdbyX67J0lRVM3F5UpibNsWj
IRHnmVxPYShP80IJEeBAb+GpW6X12hh0r5VRJzuhFOTfJ+60hwqdQzDPuuxnpTIOoqaGS5Jf7BXR
Q8jgkfNJ6+Oh8z9iOi2djYwSG6dmHJPIaCCp4S/BFCLq4wdvakUomyhH/S9TloCuwbZDzpIuUJrV
Th/bGgX+Ia41kam4M/N4R9p4bXR99gWExXIPEoeUUH+BFobajTZPIaGg39cA6RZ26RlwefV/Zd21
Vhj9akr9yf1BA+W1L42bHZ8f6JyJYGFe4c51ox7om6C+H5UV26OTeHLh6aypQNFxiN7HfuFqaQmk
G0aVjgp+GDvPbfKxx3ocMQ7ZdWrsm1YgKXAxPfFILgix5Nmx3nu4ipjrF3SfsyZ4oF4vtpXSKTqw
LMyHALThzao6se4q5Fboka5Fon6t7O4I8PirTaIz+SM6qVq1vE9udPz0QVq0bLINuOuZ2JfT3711
usLbtpTOVS8VqUmTuEgzctj0Xa9A8U3A5vocYIcrNq8e3B2t532A9nZeALqqZyL06Lvl86lb9QQx
FuxwFl3SRBmZfWmgZfbIcqVWwINV2dETpwArxiGiKQBEla213OHlfYsE4wzO57vfBXLQKtgzKJh3
0UGHHG1cM+H4n+EKb55KCEIqvEIz/agw0VdRjTHrg/9MbW45j0fNqNuEPXgSDxRwMIru3cF4uElo
uAauMC/hZ8l++dvzQWxACQDmVKmbmGpzECDIzMXxg/+jQBKrKPfKnzNYSgpyv/qnpng0bHqps4Pk
oeBedUEsFb4MMVtPj3SKMUa28tmcp3+ZRDF+IntZ7XIH86mtxJWeHSTrhSOgq2lOxvL379IbveHg
TKi2hElAM/zv9kVEak0b3oG2OUWDsEJ7T9hiFiquTkQPmgXy6LJqA5CiXgCmqaamtadFwkZIX51l
ZR0215jyoyfxJKr+T4XBnrBHhO1ZoaM2+dpC9SfE1I0nHsHW8HQDZFnNaEhYRMmcI0XjS9bBgzJQ
ZNXPELGqQQKyfHNYhf8kbg+7SYJSkvzzNvtxWslssJaiyXg0pZh3DtiqsguNewH+N38UH1w3QIdz
YJe68KqEIa5LDixa2Jl7KQDyZmsUrwwQ7Ty/tYD5Q4ywRSvNkSEl08dRcH9vud2+tYXw3fXow15N
JREs1gUOPPOLI8ijD+RHKkLRSUhkxkxec1w454rIU8Mq2VZ5rgIRQyeqTHhNLFpD6qR3qvBKHCe4
PeYcUW8YxLH1Hus8iYV/g4tkoC+OYBjjh/qYyfVSu5u5uYdgh5qHWmOUJONMhKWQ2SklI6XYsi7L
UnEVEzbSmw1PejrS5WmlFhieUOvGcgLBOgm9ZIr1jBLTuZCDrMDUExG10d5ZXtQAzp0xFQehxXW3
vzXhbN9GtyiYeDuFpwpeJo4rN17nuyHK6yH0+w1DbUsZfKeul7KRKBjajtJnDQYzcjcAhg45kUlt
6ffmtoj4E8xWq3I/qThzVhPOhrlDvyuh+RR11n0ATogYbcvuzralNmm5poFl30CVyXEoeXtiuU6L
4YoHZe4ni8+OCsVyrrduwYOv/IWWkDK/iPB5aGMueuGjZpNT3/YKYn2dvOiuhNBkY3LdSVxdMJvS
7BLzGC84xv1jnVXX6Ti+09TG/dAyNK6iyhtZVnYa2fmuVO+xoy7HaxiRu+KG5WEtZYFBzztlj9M1
DcD0/I2eE6hWg9koVsmgUenDHfuquZV06k6/ObAabHrM4KLEKZ7CZ0jlzGH1F4FVX4IGomRz/pK6
WSyCxA5ZAwE/qG//wbSJ93iV346ONsiaDpnxgeuy3GKlUL6IpaQ+Bxw8r03kmduPsGuqc/eI9Jjv
7uj2nZ558Q8AJdElNav8wZbrObsqs0VhevvWlAcjKjdumrZClS6HSadAOL9VqMHDRo0ksMJKgq6K
2REAHAFdTV+KW1SlQoFpQOcFljQZjooAjXunHnBqH9l8qbwfC2xuL1c0YDCFoIC5CdOawQZrE1Uo
Ta9hRX9XtG52USl/AEr/JacgwA40pvursLYdMpjPDEC3GU5GaQBWPll21x8O9ddyOaN3czfoiJaH
jglOGWEFRNneDYflU1ctDgfGOLq99b2QLiifp2c6Tqjg+Pf5DwcQP3UmxpmLxfOotEF/MtqLfl0v
ckPzqr2mz0LcJbgiGV5QyQg9mLPddMmUiDdochD+R2hoRiTGVbpNnoyp7tukaqhXoUF5knuICUO9
/U28UaLZ53okQBsYVFk83gA1JGJ+q9ahR8C6DZxG12SHWREKVinZhq1vcWsXbhsFoWeDET+bRIq4
soaUfTX+JrXaxCnJ0rCSh7bDf57brq8EOqhUIuIoSNI88eFEmTXz2Y6db2Jjy/9iC2scCs7U70f1
DHYyFLqNe9/MDQV5WiGeYTIwGZKIJq7vu55qQu8qZbVLM+20a6Cy18YKU6voQcMl3NWYU0n26iDZ
Gjc+ceOERU+mZh+AWlFwCU5QhSpT99RN+wkP5FkCnq6ii+8G7jztaMKCyDmEP4yJBB2N0X/xOIzI
eoc/Sri7vhjK7Slpoa/LqRiVn5pIsNeih2uE6rDLP/3yEfIpiAo1X8bnJK3ppA3KNcy22DIe+HuZ
2gXoXfIVENa3kFftHr2YxprLVonUfh7/RO+OsVqHDHzczBwphwPz2bpsQwG/z54vfk1ewymaDmD8
IZBzKOgmEH7FxCJR25efGtSOczxJq/5s2kjs4zSZVl80OK7J4AZOHgf/7LNKQr4RntDX+tn/8OBF
EwGwdY/ngzd/57k9wHIo9IOCIi1DSSMCrwwzLjiUhFnuCHWJvFfOtplrAbj/H3Rlm9FUPmASvGYd
w2DCMoirY/iPTokDMfU0cFc447nna91RRqwnnNGrGHoJ+/l7NDnETuKraU0/CDTQubvFOWIFVu4R
6HzjYZ/+iyrrRrqvKb+RRDHqZ6ofxP9ZmlS8fI5qTMAfg+bI6giV7SPhoEjaqoAJYuZVS2hoDMoV
dqAW65FdqC72x5CXYqhWWvUhDvG9ody/2xzjDW+BeWrsvA/7aQlutMuGAjb9ipAHvNR/eb0aSUzS
ura1+keLHlvfjP7qCKJlVa4MHbn12Qp1XpLeOiB5LaRMJ81Hh83U6IytheebnXToiiTKZc4s2emV
foFFSYCfOVUEf7lxVWRt1uwbWdgMCi23OyQ/dVjMxIIHIQa+tRGXqJx1Z0KExnRnTDtenyAsnHcU
Jqr6OlHfT5wtx6EYV8bCO7yiHO+MPWO1qIVejjsWRR7no3hKSbMtcMIidP2s/HOR+O9j3Hiy/iOE
5JrNqJY4AZD9qnKvcpaR5pGRkqP2bIfJTE9OEDrQfJaRqBsZKFNWnAfCjFGVq1Foc6vEf7Isg2hJ
9q2xWY+gmyf2Sw5lAVr3JYdP15r1cg/6zSX0KaucmOrV2MjjRDrBTzgxpm8cmAgt9FHQXIQ1NZKg
zIGm1VW8LabZ+MMlcxYnqSyksdxjD23G7zs0x1qNkig8KNPJ/9lKE/4IS3ChED9n7kAVDO/KTacT
79qU4pFK4GV1Emt0bGtQC/IyoYS+jXV4hR+9r86auF9gTpu/X31ZX4cF1kDbFeZWBzii8H2EO7Qd
/4IbTouzG3PF6PawkmOPhm0PPv7Z3UFwKTnoqF5M2OV7B8ALxu1+9KNXwc9AEv3vDxEv5kLXZT3Y
99q7bHZOZCaftM5+W4103gMHBv8O7mfI8kxiWYGwpSFll2B0yPrajnRutc4NOMgicV1IpfrRwXM9
xaEQ8X3fm9atTw1tVsjEVCxeUv46tPie8hKwu+X3738A2UvwZcINM8NO+4Es8V3csjjlShTgCqhB
XPpknR1S9Msb8v5T9iQG3QeODWHuSCdY4kKaDM51txuus2PwxbOcNFp2Y1VItA/OGmrzdjkwGor6
Hukqll1VT6+KlEPEqVj9bc4sSrrKjEjjAidxPrSoauPHoRw6UYahD3fncD/1ir8/RWsqihTofLQ3
/viONRqZgm4APGsE6KePBggkUug0z14+9uNmYBM10UbVC/VGa5LZo43nGmTWUxw2AtIugwXVrHB9
L05mEPL/NJ4RURnhFKcAbLSo5UYP3kgils8biWmQJMDWNRguFu+z3WUogOejMCV+GvFIL0Cgm2aI
yfdKcY1vVXvHXEUEIXMynmjWlocaV/5W0gw5F3cl2Tv9c70CfDP00BmdFHNjCnf9IfAa31ajFc3A
nT5XGcxonsTgHcMKOz6MxjTEWwg9ijE/I01AAeZaL5nYnC6eZ3FY+fk5qEofcpN33grnGUG1x5N0
gPJaF7BLkEU4h8OaECpIX7YnJ3hlaznlqTju/cr+wygKdaNq2w1aNo9++OxEYUt/EEXvETKCm2ui
IwiA84IcKsk8hl2uUzfkof4ppbM8uVEeteEjbSwjFQGQ6EVnHxQMsySHXQof3V66fINtj1NfKm+j
32PKXtGstaRStqzch8G8cdlnwYw4xwaj2Wa20LOWVkUiApUg/PaKpPqCZUduXcy2oqReDhRMt+v+
Ag+fkl7IlMIW4jbxBXCvyojNPEnZx5gMpeVA60o7ECeWmY/Kz2z8EvME2LoF4GLnjliHR6umRpYx
Yztylt5qONboYgdhlxxACSwxWdzQUnIy7s4tNNuVPM6Ygzq6Jzn4q/al98eTEyK2z3VJKgyapTci
UktcnLqlyvc3nHO8AKB8TB+Rw3o9Xhqre/DlcWUFJZHMUxkrXzNPthJLfWQiXY0ygs81V+LsabBX
FZN60dNje4RvR3Xk8KvnhdxP39KS9FOMTPafltJ17pZl87gCIt+aWJ8Fx5zSMvdZQUGcShz3leHe
6HrAX1XiY1o/BTfuPCKj/NuSaauq3a3oPTLeltbhC/fI3AHnuJuPHMi/6j3iWD6csPwgkvW1rbWZ
NofhuKgeN8kAUEan4NcAez75rgSsgjHHcj5QdgSPSJrtC0WrsSf3Q+T+ba1aauUUgvG/jf/iImYt
6sDzIQxvBmG8i1+ozK6NkQ3VXWCskzIzv3eFgFcp/6e4E2k25g/+KttzoakhP4MiV6R4U+k/qPve
YK/1f5Z2CzGc/7HYwSJcO/0aKbZS7bWQ02Q1ynJOt83+hSV4Fc4rlNF1g+8ZRckSKRnzGgXpYR35
ajy8d+maPBUqar4yJpq9Oe3t8wXR5JYtR3lmSbC8oWLdyDrdnkT3MIExhly4MIGpG56n99fkwsgP
quoEYO99wCj+IDw62OOTwfMPXLRK49jNP7Yh5fEkUjFfrGvTOzCikl5Kfjd9i226x9uSMwpm7oqp
d1aLFKSLyqJ3Uz+2b7f8TAvsvhbbrCStIA1nHcelsuGMr87hiM4QgE8fXECztmTKXD1ORShj5rQa
QPmF3zC+OCXgMJ1mhBIA8jEFBSsuD5FG2k/pqIclMjE6hC+d3NPd73KqeAJtphYN95dMkv5Jfupm
6yl85b7m098pfIsfhqw6N/21azn6RkAwxrHvoG7NMwgkmRbbDBX0OkZPQGC1ejgyggdA6Bpb8HmN
aFgFG9idSCpMaVAmwT0e8rj81ZP8ZA87O9+fn7odYt4Me4pS8HouTI9hcQhnnDteSYhpOGm7FgYB
aW33y9DKnim5hY3GQBBbN92O6rkTd2GM3LXeWtREH1a4RBnAThZp92Rff/kL9eGMBh35lgj7nM6M
dWD/Cfvn2z1ifnmYOcF7cS5dfdkDnEmiD1i64M4e4ftzvl+fHOnDbfDBPKYPH0aGGyJzl56Li1Vs
y9GLPVi+4BZgmXOeFL5c2YbqXJr+b3xjoNlE6c7Ux6ppDJGh12oDoCrdWG5DRetkCz1G84MG32v9
tTnU6t/xt+Q/r9SyiGm1D8c9oJ8vlfS/icWR3M/tTc9hf1GyZkkKeLrEQIz5yskVWZmDyMcrcQon
aPuQ0IOiJPKM8cLyZ0YiNaygp/TZkjDGHKG5hIWElDUqTiU2FqfdE/1yV1quv3gVPDwvubMokfbG
Lzxis0jk4R/6o17Kji1rufy6e5PDUuURoL6HXJcu4XP6+f5lM+FX2WpuiaFPmwKluPHujJuAkzmi
di/dLw59DLtJqgGZe4dgd+YwK5tdBOL64w0g/jeM1Gxct229W6ugIHbTUBDrbrLERRPHsYLVub4H
xtogYOPsvxgRQfCdiZShMSp++8XF56I5ImE0Q/NZ8EM4UOmmOh+ECASFVhbjvuFuqTOrGcZ3gxgR
sMcbcMCEdrQesrIxZV53CQZmIXAmFsJF31l45q8qeZQFV6a4C1YbhhBWlAFEFQcXt3f4UJZk6x95
sucU0f9HK8s6qrWTpYJYj0picpIOgexWg2x34Z3DYJ56afFS/WU+72aBzcFM/+enQJfB1scY26QY
9G4tLFoW3M5uYW6cEGYMFPDRnUwz7K1XwjJ7cDsPdIaGrK7EYmcxGRM6O8DtamuOwHXatooNNMk/
yJidKuHtDWz2h5ll0v7cr5JuP474/E4igotmHbYhegwCuU5CNc8eTnzE8XCvZA0exfG4Ea0RrniF
ttkFe0UWJeYkIfsCb3XuV/VtIEBtiQ5cnhF2DGZDWdGszUVRZrGMqz2kNIeDZr30zzdttBQD/JS8
WZhp+bopz+5NOT40EOG89/H7WsTS2JZY9u93tOUFZIKlbOyI8U67TewTXKIcgmPeZEdn+Lqq1Wq/
SPvpm0pY1gWWIh7sZZtg0/EthayPcQXTbGoag2Tc5JVg+EXrxld+kDyfTmnAJV0K+32D7+6ou1Qk
i8c7grAewHE2dlZs7lcPylIiyxskdV87OwBkx7BClKdxWyCoFTXt41J+vp5ynTQvhoy1O2D+GfNM
Mn+/zpvualdKygBPm1tm/ul/7vmWgUvZ4Dc0YNFli8jM4q5uEzONNIY0T1n13zVqE4M+h4Rui9aV
BZfPo7xclN9a9QigwDlb8j/AqPjhw/1/1QZonTpr8qwbNNCJ8Y68oVybU/jRQVIA5OMDo0hXdE1R
oSt2O2uK1OZOHzkTrjZFTf2oleXbMbwtWVqOLRSl2/CLjddBVkxZGR0G6fzDcOlAoAEoktSweruj
eancLdjpT7D8PfyxxXRKkmA9GbzTgp4w6bfw+jd0ZTYk0jZmATcBVGG3WV1rRR4mD6vR+pynBw0d
yo4ttg5PN0ROpYTZePMm268lCGrmY4eEpeA0xaloa7CL1fTq/BNW+wxbzQOtnl23axogxib+Y33n
rgdk1+XS7rob6TlPz9MUuDUO8F2X/nSf58xNVaqB5rQWYy5BRjods1fPX/apu9oFgtR0CLmTpXMA
4Lp26VlMXxeMigNNBifT3/eq8B/VDBHacWIfUvemud3HUEBt9Y9urmQoEP9epZiEGh0tI5t8u7a5
47qZup58Y5AnhaW6JjH1aeCd9eCp41WrgkFC5KFcvVbGY7sMxP2VdCOgpjW5lHzEgkSZRQR9/z5o
JEG2LN2jVrJIrja30y7070IZkkne2nWKfWHreJ8M1Q+II+EREImkIyf0y07bNcTUCs3MtV7ukAeQ
PFcMC5+Kw5IXxOYuB0SsDYi8yLohxZ3o16k40KXAh2175DG2Jpi71iqU3myQjPnGGGk31JDcFiq4
OSIWI0H4uSwN3f2X88M692vPl9nQdWsBiwbtUAGr4pVLEzFJZIVPgrL97gfxsqPPGiDzuimdZXzV
vrc3o24KykOxcqB2FAZmF1XaTI5hcf7CJh/aFIzy/KdGAPaMc6OL5ogpL2ZApVE+K9ey8/Yf+FNt
5pv0kFC+7OqES3GNxRWDEp556uRMWtrbE/UPPiaQGD12p7iE0PnyTNqUhTzK3OB/D34luXuCryjM
HO1EdXYpF+RJS1ex4I9Fsoh0FfkIhHkG68mXnJq8BqrMOaCgV2hJ9o4B1FH8B1da+g9C3C9gfEZS
N09ZvR6ewQofNfELev3YlYeX+rSLlIJwmbI8RH+Z/SEql7U4d5XOF8W+fu/DBXsszjDj8KqUj/m5
5hYr1qCZTM817YVcX1fCajXtpHlYLZ9E+O1HCSeL1iM/V17MtsBBNJxoJft45vejczSoEof01qWc
YPUIvUZtmI7r/8mQ50Ot32espN+EPYRl1h83APET912MEV3toMXhgI4gXFcb6NcoluomYBPwGxkr
XLPWEZrINxEdZJNUkPHEH8f6WujendwASMXVsHiZLUB9GJz6YJAoIgfd/J420o2XT5CAzkBA2cDI
2ZS0HqhZ7s3IsmpRQ6RYHjkbywvtVnCmF6Dy8gJO2DyDSeVglV7UazYh53ia0fp5jEDsZmI8U9l/
03hf//6Ezq39S2/gxBbgBMYoSVph7dZk//vWYAGM6UdH1F3BFYY/lW6KS2oRyyp3D+US7cEDmSfu
jlgIpampLBzghxc3qI4jbS7oqVaQ1SXRTNS+npz+u2ZqVbhRfygl2NXYtSuA/t3ubFJ3UxXZCkiu
tkqDtsKib3mCMcPfGDZwy/sR6tkRcCvPie4EZk2oee9iTn1J4ZMBcEz8kmZD4GVLgHqRN7Tqz/8X
mm6Gnbwr/j8qRjg1I2eiM/445tbQmCAzMntUAeww5h0Y59hkAUfvcCPql7qNxV17O5+/JZm6fs1j
OicBspYudjG+nSnaVGNxWFi/HF6ZtJV9+5KYOIxikfvHlyZqKdEeET6t63LyBPJMDA/y8jZfNzqA
D2q/3mrpbwAck+cR1m+1V2d3KxRPfowyxee3hFYW+GWwpn7If2tjgtKZNceHYUvt5FOO6xfk76IL
ZqHI0wUf4KPIRQ5USTdhzpIOHx8aiZBbqVzDF+P7NAYZsJgvcGB0Y61abp+DTHT2JTT2kadNbL7H
sVLAYlnBrc44B7hssLU+QgIoEkfXfli5oDp9UqPuj1Jzh3e3ALUPovQG3ZzGYGdp696BkU3evFXa
Mbwb+TocrUlQnWocun4Zrk1KBisyi74L0eLAQx/u7b/FMWNCSmubKUG8phu3JpYf+PC9utWBKDl0
U61lqFj2F/AHCWLZ/HVL4Gu56qU1WDhVdCTinhdnIwSynKcCkctE07yotWiVH+gAFpUON7SbIsCc
r8bDVbEqAKnoGo0twFAE6/DxNhCWKxDNrSF2szcSBkS3ihF15M40lqmyDUtUxDbdxFBM2jPfse8C
AAjj/mxV8y+H67+SorKdWAK13MYCLMT6PA323+9aMFmxgjMF8Tk7UMB4+hVE7MKt1MK4Wz+L4tCo
fVPKMxYeaRHM010HSjTeo2OB6RpqYpvYvDe4KTKdaZ1TF4/IPhkOIWnjMid+Nwpx6mqzuYA5fQVs
+8EANHEevRqLoTcVaKwYpeWnaLF1m13nGZiFmC61JmmGQThtSF8KnkyqCwrucUDel2xOhWVTZt3j
gQtDMmvM6kWdg3DAdSaC98JBaRmO1O9f7RLCdEovWCdVuJthrfdut5zt5EPDqqBKY+0kxiG2ITjI
OVa3q+McMTi+S3LV8I7Z4PBp9SFz7nkUX8Dgbc9pUf/VrP7JCNqKKLZpSjaoM/s8dw24DLwOsMxb
6rc6i8zu7589lqDEtp3hx2T1Z/JqL/R8x6LO536E0+15sVGD7mUJ45MHuErNZZkI9K6noVCPetTx
bFnsWBibMr8O1BSXQoaUdX1+L1rBYHnNppPY4344bMa8ByPJnlYPHODNjdEWQC4ApVDIikbnjjsT
zpD7tIWKFmaPKe5qsY0TBrZKFPd7oMCaI3d+ZokYMjh7pBGSnnB4YOnuAzZu+k71VOEHoCYo3YmC
AGvVg9FEHK0rzCbJ3Asu1SGQ6fCw58RgOxQbPWqnPyHkh8Dglx66C3K/N24tMu+IPaMvMNFWfprR
rcrj318urwmOEMnjPhKwRp7EDxjYxvCXLBcZUYzeXvoGDVlrMs3eBFZrqM32dLJu+RZr/ST2j7pu
SiK9BS5cpz/toZgCKIJtih61Rzedsvg5jNTVI1caU0CEdc4iUpnt681NJ65uN5Ln1OTRC8+FaiNZ
clx2rCK6ZlnGHVzGsAq0HvHebN0bRC491Di1FLO1QhNU0jAMwuqMGoseETpJwZRY2JQ/Mkyo5lfc
b8UuFO+q8OTdP7WFU0o3mK1eDEAb5pc0ubzFerimWQgTm7mcznDcWvPqc6g1lY0HjwaAhk95v5jL
N2R2L9MnHlDlDqQWH44FJnLOIgY1RUimGz5DtMvvyLS2Cy+zxR0oBjEv3E9Ydj4cvwXBAO8n28wa
CkDC0pjMA2F1VhfJ6JR8uw8HSnJymfa9E2uT2AacZ6yhBAP6vrDyoAg+Z5WispiD1cM0Gam6NG11
KE2yGA+lDa39AeORE63vMGBXhZZyJxZNNZY3cCIvK8KzFjLY2qv7V7ZxA6lF0whWXBerWLYgdc7L
iPkTnTiweRuGdBIh46jM7sG37mC7tjM+qCD9Onl1oMiObSEttBipZWenPP2wHG7RyL9dJFpHh29u
zx+wp5NR6E4A4QZA0IdD2SY7dT7vTPwQtgmqLqRkT6Uv0OM02mHq4W+y/ryYR3vj3DBOrTY8KTNN
ogBRN83k7+3gl8A5i2quMtOr4vODoTBTbuCpxuC8yScVYuGE9w6JUCZbCSBl6VOEzLTj1QFhOpii
bjAyNx22psIC5Grm7qkOxoXiLJQ914k4PtiwujLnwia+MQ2zvppcbWeen9Adc5DYRR8QRa7HnAj6
gUTnz1YmReKWOqlrPxelj4aw3LNpqV+jKOitoFK8Gw0EJlMO9tje7GTtI2SNML22T7/A0zXExDNT
tR+W64wXWLc5lTTwrgtdfXxjoQKTzYAlx8+X3BPo1R4BF0XeLoTeLn5IUFXVrSQpZkNg6mNYtuk9
2R4tq762dWsHn3zW+eIWQ9BXrOc+b57P6xbms2hdwJKd1AKlGF1nP7Pz+BqM6nPfr8U7QFgUGSDG
L4v3DHbon/vpIuHIM5QyNNOGXs3ApEL589k9bKl6Bmop1vwg8D+WyR1uxBeVtJNBzWJb1AorEJmv
tpkdCGBRMqHqWf5cjh2h31RWeRig1T9XskX9eeL/Mek2TzYZKfegoHhkf6orPG6uJPeWOtbhMKuQ
IATs+nt8i8pohw+AZqHFxz4hCBpOd3MGsXBRiq0OEwn3KHpPJDKXEDsE2M8JxFGOJWhw3HbBF01p
5ZS5Om8Nj7RqhxJt3CbDKPNcrRQSgG4AJkL481WlDxyWAxrG00sTwTuhFsXFJQyCil3w7wfvdl/C
Vf4/weohIXd9bHkWtLIfegC0IquNW+b2NywvqbW+qa8m4/lfr2f+QyPWOgUPmDS61pK0UxhBiQbg
yAcXdBVE0ZklwrKRc7wWX8D4q2/aHfQv+g1GrsMd62fSV6mJOT/RGqWR3nquJrX8GQ/nDGj40yiD
n+vBMtEdK109fgx/Dou9+XuGLlCxNm9WW2xcQDNH1Nw/xNVMm6e3UuKyRsey3oSc6mPQRsYY/MDl
C84bpddYu0GkF9Av7Ix+ViunpvVG9sBHgPuLEL3X539d9z+0IDXQw1O9vAiDEU37hVckNLZmpl2h
pATHgo9MCJrrc8fhUzItJ9X1iUSyUOUXEnpvoMftBjwoSxHx7eZnh+NMDYNzZWWuqUtbnuOFj0e4
2X4TUrSscDTwBwIRq5ZUYYawAdzYsNc3oJXgLnpAJ3C+mf2uYS0kAgOtPUICjmilJ4Tr31gEBZ3c
kbAvorsFRu0+3aPvtH01OQMcqYApPrVF3Y5gp9Vl/8FKH4R+kHH0uzdJnAhyZoicVQZnPuGRRAnX
qOK7W09cloos14gpemcCxgWORoUozyut7qrfwqhbToBVSGGbUytHItYKmlZ2xvn7Oqtcxq5L3yNG
1x5SYx/aFeGm+vnOHOUGUFNe+p+8rl+Yvuu784oCHdb5pJUQv5n8NK02+F3nzGTEDy/fQEacZ/Eg
JpektUQs/ExVTvM4+Ft5IClWWSQnI5jVg5rPYxVpCBT5dmkHuinIXuyid2ww/ZC/Syka5OGrgc9h
x7+cS+H016Wu1rMVVOIZUZ80haYJ+10ZVYbTGBC50kgBAbln88vG4oni6ibR/ruFiepmz5B2V7mg
PQHwyjGLHio5Q1a2KAsmHMkV1YTjVLfAfWeR1ec4Pv316JJXBHJraEmSyZ4jRwsg22ZcJticu364
tVZlphPfqO5AtAUHuayQdwbl3ZlU//h63FkzWPKdk/b+CtDIOW9FjIhd5I9K6LnZ+Aq6TtocQg3J
vcQZLoG/F7DSN5MPW4KQX8kQV7WJrTpk9eTCF6WGPtCgJlpR7aefOJZEpHlnOcjCdMCthKqT/u0v
9Ss480caWm4ZQ8DL/xn/GqvLu+W5K6HxxXvyrnUkjOvmJPu1YFk+yVLs7iVRBpKzIDsr3oBaPLcu
0iMtUHn09qJ+qfW8FfLIVksJEMtkWSRVXQmevICgd2HD7MGTn6lIsF2VnjQ7Y/khZBobpcL4Tb/u
ELe0AG/jwDGwktzLSTrNXRxQHS5B0JCsEsY9tXDx7yjtI9gqptHo4sEljeTLKfdtZ460Mbr39v/y
W5W+PmHOtiv1kPxgr+QK0Du+kChCDHrLTOkUZLxjIt1CKrFW9tLINB+bTyEMUbyOKo3cv4jJoMSU
RZ6n1eHOheUs0PRURQ9nqKZoOX/5AQ0DXeEomm0F48uAxUnI8ImheqvcvL+yGfZwjU0S3YZgEeJj
0nxYM0IlqYReg1ROlHd0aG5eVj1tvYY08SVdzP0hZKuBC6LdQRzJWw18swo/HGiL5DuOd3OnOvTd
E50xnIWWJ4/UrColMBAn6dXjFyQVOe2iIo6LpA6TV1cSQK4QMnx3A7srZH0wgBpkD7GZ55CEXJ55
sHSka8KUzGNrp28vR/ooXE5DTuxMqORQHOSTXKF/64//6wpoBrJtUgClDa36pf5x78MAbOizTCvX
msOfKh69aj82pKqenmR+FEqxDPMDlP07HtVEzItS+isylKppSkCcEdi1qRc3MMtcK9MWy4dTg72o
89ir3bSHjsTrW/HagLWbRU0MU6P9sDXnQ28aGhmxaQPxkSCsBzieQPVSKqBVjFuc00hc5chqhIl2
zwGUF4XC0tircZrM3Qeqy6jLSBq0WAyIlKyqsb49WvWZZeom2RHAxONzBd5GJ5t8dXzH9XGh32Fx
v2uQyTjpBODqHnQ/H0Xa9Er70r5mcVmLAyfxzU6srPZiG+mBOvqFIt84GY7DqbuLqvg4sYRbbIQV
ogEM7itqYqjDNfuME8wpUhPLFqmqQ9ev7J4Ktk+j/Cd/LFAJjQPtnhACqajZe/oABw7yvS6sLgxB
bhjqaLePFE3XfpaIiKjBrqBUR2vmn8g9FaG9BGLy+oQ5JYOIBc61INbvbLdm76uvJ9w81Vm1bVLl
mV6zSzSs9DojRTwiuVhwJX70sLVK5uM9tjWxEdcgzXH40ocdpxByRHBT+yheJvfCRwpwW3Qv6uWR
XQY/GCyyMLVI4lJEGochz3w0S3PTUn8Uk1QP/vUFKw7HehevqYgwYxvXOac60CLFcZILGBvmR+el
1BLFz9XV8e51qLvSVbpVkiwl0Ktbl0Zf7lQAB0nhyceyI8tnFBPq0i4lya+LERb/ccIEQgHdhWbm
z951k6pcmRMaKxNltyJ30XAAz+Istca+mkuCnfNrJMxKwJ4i2GqEPCBS2QbnUqsBGdgoXpbftDx2
8RSrxS388QrYDT43YA5f//DtCVVfGuwq96kuel9UcnxYzuNZQweKaUwpZixvR0JCwsim0hRC3vNa
r5MSJFsBvh21opqRJNB0l5gXaE4BnVzouyVgIG1P8kCOmkYb4g3e9IZva6wlVMPjO9Q6sfWlVj8J
/NIw+kwXjV7606kv6jBDx3j/649yxUH4XZc15ouAw+E+kyZ2x6A8Y2PCl1EsqpEUM7QqOERbzVyA
FUlszpXiGVJyo46SaVySO02tLrREIN/nRAJpRlycf0AAI45E6ZeEym5ZwAeroO2D4KP3Ul2WsCqA
Is1/TIt+lretXz6/3THkjtqnNL+tVPwoJOvCL8wkadArMKcyODJk0GreMEvh9A1eJSgeiG+JpMz8
aL9sjp1KDQC9ghQdJWDsZaSnZYoM0+LL2Z3+T+2EtSnlMsxQ6Fl9n2Luq+D3EexfV8ueaUTTjB26
yE8e5JH641Auoee8xGudEWMwMZ5LCO5FyR/a9uahOj8YEUwrRJIxiYBJNHCh1OwiQYtZOfCngq4G
I1Tij4MJDz2a5p2jc3MD/GLk1z2zfapqYzzHlWv/LKqH5zDDGH8QVjicznK9pvXF21IWw42eX8RW
AL2Otw3wmHLaSgp1MIX3kfglbOwCfZAdkUfJsPva+kwiLNeYJ/Wg3a3T0asp86hXQfIBRE0xit6t
Tp4MgrXHs/urRHUg8QXMWtUdyPg6zKkf6vehN65bYPK9h53YbOBlDUBKAbqw4zsVgtLKT/ex6khk
eOb0SaYSLNNuqsQ4kAuvFxxGb/Sw7r2Z4Zi9CdCpRidkfG22sZOBrdTm2lLMVXrJqQyLEntYyALS
cIuabiLp0MRZ2Musk0Ol3tKz230kTZTcU2ugDrtgEuvsquM4h+7vfkbQLSaN1E4AeQOnKKYHp6Mo
dkjV/p+5oY8xU0Ny7ASj8cCU/D/h9zvI6O5+nF0PyJwNxCmu0gXQ3yY7kMJpxmCQxNZ51oIB7cqm
rxZrvumrf0W8xVmlBIqtbOrLafHWo+cVDdKLJ5EDz71Xo8oFoMi25cMZ7Lq+0cnUwh/uC30/ySkR
ajX7W1/oVGnrmEOAyGzLdC/EXoqv7geZ22O2JPqdhGgjOX6K2eYgkWFEnph8M1opKrtG18HDQ0VE
tP43mFypShW1KtLbFm5gZP5KsorLDdo29iYVC11YJzyWDgWCzf+AIT4dDkltZJ46g0T5yzUiEz/F
DC8vJA/pvnf/9EYzWaFUre03GjQAa9bevbh+VkkKAjIXiahvRUdE9PiDjwxKmxmECYiCSzKEakNL
h/Tq+vHZQ01/MFkz/rdOWe6O06LNFhcSvG6XjRLtdQaLtviilVHDeXJplz5f0Hj3oHrf4AEfyVfj
n33N31La5AEFv9pVwIksCmwy57zFN5soWgogNytYm52jMtaXJywBGnc0Tgzu05uAXxIPMTkD6GHh
JcxLuvt0v/5z6/gbJAeNzaCOUaYJuv5nchh1YJ+rhw6QiAijwyXcvjhNp1xdn3SWW+eRJG5oTl+z
TOajYzMSH9A2HrAnp9N/ldBPdSLopeaL+xgug3wS66Uskk+Yy+B5gGXP2srrPOdAMX/EtGhlr5NJ
dlmXLWt4D8+YzjxRuqt74bz2ySc2Kodq/VSvhQk9dn+3Rg7ol3BXK38DmgIMCc2rwTzwW796p4o/
BVbB4zuAzPFozmCFlahPN7fzaj0PyQ91YfLbPhPxsKmwbBx1T1cOuHPKoOSbURbBJqiDyY4h4c/s
S80GRqX//Ua7hs88aswImUTJvMAjwRPv/bCMi+VsWVBgYGlkxFnNPbyra0f933z+E9WdK1YFE9sQ
601hlaSjqGkXhh6QjEWxQSHCM3oTt1rKB2bN1hFxomfRP4kZHVUZAUYf0LyCY00yeiJbPvRJh4/y
WnepCGD9maLSimyZh224DOvFYeNdlX/nWv48A+npaNciQUgVajKdnc07LAQZAriNFl28EwsjpYCP
Asl5rW8zMvUVqCtSbgdH5gnRr7It+LUXvLa0KMJTIwLP9RHxk8Hp2uJD05Pot2S+8v7nJk3EHrov
IpnFiP0I6MIvYiz+qPR7TBeZR0TsHrvbQe+mfWmuORhep8u8737kK9UaRT3AwYTVe91leqamGKSJ
v9fPOjKUcKiSh4FVl+ApPp0c+r9Ujm9runXDbkPzLXlHNjzVc4+z3v8Rb7oLN0dykBA2MYRwa+hk
0pEb78b1/s4FGwNpu9jZmj8HRd+OEUO63mBwXIcVHc1kh3K8DRDygdv9X4ENsOLDJMbNseMThOnx
C4vC5nQR+2Hh9Bx1/2UAfDTM6h2nCxR+rGch+xJctgq8tihsYg1giqs+ONkwun+88Yjfa1tA3bJg
dt0Xi14sRcMOgRTio/WkMhjNPN9LQ24epJCMjI0yuaSmtC1AEj0hakAfu/Oj9ezDMpEzYGTjq/+w
7VIcsCbexZtSM4tRCJzPP72ovd4D0glSPkNh1sLBeMYwxIPSqyRwYWlM3UlJ8YyoRGu9IiBv3w93
u1xLn3r8XT3gseAW+s/LpgZMdFJFD74stkEp9pbLMDYupZ7pL0JUUEEN6VjlQs3ShmNc268114LY
B239gxM5mlB4FTlScjZTjKuBilHuql7zYKy7bHr6MGG2iWe9L5KmneFQGdQqte5RxYjtJhD4OOrc
sal9OriiWzshTYUMbjbjgJlpFfGa6fxny+1XWtSuBvvVHEdjebi3FlJJi5Gkf/zORZ3pZq23n0DB
UPjClhxieJfB1WGjpvEI7FQqm4W9YLkrzYO8vP3N/6kJqoJ8pUgciibN44cX+qaQRn+k0kGU+41P
0ecojIqzPa5jsuGERip9S/BqbLIT/RrKAC72AdnZhGO9Cmnthep+Mo0rGQmUWoZ+ewthp7S0/Ub+
2Zms2IyEwUOUOzVpNSjgBknqT9VyUrcvGf7PT9ixNGzeRJKpMTvpYVJ8Z2dCjxcYEao+BX4OQ2r4
caHvYCPweQ7wopv5qsPb9QK10b3Dh8Pq1zWj/vNS51OUxgRlv25pmJnhfYnY00ysQEo3I0ZNn9hz
EQRCCCaGS2GUainB49+Jh4BCKE+tGA32RqlzkFooCQCvcyg4AkwWUGj6/nD793k72vz9ab0cWYO7
h9EIa+22F7Z03dgrShMdbDx0FRKsSo9LrxwD+YZP4d+4AUHxtizhhI7RcDc0dRVcYB+6NmkB5Oh6
WIYLGScPH1zrXTJZ9EsN8+yL54Z223FuakmRA2eFhI+h/AHXnTSTKUGCOjDpcNaI5mPwoJ0yZYpK
un/I4Wm3Y1n+MvSd81AQkqa3yq9J+dPmAcJjcI8Iufiz2zfSZ9VN4Q4C3+1U61xXXfWVaMyZn1tX
ggifHJyq/s8IKFNpIW0RB4ansVy64ULtUbtsmJN5icslmsS55recLkrTAO/tEkDZHxIZ90AaAQP6
IQ3OjXEu30h8tTNumjowHEAZrRj4bPjY8C6pPXhUT0wkMHPPMg3EEyMfQRhFop3bHzQqoRtu+nQQ
MinKbyDf4Rw85iTgRbpPvuzdMHfkdjidCrfao55MVhzpvmVnnibXU93M82mYKGF8sByfQ4bHp0Bs
bf/6I+HIp5IrjfrKWqOMdgYTDZSO80YuTjGIJc5KjgswbDKtlzDNdlxUup9su5zeDoOkVFnTTzob
ptLGSKWMzvUsgW7ZaE9aKNLaIyDAd1xebpPEm6hqN0MrAFacM8L44h6+NSqVxZWdNORY/qMz7utm
uEnAFNu98YLLm5kDDcrkr8OaWEk95/IU7SGGEjw+UBs1zcfmm9mU/PTECz4HEDj2fvkXzPzUKPFE
OFzWgPqH59zUm4elde5IWXppdpYhqobx9nHjnR6KvlxHHzpUr1ZI45U6kN0/IQmWTxYCYkUdS+GX
VWIWxLvySKosp/9D3C/SLBYQyrEm6UhX17JXWJ8/JGB/3gRwMy7wb3w1jFP5KGeXmE1nF25CZHjP
U3KD1mmm6QgvXUGDeMxmWcLOsVg9zOvF+ytcFfwqISwmz63ZxbeY4eBHz4+2mmqqCuZdqrqtsWt3
JkbJV/Hjdx3KqbphzZBbbfm+iI8NgMoR/xZGyU9YVCargB8Q+2XG9FotwKvEfSK/DfsU+dHVY7Hc
TTlbWvZH+tKM9id3N1bve3kr/iWYlHhPWsthkGjWLQGB0QcnXhFFirW9WDtc0V5SjhUJKZtxke10
xi7PBxKLV6akXjq6Ua53h6SyJw5qig6Ppk5hlCS4zEc34Dz6M7X+w67/uoTaHoIrtYNK6+I7ttNK
O4kDOU7cc/BZAX1HrwfsdtNhuGtv2Ua8fGdBCGQL1EWNu32HzGYPUMuK8gzFtiyhYXLII+2jOoMf
s1WRunwvb/y5N2YlkmuAPnMg3iTso+C6B4JfKjW0bZ+gAwCYMJHH9Xsx6J512AOIqLBSk36f3/gJ
oHrL2ieeIl9m/JbIxsKSehy6Xwx8EK8HpmMZBcUhZWY0OehzPMu8TYhAD/4kk1JqQVy0bPBL9t5w
C6RbuYYlIoTSxOjSQvEAxoPf8L/m7Jkq7YsaX7q41T1pE85cHwhhztj99uAM3sQzNYY1UCGjyiQC
rRt3vZ7SvG4Zor5BTf9cbFWS9QfLhVQ8epVcdcSfUhSk0bIjP4eNfuxVvFlbcpz0uaqdtg85BWyt
rw1JTJheIOmTmbWNkMjvnjO7YSPikt1YN4pAJwqiBcXoSd7fwpZ68NdYUr2grBanDezlYm+yBFR1
PiAFJHresJwjtkZmypbc4y2zpVyPg16NY2q1xbeZyS+shf/FgA/e6lXcNnoBiAYiYw+/Epd3e5oU
kua3tg9tpPrxP5Ozo+YvXOLlIRb2oLH6Svv+0eEJP9aCuaB1rjEqN8H6YE4h1ApqZdTmxbV1ivDD
CJ+xINFDKAsTtGsKagMl0+ZE63gLkjuaoMIFX5fMN2V9yNmL5MzST5+HmeABzjQpaQQbN3Jn3ms/
0ob/MdJN24BexWhhIT7AJNfX8Rq4YxluGJE9kJdIt7DzYPXxzjmBxVb4PMvJGq0gM4lI7HbeQNr3
E/I5fR+KyYDnnSSip4rKizeaiOoWYHYsS3QUCqkQyKibJo9vMxdDz1AxHd/ExQnb5HDj3RH81nRv
cC/jTQnWKk6DGQ7Y1c3HOSh5A8QTYPq0AHl9p7FBTkjTpo8K9Nkgpvmf5XvyUj2Mm2nqWOGNR/Nz
qMKlwYw7rmuwONIN8yJ7oN/CU4fNfmZmO1qaPF0NP6s0tQzOjB2ipK6tG5t+LSDtQ6DkfxIOfq/k
204fzINMug1RefwWtxWvSQbToMSe80jFINhpKLS5KSloUfowXsacPLcd9BV9KTp+wd3mAQ3p3nft
CF99azOxFheN+TL9522k0BnzxyKMobwUn087s4FAxAgPliMKKcXWO7Fvw+IOZN4/c/66lYhVYrd1
G/1D6NipzvPReXnRoM+WJmj8IrPekU2B+6oisSBk4GxWZr/wUs3I1wpbWm2fgg/lVl8PT7hWoWID
JAjv1aN/ekmctd/dq7racNk0IG6x7MBqGSO6sqnsLqnJO/Uycu10r4NhoO2jSDxEwqR06FK5R4PN
mDdFD7TLWdAmdPAvQSkv1w60sgIqY1zpiRNof/vqQ02xfddVffBwkd4k38dg4AXFKml1qv29HAKG
+cG9r3IBrWQvKsPuwS5cSejDgiw9a+CGclA+O/Lj+i6oIttv0omdeQamXF2yYV/3FLCW5P/eq6pn
0zj/4hwluPtzJ080Fq+VBJzN70mO/erluw3X4bK/5IYob3HC7lPZUkdEtpJm+vAr0JZhwae+aFKV
WOZgseLc181bksDoFEuG/BZBncSzURSU3yG6dYD4/F41kZI5mxJebmJszw1vJjKGOresEHj90z7x
ubxRSvD/xwDNa7WO4wKykWtre3hWTmviYq826Ab3rjpKb6bDXELxCRo38TXzA9MIrI1WRDtIZYM2
Qj0JDzOP4hFha2ZNSlTn7xAoXmQOYvxpCqyGb2pyOIa3RB8K4GNPUj/haUe0GhxOjfaoqjQP1SI4
ktIF0ibatfUV9HQGGkwWdF91pdg4gPuGN8Ifab/KPYu5nUuQsY8oXPebr41J66yuWzJ9PP7uEKN1
wedpZp12LYT4B2RssnuX1oIeLRQVm8b1Y38Cp10eOaxz7+OzZ5/5y8h1g4Y/kdWm/+Fa3O/2ymfC
/2CYH0NWlMWc8BEiGLKhnG9Rzj23G29+IGz0KSbx+94KlOiX0yimPQuCXiB2q5k6zMpujx4+hZUU
HfJiSBJPvKu18b/V0Lrw91TgbDebF2HZ+D8RswnRp+EP8sCsBcuEHqa0uV87GNwBpD8aeIcBSmoR
dh0/wrNjrbQxGs97XOodahWaWQS7IxM8gjsM2Vp08X8Cx/Rha8ngBb08Aw1XDvR7gI9+gB+Tepqv
BZ7B9EVDcsAHMpN2cZs/wLNkMyssgQQs+tkh2fwbI/o1XPHRjUcaGjEwK/mVf4YuvALnzaMMwG2b
gI93SqiO28BZyqiRA9clT56bdqwVzEebLyRDeWAZrny4UzP6VppMifj+ph7aY1z5mSk4T+m+skzA
Gb2tIiaeUy5G7pPY0KkPJi0pEvQnZaSqaIbff++pI0h2OyA3lmpt85Wxl0BwwU+emfhHPJeEPXyC
gJco44ik03OuhBNVem6HElBlaSgbLaaIH4TXztAHFIkRYXGKEAnlcO5iJEJfV3eRX/JMSp0TFkUi
SY3x44NRDH6Pr8N9Iti2YVU6hm+V5oKFBTCbF6Kv+LO5lO6aCrVr7T+0NwGhA5GuZyWFuDcNhEYD
+PtWN1NTn5MOiM64hXhFbz5kLeFDHRcIazYJ7GtqBrrIJ+r7l3ndyFef7rC6GxjolQmP7AXGMTB8
rBV1sCDefOonxC0B4C7E4uDIJc0HSc03WwQDTb09wrMyj7B0SdNNDbuMaebD1YuyhEcZOlIahU/B
Qeh1M5osxIbvRBnZS4tkHN+NHwS9pzJbR7wt90kb6aZ3minRlxNylGtXKaoTVfzDCxcvxeWFla8G
XEEmkNK+nNGJfAjitAShrtXxMWRjblPUV2ccRAlfnVOcoqoQstucoOo/R46Y+ryM+cc8KDiz9Mgc
J3wD3v+fk9TyqhP2UIXQel2nhdLW5JozCUGDLLrWc+NIE71qGS5o2WAiPZdoQixtEKX1yWnLJ9u0
xj8Gf8oIRSOZ5Jqqovx8PAZPrTcK9MOPpduB5bl4fQIgWD9igNHnBfOxM9oIdxehYXwgNQOIxXJZ
bWInjeS3czUPQ8Az8vYgi9hLqv1GFAEi8AwGCN4RZ0VlMZLLe/s+ERywrmNb7VWT+grFsUj5H8vP
E4lMpP86vB+Ar79ny5270vqRKONX7aktxcd7bapf8S4PWfFtqi+b9KxUuo3pcEQSK4wYGww/ZadY
QUSEmBs0IlFPtIvVO3xAijnd/ifhPYAbfB48gAYdR4qigXD8DViB8PpBT0pV4CXfwOrF91Gn37Bb
hYeRB1EpUICqOS0q/aMotxXm9YwxTXD5ziJx0nvb/wFMx+qO9h1CWWPsWOZb0k0x9IponXsa9bVg
XAr4HtSNOAwT2YOB67xx6LW0j9/B+WyMX91pV1EICeHus3eXPAUJBAERjJ82am4r9+PgKv3DZmd/
eRVGPbE6uEnoKef5MUNoEB7c8gj+/Jv6Kleqp8GZIs3ddl2Iubz68z2JbGh617LJIPeUXppMIxJ/
HmkFLHQgGsMWl3pAe3rJDovFwS3R5aHB2vmawdlsUchCatMAXfVj851eVuy5D3RQ1QRFDk+ElzwH
PLEvq7Z/2sObUM+secOhrQjAnnnEd8WZmsRezJqsjcJ4Q6HoqtE2dEbv78To9il3hvUZ+PnyXFzl
cZy1yRBcdTI7RaOkxb1Y+4mOVPJkyqfYEkHJPxHjyCFPWB+ZErVlPJOsKFMtW7X/Qozt4dmr1uLq
g/UBfIue1ZSO2W0+jKD7z/OQOmu10US6qUv+Lj/pN+N9YblIpIuzOXcDtePnu39qUZlOx2yU6yUf
ELCg3vsZQuS1yzTqZQMNqmN6OLgc9kqN5WN81i37NyIun4zM6dp7Sm5GLg1mmwoAcUg/J6QGPHiR
eo00QG1T8ZMTg/io21TbIrpOAl8zq9h/vyRqtq7OWUp+9yc6s8jNmvGju+o0x/Z3FAyPGDHBmXcA
oHE/mj5neXYPgHcdemBswxgHtuOSnUxXOVRe1kNPvAY5pJdbnYH9dNM98oLU3EnhevnwWdJlvVqN
HRXm+mcjxmb4wPah1kqnc5iFRYqKUTPVsIw5xzlo3NA7m+gyIErlUW42Ls2SbP3vVLrDKgCZUJ1s
1DJUWg6rXv+U6JbA6IZ17m9/n8b5s2puGq/oJX+BrrUJVF4AtQBXminTaubuKMTPLUsOcsoXXcNf
1yjeKWeWcJsiTqunMAnK4GAzMAwwe51LCTA63LKTHOBDBynk3VdnSRPsRcmKSk5zYRHb+fsbwoTx
EoENt/WUnvmBQV7zZzUKGpeVWzRr1PGHmK2NXKvPOkPnURhVsYVklSxM7Lf2Wyxs5ZUYDbFnp8Rt
H26hGrMlezNW/WGD7YYYhniQg4xIe/nj0RdPdJskqUjV5D9f7vzTCrufmFLUFNekVm9jDwpsTxXt
knX7aqBksL7Aa6tlWtiHe8YNUJJOor6TVK4mtxLDoPuUb7xFBg4Ntz2bOvKJrCzlZ/q+SS/j2tjv
Wg9igQ5Jw8Lpm3f2lFp/6kmy8TuQZYxLzmaj7BsJKt2dG1qN9+c4gIUbBd952KNo6nhTo2Dhi7BK
+cwYewpDznWS+e1GguYDjtSMma6Mv/LaPO90Tv1wT//EPRxQBgt917NF91gUNY4RIY1RxDUu/6yU
naSUD1eJVDEuRCF3Y+uC+MuceJBjWQ+Y6GCphfqrR6KRAdvx5URmJ+twLDBREnHdObgdU6ofQDO8
wnYmbJlBGRZ6MdKnN3fQuqdLREyCFFTbkPaOOuIqSHy5PZf0Cvks+xXxCBfDnkMNrRk14JdoYs4o
RxeHgXIFXwP0DkGERYpAfnHhUEH+x3Z3958nlypCDJ3asbnfMw3HfKy/1PGE3Sha5R/+Q5D3ycxo
OG4PM5Eyh7jKUkFjbqvFsd2jqfL1RBB0UKVe8JAkZdJobLw1fLSoKNTb8eQpJ1MjSipN6yOdEe0t
Z9wL4v6XW5weiAJ2sX+BM3XZ4Op9NwnIIy0v+YoS1CZsHe4MS/pSvV+8FRqQgtHjZ90bRbS4kPKE
tTNZexwS6LKUR/w6w5eIoNPbaBR2tUSZ2zAEgaxAjrnClPdgch+Uq0jgvQIv6FCZ/5cgobk7GLgr
wZX9sysPv4xxDxooSR/duxvIFkzSUVJk6DKH24qh6hGKmHidD46LVLUfYfEW3Q3UVMy/YYd/LC9L
UaNDHVAlwMKaWYjdkDKDRc+jl+DWlqnb/ndQ8eS0lTBaW0gZKJacRWtZzbwdEo8ulCHR10qGMyPL
gfvmHUBLteF3BrZXeBuVnxX/FwOaUqvNpwr2xPL5R6pYtu9uyJmMTfFT5v4eiaym5W7UIGf4qbdP
7JCLkw1oC2qCtCDdkt4qvo1T2HwmhlrqIXE+/7tJi32Taz9dfcXKRRLjuwcacej50tI19JclvVbO
aEyQ9l4nzcSxgako1l/x9dcEABorEYxzPXW5sn2LhoAaJI2JLMCGoY3sUyTMJxuUOSvmTTfmqHEO
mQ8STWLs9bPBpAC40fKhhtT1chGkbquDX1EOECBbztmLJsgKs0AGq7HlhyLmOAu8xpvK4ayldOVF
SN6Vmp26HWkLJMsiFkCAwgeJqGIiHGDXbe3x+paD4wXni2QDBaVUarsVKW1hmMgCdVRiMB4535d6
Dt9mNl+u9BKpXNPd4ASzo39h+ExJXBTWBStXz4Tj7wgySvnXA//qM45rTpup86eivu2wpcuqbZQt
B7/Ft4ke4o08gvb5ie9e6s35ndG2MUKyxNRGOGRPER/9uwPbmRFlzFvUfTFjd1AGdrmGt21oC6Tt
TwQUDC/LhvnOeke2qTiVhfZRXuwEkK3h3QOkh6Bfo/KxoGG27dxVNigBUyLe/JyWSMNN7r6tXQ8X
rlR4S6iDdcsliIlGDppDscptA/x07U+wAKSU9ALDpn1TyFOqIXq/c+cIJbB0G8gi6AWTo2plLwgp
b9VAcpfv/X+KAJhsVWXvJZ4+ME31eA6BwQPNnpQJ6R8vUij/9N2Q+uELfhyO7rFBVBtqeybKSF2W
pYq81UH1icrYf0VOKGDVBsU8d4R8G4Rmi0QmSG36Xo14hQnHQ7qWuzRKrCDIAjrzFRU0h5DpCAYL
p6Qt5wVMrlL047PWtli8gwqhs9jJIu9R2S0WTHHDeAgKaABfUQQijQosbpnnRqIpdGCAYwyrFPXD
EcfHEf8F4x9iEH/RL7f2i4wTPz/8dKKl2PCG4S9sQ0Pzc2yFdIw9qBmL66DsTY8EeRF0Js1mCtAQ
OvMhOh1yEOHobB/kcLZyJVti6O3z4vlfEJnfAu+Y3DK1VuneR71inC4yhafN1t3kcC85FBGIxjws
xSS/Pd9YVsVl2bkr0OZb9UeAffRdLNauxkCImkS0i1+WSDCj2fF8N99M84VLJMqw6gQSKGv5Vwet
W42MznxFRMTU3d3N7O6rGmFkrdbIsA7mrKR9RoOx9pYU81Vuqk3JDYqwP3Jej7e4zHU1tpbXwhf6
uaE9A1JHcbFMA6Hbkuw6EFsek7nD1uPNobU5LkZE8xd3PWa0IaezkYKdiLpBeEN9T37d6+0eS0gr
AuCUrJSItQQtIZa8bxapwJQvYGQTi4GqPbt8QTXRbghzCfjLHim4VNL23Kbbs8ba0u6Hj2+QLl5Y
1z1815i4Cb1lZUeKe35Cjg0S6iOOWAGXLQzusoCERgVAiCvRHTV+inkyeAg7ydLsydAQIInXQpc1
caM5hJTAHH9dXf7zWa1lDyekNgen5LOCCrqC4l+gJM16hfRTE7vd76suqTmSF0EBSyPBvjRCFP5d
v3/6g/gn4M01B1sd+QZJ3iLKqrzI//if5i1y4cmEbJ0yIC039Qrdn9sfsPO2g9r6g7FtHM/b+M3h
ePfkybyajmOCbb2v7cZAY/AsYczHTZLoPYUjj4YAHHXY/3HxOvdr/vsHk6aEqqZFffDu2go8dth/
VTbSXryJ4dPmm5GXxOfrJQuPGti2TQKh3UwT8te1+rfPPm3KlJxKF/EQmm+hN/hjo7PeLR+Pivwj
QXFNz07xSM3vgtzEBxoWgX9pXLDh6GSFkjvxbxQroAgUZz/xU6Z79z1RIfYePbzsQnMrZj7DM1Ot
0KCSQmB2E2fkXQrHDZCs/EZNSu3Mms2W6mHykaidTLwYrsmjEBQVtsFo+Komqy+9q9LGXb1RZ4og
MEKZo8R3c80DcZbnZXNjQrGEUfc80trILitu8MkzGjIGSF9Lwf4JwrK5Yj7UOtKRXP/26IbIdeJ/
WLjevNlUM1w/sRvvB5eAW94/zE64xJJgZzGFfvy4U464ksoz55bLXL6ntfn25dyXFUovPtGXKSpY
C3kuro9SzUVHWRiHFmNWivVDMCTNWrtuAMoyM2ZPbLNmLf8mSs9nN1jghgGdSU2fNeh5d9ZFkMvx
G+7ukK8K4msHobl6Am7R8RU11Mno79Mea1bquCO4LKIdNJWvykDSmNPITVa1AErACYRTQzDjqPJC
sRzfbvABBr3+72MR9PbeTi7q0KUF3zsxMzEwyOjmZAfKQ/wB45YwKs37v9U5Eq/09g1GIcEgIxO4
BZSexmBCaL+Navle0j6TKUuVgx4tCNnUIpptjMl+d9z6fKzvwTm/5novcerptLE47abb4+JcWwh/
zCk2GTBCN28MZO8sZHW1xNQAWIIWuiIo8omHKgkJFr1teU6Vh4VJkAW7CfS56u4KfWTTkODADvLX
lKS6RvCbxAM2P4UEw2nX4pt8TPpwmzo74CAfqiBPaZDZxLU2hGYeRtEBMbV1WkywWthPyKV+vR6U
MSDGjFaJLWDgGNmP2SZE2lCHkIr7oF5QicxONJmEgb7Y3fINqBGQQMoaia27GFMEpf4HapE1BvFN
zYFpLnZof6g2bdiUYMEpwHHjtppKqU9ujWRHzJ5e03aOyrHv4WGjzpdmgLteIOwmMFXNKhIxBIK8
CqBZHlDC2aJsa6ylA+dRQ8owzR2mdetoF5anQhLNUREVGL/5RcskjJGI4XZdLZxNHEQl+wNSpIM2
Qft+BnO9ARTDswm5QU90wJ5yUNupcQWGmzvrXPYD6aMiPg2iPPK9nUiKStra0ZKfF4O/1AVl5OI2
I/y872221cIH4+ZZj0gqFWdIqR7/2GSqXZHliYAthiZD9lNGpRkZjx19T1+VjMM36ih37VdIHtmM
/Na7cJGWD9lMJIoc/FkCQkkClwcP7tC6NFRAAyZ4iUFD3mXGp5sFy3O3qdcDEER2HfLdsQEMatRb
8X7kyMWdv2+rwMaSBMuKx8MMq/GKWHdm2jd3pxrvoPww/Y6IMLXVPaCO52A7++6CJQqZn98DBdvf
tO1ftLspV/0gFbVuuPvl47JmKP/HZwTc+21Lq6GcrcNU8SFuRivtEa/HxFuLORmYeqEjiumjIi4Z
MkpeZBDolFxuqaK7kX1aOQfb/BTh8uUoNZ1dGGe1QSRCbCAxM8lerNwtvZtd+6o8utQImKaF5YMf
FHS2o8bZB+R9exVlP9ly4VnTxxSToFogbYbBfE21MgyqtrPhlCB6dKD86/L9xKMTMndSCW14+JOD
j8Jk6XpfDdgs1hOMkCz5XtHkBbf0oWRzZ5RE5XrcFqe76I7q+Bwf2FVGZ5OQuF6FoxwcLzfNtFbI
l4J83NT/5Z79V1cKUA/HHw6Cis5XEpt/Nv97cEpeZ8VDV4jG5vP7PN0/nH2uqis1Ia1uJNUWBqfx
SPdcnpMXlc3qMVb2/c6LdGaR4Mlv9pzULY3of4wBAVydviiNblzNLHJZK9s2YQUSlLlg1itnHjck
ojRSqdMEPs/4Yd9qsQr0WkEfL0y/79QhGfEGDhXspF6OvYICm8gTv0gv/c3eBsdJp+bE5JRWdM+b
8nsBZnz1g6bsRyOINE9VpYOVFs9sm6CT0rBmOYBJQcCed5J+HUjvUCVUZ39dUqihB1mrcbOesPGf
zanoU71EOz7NzBe4915vFflfxsGbDlMSO6rtN63yAkc4zR4qsImowN+eoeQVKf0z+yXwPVheDJeh
OKOaYY3wZ1NTmszp3jNQtrqYmPN5tZ9RJ9K+vLGCQcxezxPEpxD7qHfbVbYHAZBO9LJtaoAmjnTr
aAGbDHKo1sN1HVrGMGl0yAnMDBA4NWr2jb4O2U+NH+2uPzSv6JVmX8GiaWkA6x0T3A3vwuSCaCnG
8V7/sTdUvwzUFhvX+UjvB5k4t2gPEhYGfqLZuIOPqCAiiMiyYgN6xAJY23GZiAEMKymVT1GLyWID
L9UoT6TSSWYxwX4XH6rzDQNrAw+TR8QwOyHd3QYVp1qsy11KEmtKKVinwtkYWVIE6fO0XrttzOJR
MZgaQgzjQx9gKjkuhVEioFUQBtsjqQwdxtN2qs6e2SI837l4Qvefmz91rU4XQVBceGIfIN43Eob3
wzvfurrAG4Q8mieEM4DQug8t+z7oReJhuIJZMaycO63qupod8tZNnmo1qmC54M2hqpBVo6rTW2+6
LdUoZR8sQEO9gDzBwNzMzjtvH+6AaQyKLvTkEqUbANJKJrueLypZKXTBKIXmFpEu1jFFJUTesBLp
yQd62/60AA1kIXL+HqUoaICtZegLVJGNRmjHlwzaSdKrnRjZ8zlgPXPXCJZk/D0dKhRnB6xOmHZL
AR+ZAzzF4JcYsch7enzOYcxz3tD+ajqkXgEnuOxQ7vJUud16ztr7w5u+yYFJ2go3vPUAqw2SNcER
2yLy4f7prDxMfLrv6oVSJquZk5OMJDuGDL/NUuyhQgULQa+xHuIoQfaq6it3CKtBqbW+IwLRvAt5
kQzrf5J7+5Q059S5GH/AABOIzScwcyB1Frsr3CrII1ztazmkqCZurrRd652WsOQzaPEFb3pd01Sh
VwEMMd8HupZ1mqXFlOwlsU5Ii0GdVn9t4sg5JB8Tyl+KrA9bHHIIqZK/4sxFuUnSQSsf0QtX9wOx
hyavz46MmDuf3GlnqKxnCm2MmaJdQddEPi0K6BAe2CmaADMnyjHAdMiYHhrtGzb98UV5/jTJZgKY
uXWOdyczmsBklKFU6pgcZtcGcINQO23COZDJvomJpBXzsKFvddqdOvbvQvvlllLX/ihLfeMV48rH
O4AOoGV+LAx0DAfFv3n32CcWdo+TDuVQx+l0aQfo7SdelXP13NI3hjZf/jvdX49h6gSTJxCLg/bF
I7sWkEvAD2kiRpYaeOzw82oeP8HpN0BMqfpfP0ZZsBR4p71kz+0Jqrv5lJskz7DdyXTAJQFd2wPc
Jtr9wtHcb/sggga3F6UrTwjp+TxZ2NU3K1DdVUSlcvq1W1LILxoy3zdoFzwiBnhZA4p1YP2x0Ty/
saj1KXaZKna1dLJDRMLVUd6jCgnoKDCtjT3VUpHeu0TBgdKwAUtmp56jEihOG0qbhoOkyUVFtYBp
BdLirYRfziQDPgqZgv8OHIR6dLUbLI6EzJFCMjtUsVEBcB6kbk0YOLjTWY3yIb0E7bQbiaXLlRfW
9GqDl9CnwYQdnQGUPXDzbE0O3kWQTMeIzlNle6q5Dv49534AA8++e1UeGmkJXJP+6jn8A7CLe2ki
7dJs0kjfsV+GIS78wVLES6cMmNXt2qZxanf0p6MSsFG34SKHURxZv4ab5NCILTPnVJG5LeLLtTCL
xH4tst9ojC6Ve0Z+5YoyeCyCb6BT1Kzbs20NVd33JXwKKFoQgsHmaOcE+Ii+tckCMGlIssNNOkwk
h6PGfEkCscUKZrrei7yeemwq4Zid0a12bwwhS+FLkNlhFgg/McZcAMcxLGAJRflTga0h1ZhFr2JH
1pwYyaDt61sT8qWacDQ7U/gXlVKoKattK+cjiKvZ0fbcjIa4GHnAEbd4WmPWGY+EvfkDHfBlfi5k
1/1SYvnCEG3FkqTEQIx5vQRG1P4dkXYxu2H+pNCgvGsEgYvc8TKalqd2D6kmYz+mBsP8gF1ffNlk
FxLubOocmzAfmWVRSp3t7zyxWYwJTYmkc+785EsubhnQsHMnrGGcBSpS2VypePb1z7c9TnBoOkwj
CFGXuzpD6CbiCV4K0d+esnVLb6tUU0nmJmOyVwUgkSCSLiKaUf6Ev5N+s20RmfoGwSaxOssfJyRn
st6+QcsFPVaiUvZHtwuZXUESmRhel+ZnUJFAoxjm9jG7rP56/Vwgs674mY+zmXEON19Zgek0RC27
HJyGqNqFKGz8NqZoDkAbbmOGChs2wjSqNBQ8levkH+EGTsi6Qpe8JSipizR2tpxKzq76s360ZAuC
dWd2I5e7SqK2S+po8BrvStQeY2lR/06IWtWXysEIMDrSCb08i27NQfk30dRJF582yqSwEEvPyKgR
I331hCPhTg1TbPG6NraOo6oDQ2CHWEW6OMtHhpEIfXRVDqMZSlMuHMf8YcZQo+6S17eUSo1xmCVV
0Grk4Ci0OHCUY124ceZUKa9qYzETVvqRjFBYToLW9Prr4BLKBq9Z7veWqbjXDjD2n70mBYSQHqx4
GOzsP7YXwdfm9QqGeIfhEc1GHqE2Mbdi3OpD69xsal+cCgFbQ+i6GilijpnZnQPK6weiFzsgwi3e
KJPs5a1BR6aLv76RWIYcvtgu3BIvistczcShaCV4+fYV+uoNszA3jfIDAWgiJ7jwdNrgUOdCpy5b
jP+8WDqQL/30jdfF8gdyerPHdahh9FBgLyxt969OMtOzwV0vAxgiST5FwkFS+tbO4QRWCGpUtcws
+k3OPxUcR4ydiPRgjErdEJISscXJ3y2H2aOibuMcSRBU0C9mLMU0FGMPRcQFl5BltKprG8D8Ba9W
PN4Sxg6Yx35PX5PbCWbIoP7sLS+ba4NNy+kbt6S4HFRmbtHiIcMZciptYq+Ew65E1pGGI75Yia4l
jJs99febpOs7huRcHs1tK6B7i0dWjfkGBfclx05F7+KlvDeTG3XitwxbbJrjmUi36OhIN/XzE2Ql
eg+jMABu/I00/RKwO6TVKXNSfXG6P3qiKQ8vs3NyInGTMMiinBw96fiwumJgv95yGFVbHD5Yz0l2
eMS6S2VxGju8YShDIZJXOuXjNYNs1Re1h33D3xTCb+kb7PHj0MKDKPNmDiZpdXAojJe98XXsC4li
krei3jPMdRPcozfer1PE7HgKyzpMlPv2PtTHcVJQ5N6YF8fWQAxRmQqTgHaTXGUbQP4oCDJkzuMO
AcZg4yyZE4ruNtcBDYrXZ0NAXcfPXYH1hRw91oStYfMJ9gT1NxR8ELdcNwskUPqRsbHPpTSLibBv
IGYf0zeF8TBOPNbTVujxNkrgXMzA+7VBNpaaxi0UrXS1PSujyLrj7VMil1rqeRFKWCj5+vJA3lON
u5F/XzV+8YsaJ5+Z/SSW2xNmBZz1OlVFmkxo34C19hSohkrkk+m9+ACQ1ej5StuyVLvGV+n0jaxZ
uLnwtMLKaBYjZmH01sWEW8r2DSq0xMeMbXDRWuA2PMjeXblOkWhMiIiKWwbxEq/mCSI0XYSaq/r+
32lUPVmMi9FEtcYqkYzQ39vXltIZUCUWmyVVTbixcTuBp9Qo/3rU+c/K1pRnPHKMmTXmYZfQm3TV
GdxoTQFIWGXZQRinHg33AIqNEpgzRGZcY5PD8X8P21wrBGnd/jM0lwc7sGZfM+KLqtp/UxmZUMSy
C/KIW0YPOsJFDRESPUw7A6hhzgj08xVeSIb88xRkUBTr0HILHLRzaBUkwN7YW3zfuAo4zseDDbhK
9kDMDNUQaNNzIix1QlfEESX8vynkrz3QtGypWG9qmDb0dpDo2azviJ/JSh6Nk3ntgfJ+F+FlPZE7
HjbYEnV3/Sz3k/hVamPBmNnuxQjKOI/CMIX4qaC0WQmymd1ETZNH3no8wmRh0u0fLl7EbLFj1X02
O1ZCX798JqSJaIvBLdH/LNwKFM12e0Cx5XuD6h3jk2UaochZEeTofidlwQx6G0i8cqMUl+8eXTu4
mjACQkhyUFd52vIc5Y6jY9+f0u8XJCp4NMWW/7XLOADR0CkhuH8ZFQKx7f5+y9AD1daTSL9t3riG
KUOue7VK6SwSecAScE/TjWO0HLB1y8K1Zp5tV2WTiCSj1P1KiRBN7olWYSw0zSuI38ophP55afEJ
t8PVdS6CtFhA7qQ7DL1axx24DroxBYlNCsJ22wF+ScoYpkRZHASfnF8rjyUTpDoJ0DZxZreeDECB
398lXK3uLFD2yDUNUGnYQgHBLbGcglW8C3DLxqN6O4PdvYxmP7gs+DIDxifwDekSY0pVcsM/aeBE
311kUc6rB7JyTprrkCM8V4G7OFUUT6hZZBE5GskaBO091bPGP/uWbyl/HRKnr4hGzCYIDTRBHyqR
Gkin5slNO7VR4i/bBO5i+p1Uf6xk4FpJBnxhhuI9yVJ2XQIf13bbXvOdsD8qytMC1E/ysLCO4lJG
eNKnqtR79S5Dy+o8Mr1DbHqNGA5l21tTXdiudAw92ijbMTVSKS543PYJYQZC6maDuX513vCHULD0
ckZaVy4iHkP04Dbx3F26UYssxiCBkY2E2KkUIZJXZIvtyrCcySdq5NakhmidTnT8p9IqW6N2ENJA
rU5r7PaRCX2ZvE8E2KaA6d5V7ClmaH4X10VspkbibU8dO+ZGld7uFvkJfgwUBsaA8J2fdh/6jYlk
glbAVWkzKzLqEr+Pvt54wZCX1hsxGsFWgUZyIM0EgZ34SgcJ2kuhtPZV/HOfjW4xGKDFBcHpjgh2
qkAA+VM5xNQXuPjrHr6iHsWaenli1rPDKcTQ8+W8N9n/eSSoIMEc8Elvg30iYFCyUDsWCA23c7wp
gz2jLCaLePpyvamwyjwJEM244U6OhVlOX/wu/3KMeRP8K+wo2q7Ddh79hHWPmQP+YSwrNGOloq/p
Epa7SZw1f3eNpyHhYGh/74GXeBLhnRr6LnyOP0WrPe5iKcJdZJtL5fKWimMqyyu9/gx7smzUVDIr
gjswomgw/9MgXZthhwsc55CpfdGfrys2H0blZGC+XRRRrA6cqD6QrMge4JqLReMXvcZUui+LIBtT
RPyiysIjPAUzeyNBIKA4G7UeBfsz9jSIXTxDLhAspo3KN3lRn9yTohLkjGuhwQAI4BnFSK6AEZJG
PAopsUgbqLj0ZYyBY80I8m4uuLQhvd9Do7MvS6WNWmURXDZopdvnp9UGyd4IcgSeyWJPJcs6Dvx7
4cwL0aywtXI6GM+4Uel2eCBM2MXiuk1nOp6GbcveocWQfKH1jyD3aNQ0lj2KNmqTkZc9TrvEA90d
h+eta/2+zZ6knnh4bXelDFNfv/zZioXbs/0gsvTW0OMWovDLV1HvPJU3ZeNORSJWvfEpj0EZsvBK
4GZ1m7weaBMqGamBjUsDoq0JAEBEJa7VqcmFyTeEkkryaEkT6bLKTUMnquWAWx238ndPA27Mb6PH
oXJ2TC/i+zXijC9UcylOF3y59Wo1wN5rDjb+JPyAF2PmaNgFw5fn97bL22gC/5OlhChB/Ichqt6P
n6x1AcWgXr51nxxiAeGQmi+1rjTuZepqMvHrKTrxC2UG/MIo4sYVpY9wZDUIcoAaHom6JW+K/XnF
BJK4LrZ5hjYqEHFd7L+6ELXnMbGbonrLEjuQJEgn36EkBB79+Yh03RxzeoJOldAH++oAx1wlw+XB
IJ3L0Ld1AE1VTooatgj/Jdl5lj34ZGdImrU8lMZ7IvTfwjy2ho/LQPa9URGpA0G1AciOxLIR5lFg
XrFE/WkbxkxbH49I3It+SlzpZ2yhNGCIb4l2870Ag3TCxDGZ21J5tH08iGBz4vg3e6vXHK8NcqMt
gWTiy2PObYlAFt7KjsJQwUmAI//Ewq7GRMSoIRlD1Hl/45CHj9nN8lHIWQJIvDrl2MQBhxqsGsWv
QpowQ+j6wxnQ2SqDBuarmT/TbzCRN6Xns2zRzbFmh+6R0rCiv5+W0DxsTShm03nWCM6/R2zKfkZc
l9ZZGIXIZ2W6qrwp2oD7uyxLB2so0LHBL8v22gSuS5Ipmt3E5MTKb2hmhy15b5g8yLWB6Vx9fBQr
mKROOLngnUtaVewQ3fcAptKsMFnek1xPKV2bq/xzV3rp4CFSeaKzUEvc2loT0YT3G1bU+OR4nFcl
tqUVOZdinSe/LoIGIERDSgGYGXLiUJNSlQsMh+I61QxTm5jVDvs+/hzWzwiz+y512Sod3y2gcvNO
2BitvWkeaqmwg9I9oxAVjv9wBtkbVVqLQeQolGTyRJjOMxVVoN/5BSKUS2wyVmaA2LnsefwkQ3R7
VsP+uquN5wDTlJPh2Fdg1AAxCKM3o/jqMQ/wTnxQAQmjbsB66WvlI6V7NabZaGcWzyjo1kyTn7Xu
UBp2GAKieVwjVUvH06KHIp8PodNZnHQQ+1iTlzCZGb5VLRrzgZpAccVb1VRAx+0Q7iXrxEUxxYNH
e71Mz8NZgjrytth4KyFXAFl/A3lVEzcCBT2rzNJ20wZY9aae8lQOBD3J4XAYH4P3qD91Q1/8zSSk
wEnyHAo10xjt7Gf98BA++jdjtZCoBdISg3NMMLxC/kCP4mKsLoLncniGocZydLgpaUmAtWvvrD0J
rKTAjG6sI4i5amlH9S+fbccURzKUMYlNuLm0pjL4WfspD0km3e+0qUTLfqDwp21yxtsA10aLg5kZ
F/U1PQHWn5LYiCumZRDGWMOEAWCq8M+j/ZJaVoGJIltY/OAAyUb611uqfwk5cjQnKUvTRFMUsscB
Pck9vSNU/q02iS3hF5WyiDxptiWtUsNh6iciOrwV8KbdTHyFw9xcCWwBBrwuumrPufZ53mQJGtD+
GfJezeu6hfsv3GTovGPhUpJJt9PclNWLDCG+6zH7E1i8FruH2pjnNh4St0LKldbAMfsL4qth+OcX
YDnqq3RVNYM+oZP4JHqW3T3eKaTZkPCAezs+rPTR1/Sw9LU0/BAIEK234TYhLYPYfqZfnJVUcM20
gLVbsg4RYGcH6d58ah0UlyXT7VwpQTpfQBnFGYIipmSk03dLYLKwN9wFGneW9lF+A2r9/SO2nyq/
90PxzmMVHEVUEKLVwqKVmTsEqdh8gpfurQ9VwrYlBpfsS1sl3iC0nDNBZqeShvYP3FRBWehyPO+X
To3bXWEVvRoeBIWf2X9NobUe+Ng1am75HOqeJdKuZUeZN+HWX6w0mneh3VppwbnHoJAKaDfyk3/h
YMyzhMPM7A956kxJEYxA9sCC3WtVNdhKHBdGoIcEGLm4xfor/LLv/5JNyeLMqaipe50ocEmJSUaw
/5YsmkabIxeVjya+obIUdakH4VR/4hjlNb3nDBP1kB72UnQcaz0Fib4hr/l4jYdQJKZqX1ZJgdiI
Zjs730fkf4M90EjG6jQhF8rkfz8htxo+Wad/TrqXQCO9sHXhcqUFvcPOtWBx1z5WPGbEcQb16y8c
srvxYVWupsHq1V6AAFaSFA2SQKND6jIJ6dJnm1Bz2Lzi4ytFGabnZPFFGpTunx8OQOl0FI4upkLd
HZWlNEmRuyOHrgpv4Rk8BVxEntjfBgEqqX1ARKUL7xQO3amp4uyJIsa3pQyGeYB0sQV/lUmrE7qw
ebnXwWh7bIodP1EvIDFpuIuB1jSXiDfn4fzakUziQaXhFbb9DNEaKQmjkyQR8iK7XwMLGEVGMV2h
0gz5wIHqyja85afGph0SEIC0CtFpzTP++tQjPgbFCNjmfEESQtmTTzd3BRi4Xal1E5roA9HVJHU2
55dr/DXZxgVXLZG1wD75NMro/UoWsevyI0EWSV27INWwKx45FceMJjcbHGuyUxIoHA95K/btfQr4
I216bkqJ2Cff1fFK4bH9MSFkpnAshm+uRmnP9+0TWKtoUfqZneGJbccpWnchOTdZ7h+fVqyb2TkL
WNqMKTslAJ/5XsyVgV/3kji/rdk5VNhB2Ek/3xLZmXyijNNja+B8VcThUokxB91iMcmfjwTwhMOk
VvjupaisMYze5cpH1tke3XHVWCUTiu6j5z2XHVl328uQbDTPmQco4GatWNLfDd4ShkTeNKEI6rYJ
CrluLM7cnpmF51qhVKvDDHiNAIDojQZJx7vVxCalo4zwLYcpmWUCGpEk6chPillF1hBv56QL3pLu
4CpL20263EL5U4gaKIsJMy4qdb4lqmmGKC3d7U2OISZgluY3jVS0zZvly8IDwB/e5l1y4wWXcGR5
z+qy69ihOP3j/T6VPuzp7YvR7toPLizf2FvSu4B6Bg5ZMz/ow21VVG3QAVSD8rB0JFJD1dpjT/GN
HsIReajtaZkhw9kEm9xxGc28TD2Ann6rfHLDBSI5nJFsCLrtZsA3svKi56JtPUXRaUvaTYZHQ44X
bZG57xIexmLrYfj3XZ17S338ZNSLO5jtJQ96rh2FcbhSSm8GY1Xzm8dDxezmurKgDUilwC13sdgn
eDcdKvfgP1dqsLZLbEB4N4XdDMrSZ4z5RCAF8XDz+T+1HL97OzbtXnBOMJc1rhlh/mUlhHFmkk7j
WU6MildFLvaKrlnZXnEf+g3dulMPyQYVn5KUFTne1MTdtTrSSKvM1kCqyk91wAgfNJIezJE9usHW
b3vI8IdNSvYJglugYbDTie4TIb1Ir58bN16WfRSCo1e1yWEOvDCnIlBQ3U3h0z/vVLeGP9CrcYua
7yfaOAhtWsvWQyPGx7AjUT36kt65bD3ODTg82Bgwk7XklpgiT2Tv0tZT2L3vtpGw4ZMjixb/J+ua
Ad3HY8eMMI2KBtohQK0+G8mm9dGGjOEGWdc0TxMA91y+LVVfvrNQyU8AENK7SvkZQkl/JKWAvCnK
pcqOJSIvS8wkPryS1N6D75h0q5uINYZ/TfdSrxP8lYYWUNo+f2r8aIa8jrxuO6mhgMcyQRqszfJz
mTIN0BcYAwnHbezE8SSGgqyUpBvTt1QMJTmbi+ne62loEK8/kfrBLyITcavru79Dtf9ATkTJjnsm
y+e+Vril5rua2u/WiHES4scaoRzlzxhJn2p5pnc5PQazVEDfjm9EjjF/TgQEk8Oefdwj4ZHWwWQS
pCzIgRgBz0mhDRUiTw6qn8M3cc7lYm5QlHzgw+17ROduyVD6GRxC7jnTpYSme5IvDk+9GyOXRILp
B/OpOet3c87O70Wmy2urTTIac8awgnScJVhUGT+MscUUqjlOJhS4x2Gc5Ix3ubKo4bfvHBxctxRy
G0go/griWiIdsWfNSEByJnc8tx6ahN9JQeoZnGwthTjQMhdziO4d7vO/84QHybBReOaixCUP5Tzt
ooU2teY3bo7E7MpjqW6qlHU7vJF3hpKBw9qJG11Q7Y+3jh0lg9wqa18yYoIqmZ/som6YZhf7hZxP
iR/oDyl1kTWRf1ziXHtGru0OxuJo89DO5vCLMXliEuoQjeBiHIDmN7ge8nO1pb4SHeoSmGsBzPS8
WW+oS5silWVcUJE3yNDnG2L8CT6ZNs9pffqjVMqaIGtsMH95kRHkNheaskqeTr+FhCNd0CWKmCjG
YwzPddo29/J3b4AjkFGCNsBdNWVAQHoIfNrroYMmn8E43KnD2dXKBeiWbiiJXtODetSyO+lPeSs2
MJ/1fiNlAPbYWRXZAcTp3tduuHoRRraNw/nAHfvZZesxqi/33EhKwk+GikF/QLV0VTjvULSp31YR
aWpONidiQ16vkxxyShXwEeVI5IIQulfR51qG6LdvmGiwGH37mjDH0255piO0u61MNMWxwgFStscY
d8rJvOxIr6vDZcWu4BLg4YYGpFC/GRAjO7hXzN0MhQe3aLJ4W5hMrjKd7CvrMfP3FVfGfygP8FyR
SzLhZYlbdElrxUuozg81g1THwTqWo2fQqMdJgyVIJtDO0cUMK7N7KjnrQJlNc2lh4cvNVrttwqZK
lg2bdAlnnKfuN2zd+yUMaUaENKd9FtomnA3qoaLLCfgr8MEiw/VD4bm6IgQdJXMvNhQtIegrPxUh
vbH1LYApY5Cir6mab1/LyAFL88Qzmiijmnat+wVmtIFq/ZsC0GqfS4tlO5/E2nnOFC9KBvIy2paD
GdyFjqRRQQo8nbDttzyvZogNSv5eXTGzYBbP6F9/6b1YKF82987G6nSB8AeXEvbYqcfqKBa0OYgm
Fe5y7v2ORE34yjcMq1HJ4L8DCfy9yyea2w8JlyymRWtAkhEqTDlydx6d+oUxCFJcZbDpiLZVjqje
4oclybpBtooP3xqFhODa4raZHMD/6MRr0gy9SW9fWhAV7AcjM0BwWgKxnl0C/milwR7pFk1H6wSP
Yiy8wvvvRCznrLtijZPpxI8ZHH0zbeyfj9j+zDBuaWPVF3f518P/kyy0NntfJ7z3JgDWfanjZ3YE
lG0AxyZ/eoSovI1A3CDUOqh1t6Y3jyx25BpFjukxuHG5vXJslobZ+j3m15Z+42snIn9jvIldhRyt
/ZDYlGQhvoLfcZ59158vQZKkIQ3f3uARA43pqXYSpesMbVLHjntlUW85gytsy0X9DYTBJ4K1Xp0h
R9gjJKrkAA0hDad2fnfcarakTsqpeY+AvqjOxTpv4iNXjaV+qo/736Ft+i9NC/R+8HNn2IasdTbI
leBveasDMr8y0tKoppLA+89/AE2EovDVAFu01oKfjW1MbcmSiZkgZdyMxGHX0UM7ZuWi+SnMTtLy
31WSGc04euvsGxlOL/AgzE457VjfC5wBhugF/ker4f6mxAvELCfBYDeQPZkEFwn5JW45YkibA4GG
S1UkUXWe6EVI/lAEqAtv4n/y4rmvlz/RZSHZHYhpZdSXsiHwX6ARsPwdz/l3BZ2HUKB2lJK+oYeo
6JImE4fVF5SEPO3hhIXupGh6kDmOnjFVmYHLbmUqQ0ucqFh2oYi2M2bQoHXMZUTpcQOfwuAJLzn+
Io7BbVfWUomlaK9w5kZfcRo1Fnfq2883wg63L0C1jya7nNCfN5kF4ZcuQa31nyp8wPdMlbFZOQeW
2eX95bggWCqKSyvASkXIHmfxHbGjgrJnLTeK1z5gL2YYF93j/l7y5/s9vxmviv7KcUrzqMCepmWA
tAt61c7YD6zFeR1696c0uVdJF58NcGVVR93Ywd1nQuQrHgnkcKSN0IKLColy5jHyZE7m5zs6M9B7
6+oR9W0CTr66Bp9bqkfulkC0jOoMxGonE69n09DRuQc3X1zCi3Zi4BISai7TeH5MKb5c0PjS33A9
t+MRuHQJKv0KE5lkEerG4xjuw0aLDYKJc73ZA5ylrouMHrzn8kbOsAleH+96iUDA5tn4rXiRoD8j
Bc/8NfZ1PpLkCZB+axco0SZQqpaR3JYoXDvN7H6KMaejI+OJDHLM7YboxCtK52uxchPb8Q0QvpRc
k2GU/hdqk5t4hVB2Zzt0UkrpqLqORgZ2Etsl83APMFngfR63phPkngoMMgvsQM75tUYsM7KcnKUm
NWAEreMRFJEg+auYbnb6b8XCAj3dsTOnQanoHC2RU5raZcs8o/+fs5gTyo+PxFPFhcp7z5ySRPHD
2C+VMwdgBfojNeARtC04NsPGHKGSmA7fhCGtHVf5YqmWygq3gfLOusnu26JY0ImMeTFBT+BWKoMc
HojL7hB2b3/4GV3dl4StDGhUDiCwF5+/xGnaQ5PvgHsaZsjZ/igQPZaUbFc95+vgjEtGm1p6Fn8O
tOUq6jOrQHIXf7NkOsp+Q/0pCMigPMXQhXc0KmtOH1hHrkzPtUvmkhOdgWIBC4p/RJ1gBRcTbNiv
lGKDHn8g1p9kS+10vNhETej+6oHXi2kvynVZ2skW4g/U71d996PfNDA2SOu5py2P7nFVm8MbNMG5
lLMhv53qrWGaHPuKkcKzBUDIy+PqgDM0N+bioDuOKSX1kS01NoKx2bhDC4wm8vH8Esx80r730s2u
DYH29S6UOxkz7Q1NHWN6YYnRUoj96bucnn+hBeiphpWkHbgXvxwVB2zeAfKtbdMQd0xgDUf6Q7HE
TCKE/g8o4UxJDxBleXAK0/mUsQ7+F/8q3hXgoOogRXyLzcyuGDT5PedvxDgYNsdyijED6scLzX9v
1nRm9f+3uDNInEiFyTXjHwCXZDkVJekgTL3H7PVL3HRaIReg+rkLx+JJGSz/SwpUvF/zI5lS9/aO
wxsLsBgHjGzeW73VE2L1Dk38ltDc9uH9jvPP1RMna8Rp8dvt4KiczRsWu72jeZWGLu9efe88NRr4
sfZtveHL2rL/4z5YY8es0vG8iNFU+yyIBSuGFvLclsH5prpW+M2MsK9qu5Y/rL+PZPuSO+vZyDYr
81YwkrJWOpkCiidohbSqE/ET500AbtoUU2oElL0hG56BmYBAqyE+4RniamuHWbwlbHbfaQBcPIHa
D6Fv3MR8lCcWWnHuoF8a0OuN+8Y57UhR1/0joe0+mcWYBPJP6ar4evtF7IaV59XKbkGeXJjfAb8U
ePvVMsXJgd3D5N862zgflcY9a7gPzHWyYA6lKoRJyZtU7Jvgiqk8M91l9eyAk7DZTx/krA5J+Eyp
RYFV+DK/G8SXaoVrzBuMEiws4ZfzIcnPG3WrQPJTAPkraeO33PB4DoTDOjqjwFnsK30Mz22FPVTK
0R0yeypJ7155+cHo5JUHjvBL0a2Njuyfl72PMmqb2/pan6jmlz4sO52WN4MtTbiKJJLUqf8A94rY
ORmrOV3Jl3zya8sm3IKoVDEH8k5hSL0qXl8fqR4A4Sir40KFfbQp0PtRmXEwk+gy6b+w2ILdE7y9
lYp1khRA5Q4B+5U/ZXBEbUr+rSac6tcJwPe9Rhr2RKq9zf4bEy7SqQeSdMmpPyhqXtjZMQYvQkfN
GkXjN8zUliSfhbIfW6ZygYmCYY0TIgOHYYzq+6KksNIUeKXlCxt8sXSZ1zGePDyUYIcFttAdYfzH
Ld64nzd04pDr4+0BC0wAOgB68XtTzTaVSy1V359aaGfCXefNRbSoEoqq7OxQWzkq1zQCxqCs3ITf
7oKun8ES7O+Ff+alZtdk7Zgx/0u9ZFsk3ciq6aZURLXSFi7WB6ZrZLqttq+Kj7l+WpoozyWu6UPz
EGhO15ncIAqy+QFpO6YZbfn+z3ys73qtF/UhRpblMws3DI1jB1+Bm6+9Ff4d6/AKwZ/mNyh89KIr
K9SLOQp/z+ffX7HmytQ0iQ+jhnRd7vVOBEia4LB/sNTcq20LtYvwn6mShlmwgads/UicgC061nlq
bIR/fKiqIpjT7PEGd0Ak03ejyg4ACIT0GW5KCIrLOcUqMkhHvt4ghZUCGEdve3QOcxMtGiD+Id2K
laVrDmXjmextkwQZFyU9A+1BpsGESlJCCxda7daLCWACWiAj7Q01ElWBIgd6k/7GzmYWcYpsRvzk
bYYX5Z5u4aplQhxdH4sNjMiB8mpnehm0qSGFGJ0Uf0oaQhpchkOJwxvDWbmMDrrWLD3OfoeMTW90
B7GmXDlSCnoeUOllWWQwfsapVORnkq7EI0eNOgFeC3uABzX2mVbe6AGyRbeLmlwy+hDI7eJiAptz
rBHWeeTheJqpSMybozJ6JXd6WQxr8CT8tI8jsp6bERGpxX98TxvXNsDdtbSd2fyKbEMya7Dfw3Uj
+iV5hTfgoUMLsXwp6GPEnZjt/nYroikjbXuceaRQLXYorLd9olPvddQl5M/9v4SxHDfMc9vjXUtX
R+rZ4nTNy1gT2aFbTfMN3aVwZUf7twWCOINUAKKf4DHV4VjMdYDJQRUwj8lvXL93tv5xm43pWjdq
q59TYXJuInMSEFDDs+x4tcxVf/I/SljCPEoXIWc/0jdXiRj7MU9McN6Z4cXllMFgKBjIv6+QHP5p
a+IzCEIID6ovUHnvu66rR8cHjy13hV/FCHWSV1jQX2qzOuEHoBRT9c0ootte7Bwx92M8ma+ON8fB
m04ilxERUFg7ZmySqpCjQYxRaKmhI1FyF9z1idFeT398mja2/vhlaOaSjiBY2S3Uf/QWjrv9GTEY
3x6BD3tr6uTNQuiH+XpRenKh04NeLh27VlO14h9vriv+dhX7EOvcApFS1U8N8oasXVWL3x4aC8x6
95UUfMU1nbAdKYazpOm9fAr1aDzQAL6/pNr0EaqxuUAltjoRfVnpAmNakMmy/fcXr4wHfLo6t6+5
c2cwZPyImiAVOhmtvRTqhH/FhL1zI23/MT+s/jzJz4GFpaJz3OF+I3A1tpJE4bs7tx+cZqmhB//A
c0o62Ftnd3Soyr6wTfJd49gMj9fpIlHQIB3ikQtdBbMDrcIufXbljYb6Hosa0dKn+fJa9B6Zm9vS
uykC8GsKcAAiUOvWNLWl/Wy1wo8CheSEp/1N3QaP7gJDdFe6JUV+ZHeIl3NL23bmhrOSQcSZmC8t
TtjkAcNI9jVAP8jeknbUDoMd1RKx66DjyvdeH9aj0dts+wll0KFadyZxETcMj/ssO9397Gqk8Ab4
tf4DFtdbUB4X5HqN1GEVDxLyKMegjtEYQrgOqPtRJyVscyogsy4l6uyV6j3nNqBucvUvE3VRLkL/
0p3sq6zRhDG0ylZDV5vybyEGjBhRmbWUITpuSm+OIwmFiA4tjZpVcEZALrLJAN7I87A12GOHFR46
mjNGbEO7AXn55WBF2TsYbYkq1rzy3BELd/HspSyCfywDmNG5si0Lnuw2z9TZGKCeH2vMiwwCLkWI
5CvOa1xSnvaz8bAfkLxxOBAKg/yscxv0XZmgm037b3DXFObhSbp9981WmYj39Zzq/PdY5VtHooXz
R9DxGmcy0SJzYgKK125yYKZ1mTKOCRckHBarzpmjGpgLczOw3g6yGffX+6uQ5g99Y5wkxE0sypI5
8MtxUtwFhDq6QHEQpONQVUGLR6BuwfwYdsdvkhy8y5Opb3pLdWEZfD9GEnU8+JN9CBaXmgmM6R3q
zpmUhsj+/wRMHqyhu0d46pBVedyCrtHV6rzyCPp3b3XYcv1aoDnLnKleWoZbBA5yh8aDEIIqMflq
gOxxdl9Z5GjfZpwXjRIy+dneDm2u3+4OOsWut5o3HD8ogD1BbQkiMwiYohKU6LtM+hDd/q1li2t9
/tOncekbtB9lhrIVE15wzxHDYXQQUVXRM0lvndMZTzLlZ3Pf9B1CX6DX+8eMHBAeCsd1XrqPSiEI
2mHCn8w0hURxKNrgEETyolS04t4ObtEFr0qQEXuWS6Qpxl6yl8jj/HNFdZUeG5TpQC3LypBRLUVf
sHBx0AaqEPL6SvD2/BLbGkFlPZsnhzSI91BJe5cAemVp1F2G2J1pcBTu8NGEV+PL1GQhIjyV7XWE
iZuxi10Kb8jlCHR/wm0MFw0ABrSz03OMIXG0kth8Nsz/AwBEWLw2yDCu9FYTU9Ba/7Jq0PaJOnSU
PvM2wxY/rYQCQcN+ZvtidYwYgQM9s+cdodT/2hPAh1S16v8GwxfAHRSZOruj2MY7471DsCsiB1kd
Ujcddi8Y/yixgvfzxs6YPmyGIGQrMs/mbPH+nHwAVVY6ZeL1A+CHQLrJO7ChrwSK5NjkMXUT3Oz9
ELUMqEpLpjgenIYNSm2fC+L2toB5CbSnU6RmFaumlSKCxiskCKHKGo7aU7LvNUaKn/tmUsowxM3y
ABB3r4opxTs9YDrWOaMznD74d9GKsZOICPvneoSH/xeUyKIo0p/UmwDVk+BH/oLnwGUGeoSeygH2
+wPTZbDfNTUaRFeWmmQT4xFFI2d79UPG37z7oikwrEFYE9xJI2+ia+pK+iCalWYLQkq0pWglXM4n
+eyrRNij9DwnrMzjdSseMDJHufdEbE25GlLcFwfnPoeeim4sefpSOHKmRyI+oXlSW9H6I2VCGH6R
ObWJ3AE99WzS5SFA2zGJytCcejzfUEHLkezSY9g0T2wBJ7JXyhpY/4DXjiDrxVIQf74pf86+K4li
9ACus6c+zc0n99Y39laAAGwD1Da5TC8fLuFBDwOHpn14NM8IYW2qy9KeOKYZTrkH9Wx68i89lp3d
xilYWRklML0DS4Av/yL30oiJ4agGhi2y1UMe9h2erB37L58EpQNKxw58L/Xdd3ryHLnUMu5bsm6v
sm7XusYXrXBA397OGA7PugqhZTr13zDrFq9N7yI1FpX0Resl7vburd7FvnZwB+0Br1EqiZfS6qqg
xuNfVTtEP/dW3428twV863PEhQPgIOu/kIYDH4PwMJiStiCEKBMbUX57VvyzuJ3IKMVLaVBLOClq
RPOFVgMyhRE8keIbLIBJgpT3L0cmSOlm6qZ13+zL7Uwn+3FM+OOW9Iu8wEf1QzVbf/Tf8RNHaA14
fV2KU9SxyJcaqgXvnanyoMbub5SeQ/eR70HjLQbQeGGV2c+Jo4rS5sN11ZVKyeL29Yx3vshYr1sW
qXMVdrgcMA8ob5Jqs0aWgmkr1mi/uOtNqLWrZt3+BdBquvigCXcvLOjwGB+wma35nsfWH4kAdEHr
7ab1zkoIfWS3GrmdAnrYTZDvOknAg9WbRlg8LT54U7hQ1HgFOKZPCwScAayaSBat2pon9ISdG7CM
Vfl6uCYNGa05w2qF2R0/MCdvpv1TrPqnYHdZxtipSLrE6mB5tDWj21AY5JOc+uFFPXvTPxm86xEr
/r7JvIR7D790sNxcNGpy4+H/fZqBhB35cuvvYCOUs/B37luulA/hJPgMg99zw5i/m5IYssmCL2sW
uQ+PxNAHYUvGlZSJyzlVatzyb7Cuh5B1ahT4BVBjzkYEWiZFgly5Iv3o1JheFF8sireCfR7/NVA/
c8LhBasHTlhvXKZu7WxMlE0p2N1nO6aa+j+4+69iQSBVHbw3UzePeBWTxqutZZ/GwRUj+vGCD9hm
NrzJLhmLrH0uMc5V4AJke83IjFFUZXM5bRNOVM1PXFeA2ge01q455JNlg3eHW290V+Hx4UE/eo3G
7h010tpG6+yhlVhLBCuXsbdf2FfuAXoUXX2STxwQ1FS2OyACyC1ZI0YqRiUZIzAD4N1KhGVhqE/B
kA5RnkdAidxlwB3/052fljKHTqvNobBFfahgbv3K7UIRWHtMkHyPWlMeJK5T4xwIMp1ryptWzT/L
qfBPrQlTkuSipFAktnbAmtlzbbeNlEhOZnil2a3c3aELY0TKfa5oVSkf4aSjXlArhhULZP2S/Pe7
o7YFlZG0IvqQjEG2IREgO1ewwe/bViYzdXQZabsL/3j4uf1PMRrpfSJYEdeuElOvntehTx0zaGsJ
2+sPbNr7yXnn4NomRig6cTEJJHg2ihLOppR/rqEpP0V/FewsCoIDZnffbn9f3GKpgCINaLRTCwqB
z7SWMiqHswWfdWMoMoaWYTCotAK5pfLl76nG3+PpeolJwhvH/eJv/aFQ/1wvpSulHu09enaIm4Ho
o3b6ebLBcMbanimbVARtZx4FrlrP9wGoa2GjILselNalCQyaT1+vTMKRaTQUsIlhcwH3hDxKq0my
X+5o2V82Ih6PwDoEU6hUpI8gMvHObVywnQaUu+zUA6NCALWGTi5oU2sd/sNqEIpop/6cQyg2qFXu
6U9lb5vJ9JRRMIH2YgLMyD/v2VxrJH/FR4pI63jCMsb8VPvMlgAOGaJWX7dw8Rh5wxN2WnHQjkeo
etM9uXC+ALCvyliTj0n4DUfwUUPRhu0V4Jmf1BmyY95Jw7WbBpAD6qD3PJERS6LRE0mC15kXEg5q
z9cBrgmnGiWX5bS1ra+Vilhd/ckMUbpmIUAKHKU/STTkmZjY31nAxVEnfKgGWj0kDFtGzdKgq5eW
l8zPUzg2DVSeMWjO4Gqyl0ux2+GCe+upOOCKcqJgKVE5+rqSOBzwWNyDkO/4kx/AMWevn/huJx1E
t4V8ddRnqE27vvFI9zUvEXB+1FNgsUYye9yMx++aXpGPXvKs1Mcqu0+fTvgey0RHCcRsy97bOivb
FD6UJZ4P3lJ5n/l+4fVlvbqKTyCzxb3k7dp4ryHi9NmWUDh8VsM86oboE/jN3W+wXp0TZ5f/bAd9
fh/elVxfMwDxRzMAVteoCHb0Hz2zTTb7xN9x6omemUf73V6NFEXj7v9yLz1NTVR52dYZr+VlE9yt
BI+ydydlDvUC0Mkn2itskjtWCxxZD9vuaxy+z4V4JkTK8znJO2CD7rZoyGtidFFvNXgOyPtmdYSA
d351D6mnQPpgF7NuBSQYWbiOIYD6gaYXsBCgT9DcSolQ63ySUwdQFL2rjvxJNa0HbxrxKHfCebEP
5iLl9IO2PKz7VtCNtzHenpkd5FUS/IzXx5Y552hmG/TxQeVxWLcq9EF42y+tC3BgK8cWjrYoJYcz
fYYh4or1V6bdTyueKHPXuK5PTSIldTW1V9HNbrZfnj0TYarEzyLlcTGkhCEuT/3SwK0UsyUretFA
jxAIW+ZMo9CqHZQuG8LpZXjhOXQYurvIrmZ6gW1wadK4H/hq4CFBmsvYH7cePsrH0JExuKPN9JHy
jwO695EHb/IkJ4Oxgo67lwS3CUyrVMlMT92KLvnBzpTBFITvUnUNYCKCDkPwa9I1+ucoPuKq7eXd
8kjCVgHlT9XMwlmw4bID0VUGC0ojFISIHTWAYxJG6A+F7c1mXszAr+QA1OYYOeXK59m41BegUt/q
9kD6+amTc9XsXYOaIWDFM3mS6AZuB1jWz09Syj/lgC/YFNZNCPGp11tsbjPPMdRWm+qan00amCcg
enfe5E49O4QG4OZ8EGsTYx5/iVRauhNprEUqRLXkW/UHojvnWq+A++iFXdmpYzSGlfjq/lJa4G64
3OtpwXnWsS484cmWIjJV0YDOB38ck7fuRh/K08LEGY+MoiVbQSh39RMOvUfkxV5yU+6r2k8J83kb
QO77hDeONsg6LWTnjKjtvu6r+7gs6mwGLK2aeZqR44oPXDH00di+k3VB2UsRcC+QTHWt5B9BZ60H
WvxlFoVZAeizLzAl4bJGqZKcie3s2PrHAPZ/ppMbfv0I0HYlHT5v28lalyfgJ9tO4p6VT/YJoZZn
j7YLQpkM7mnYs3vExmaoqeS3NMEX/4+kTzdErev2/7Tm007xaDAR3PBQBQDEweGfzwMp/UMLQroT
CWQpk7tTqyIAVukM0tjVxMi9csZpPhoiNadIsaAITzQSRRTgUozRnCa/FZr+QLfDx4X+ZJrL5v7B
5b2PZtsuVadMELXi7z47IdyRHTXsyn4LyTS1XY79HTVaEn7rFDLk3xiwVld0hiN4wRLK3dHu6YvE
szjnqKBeOujZQIlhmnlVn494/D+bXXVYHRvWtD2bySDpA90RI0ZXyxDHzColN/OYHMiDWgc8QpiE
ZFMSeUUsPIcUX/sgYCJVZV9CY6CfxcIFqCRvkn9bkGAfEx1M3CjkXhBjt0uCAIoWjuXKSFWcGpQi
vldbfs4F3JNrkbFbQb0sRyELlGUXj93xWMbHa4nfdk9TZ39RTzRCj78OOdOY0NRAHoeooDaX5GA8
fh5rKY8WQBHlRzSc8zulO+L5m0M7s9KmE/iixlJnHz5xa+4Oas00XkfDuPzghcoC8Fo1AKYyBvS/
jOa1GCn5Q9DAPaz1As52kmr+jEdTuDKS/nJ/Dm9kLOqE/JYxeMvIm8gFjs4hP0v8SGVsWx0GQf7H
P8yk5k7DD3/2apRsBqRauJUN+WvtKKJcJx6C9XETwMkHYfeCah2IyqV3MH9eRDegXWa/AFw4Ka8p
Tb70vREaxTU+ez4Z+dUfRf/H1JJ9W5RKQKq8S8zGfQ85g5qb/NeC3blMLsrvk/YBqh/bCOGrFUww
h6XEzpHJ5Vk9v/rrDOM9NMXUKpJ39T/OqDB2annmlM3eLoDV3/efFTd5naEi87Qy3cVWqkUQTzCQ
MfbETNQfQxyjHdrz08CmCtt5xEeG9VlxuDa/mP3l4rGFKb/ZYy/ZUGVTpdLb+QcsMynP3cwE1Yhy
GD+VagqYZWSCfdCAfg5S6fGB2pzARhO7+M6JNPt78MwoCNw8y3iVocvalF1CFG5lYsJeULXnNFsy
hZ33SxqrZAvgfp4tCY5kvPONvY9L8QZhZjJXClo73r91/+PV5tr5k1Y4LMdxNy6gptQjgYEVUTo9
9t7GFQd4OaFA4IF9vZa7VL0neVuqtc3FJuaYtYu0ufas3FcLzlxdx8Nqx1jofBAXoEJqS6dWa5ba
0uzFjZdbd6b5ZaxnVWjU9UQGRYzCtwZG8/SaFHvZJl+wcMtUAwUSFuZb7JRyOSU+ny0WnMzbYH1A
JsGlZnlT+w9mNIxsQGmLOHHMfOdokZ4ZJvP0UdZslCRfhpjd25BmcCNpNyP5vFahDUx0qyBmXLDk
VQkGLoNouTwC9yrEv9olW7PRrh5rJTU4DjvhI+HgZY0OuIffgvjI/UQH1IuhAUrBzMvetoYJDScl
tOVaMoy8Kp10UfiNBDcO4xGGzlv/JjuUsBNgSakP1l2W5TUt+7eZWVRI9I1jsqezJmbS/LHCL6B+
tmQsMWLBZ39TGXdchFIw8i15QlLogEI8eGpH8KuwZYvWUj3ag2gMk3WXeJQTD2K9Th78XOS+kGUw
R6n2IfthVfgsolo4OW0DSg+C9yOZ5wFjsfr+P2mQ4Rttpy1kmgD0mv8O3X0NaJkzDLwnyCcrKp05
2csbnBhkhuDDWJhFUSqzxRCVAP2Th8p35crvGcaFtmoo1YII0A24OeMIvx83YLK0gM2nncNLqXRT
u4PFysJH2z1rV8hstxs/eWEJeUF7XCbNo1ekklF1jwuT+14iZ+Y8Fjkp/ZgKT24/c0WvEVXNCMiO
RvEaj3LkZ4WKZC/n9EG8yvGphGeK3pzdgqrmYmtuMQ7hhCQqfoZvbrjolLej33kU4Kf0lPqu7P9N
DK8lkaKkc8rxYJv1a6PDlf4/OH0M8dzQYXLQbGq+SviepvvI1VAc10xFlq/AEtqOEpzxG0c6xniH
NjyyCB5QF13uidr0AejqChNsXoRxWxcyKruvhAjjhZecmiG8SGJ7nuelCBRhFMellLJP+97BOAVD
DLXQ+s3CFup0BEnzyMouq1HPiYaJsuYG05ILwpkhjpq5e6JbWcadJVwIHdST0tQb4sP3echewA8Q
kAh36KSDAeZL7jG96j4rI1wd6i/SN7MM0TzzXnHPMDGIseXmxLYpMm0D5297XMZR4VoyF3T0zzdB
us0sOx6h7BCp71yQXljzoi5Yw5A1OBmMrlMqrOUyPaQ1cW0SECEU9GBf+WdABrRMpqS7nJ9CbSmw
H9R0xon1fQLxlbbf8+d8nBgtlRJF48kCJVmpc1VuMbYVHdP2VogXIz6iT5z43IT08dlcAmC6ZT0Y
EfbAlW2Pi6nwXw91TM2Img6MFBVUaw/FmmsH/GvLyRblI944S05OJihdRnh3PcMuNRUDDWHOj+/J
cqWXbEiUJ1Oako/N328hcp1uFp9XbaLeVkR4dQrwResR8Rpuw/aQQMMqS5tY8bSW7+dDp7mMjHzl
2wx7nyib9oq4U2nIG8OqdykpV1utlZvBqXNZddcntYLAmYYPpvxCtLGjaHDN6/HVIPy7yxlImOgd
i5baG4BNsxJEiOixMg6j6EjGjJOyBjJcPRKP5FjlD5et+HAcjPdknNkW6/ISAh8fwsylkcbwiGyI
9mv6T2dwaxwAcHas5xKH65aSR+noqEl82JTaxKnfy9bqz6IScBUl+gbjxhNmLhOy8YruL2ejhwwI
Jk3LsKuLR/z2xp7lRQHqPfQwMDUqldrs4TnMNvN2Jy43wFeeLJspCsRsQ0FapVYehARA+/82j59D
Gi9+CF6bknph9Ou5tMXnY5at4Wwk2YWPwnG6FmpPINpTppidY1kxKerDXLD3dXwuwsWLhs9snBTT
VVewoZ8xBmtH1AD/pT5NclH1Q1t1P/luHm3wBHyvZ3NEvWe1Jlmhc4qLmtPs/HF/adds4TlG42fY
QpOpD/fjxofFXFXj9+a0LXwSJdH7TVBwGspstErSNF1CVKDMD7RzP8ZSqzYMCEOu+Y2mQJtSl+jl
5y7jrcphta26ardFQiMf8nlODayClEnep7vTjkpcUKS6UYQ4mkJEJtZ6CqyTxhHA4Ql35/mzq8Z6
kZBNIxAul97d9KUHZ5S1t1e/xOl64k7mMUbmoXN3OJTFz1YlVQnR6hyO/4FsgGOSYvl3/w9mvI29
aSNVBrbZDPhlADyjzVwvv3gEc88AbVzciInslhVahMCgu8kD2lAikKGCMVDYLmJvK8oUSghQPkjS
YePxbNg4vQ5wxa3PLaQp5CqF/4tSs6J7SRMFsprEfy7lxtEdPe1pcwkIdIfRAMMZNupDhVd1ZwA1
N0Jc22w/4gWfNas3logyU1nJ+vetCl1yJUxA0jw2QrS5O0kO4LyfGRW5XgZC48l0ZRECkXSccStZ
L+rar3jJ9XRxCvWH8/ynNzXNIYsZM+dwoRj+aLWya5VJzjXzCerFv5Z9pIEWTpHc5ihquC2fYNQh
6jI3LhGRIfjwZfxkOGnITREEEZLFhC9bAKSG0a66LGt2Folh83z6sCXtziAWoYmrzIgLvJ1y7y+z
F7RLnNElHHaJdp/o3/tJBMReaQMwnP353xTDeDtcgK6d9f78C9Viyl+QcqVO5FMP/VfUEDrlilOz
34a7dcBOfX9FCT7P/Sd015PZryn5jXLz8er6wswAD7eJi/YWF0wwFzvZ/kFNK9MtA9TKth3S1395
PktKSNrf468F51FG3l/oT10ophCT6AhvyF2+qmY1h26t4H+LE+up18ior6lWIWPkxMDDhGhdBTsF
xf7WtDo5NjaChlaT90AJNRlhDeXk0EBo/AZFzxX9h8RPKf8hGwzt1pPgoCTjINtiH0vYMZjJB+45
8xTSfi3Nh5PCFtLZmmkiQ+2pgJPW9h7VZdYvG5EjLVSyKv+r+9BDpuKT2r4LHeYpRcbUGZLraC8I
y1sKprRHqkuvoaK1CerQ0HnXDRiDIQjJVydIY8e4z64wqwMozbOoGb5rVrChG9dxgbpKovLGQ3WT
w/QFoAcAAvmENtXQqwcHuvT8XIVCS1yLPLZj8IxOR6G13wcoBLGlUCCjQbJAQ3k0d86s5aUj+8UA
iXy+3VNK63gk3RG0LlMD/cJo1kfsazswl8sYROleHhVG/Lt8uQRj2uuqyyUMhOvaUC3hj/ke0qnq
ZxfKvu9SUL+NKX8tvuSTh5HZnZlwzbmHWLfnP16cIU9W01p1+/jfbzzygNdwwXycMfN+BGIMzC+2
VKCJRE9N72mlHW3mNxZ/WfMetG6BF8eQybgmWAh/5BMtD4pOr8bBs79MTW96mRlm+zQCBY0rESEN
FCdYR5FyCmcnIfkaeXv3GEce+BaE18uRijPaYtwgJKgk7D2x3jgl0pJLjCM5DXbEurQyKvadlS8X
WBBV31mcsDpCmBZyFu11abPOfvnwqLZPpYT8rNOlbklmDKP5+eI/VhmEQoZzGkmHIvgiRjXFMs2l
1v8xcFtFJoB9BkZ3jvvovEjkh1JkTXHOEoQP+acsGYLqLWykNUQ+TbuH1r38Y2q0WWoWmo5mrhv0
diNa0ePyK3hLmop+it68oODXizOZBJrbKx++GqfgDigySpYRzc++04B8wHspBmCO8xbDEDYuj4qN
K2DwoMWThIoMfWqLlhYlTBBzVonQ3XgzxJ7Dl7hDWqaFjnJSmDdQdEj4QnVO+6nki1bbsZzoeqR7
FMLAv6Vf40ndy2rXbEo/9VoYn6CiT7jFNKmLU1dIOhXbN1N5sVbzr3jvDs6QUnVZR6g8HAHP1T48
haknYAA0P7cwUoJ1OMyZKrdShF80Z1KecmzC8ud0y/RlhhspBnLRuaZ3KCFIVoeqUGz48OTJwlPM
r04jaxTzwi8QUMKVwWieHaw8ftgdrWNvO+YG9X+aHsJ7b5qnkZ3HYrIR7/KzPfT2xXeq/+t/t1e7
BRJOK7eLEN4xHCKKpp+kZAEm95Ck33419Mmx6eMCIPqM4XCbUs5gj4xEPqHX0I2StZpm9zJi/+2s
cEtIvz0q+tbgfLLbb0ChMVKytWKZDcSnBy7RNN7BRlAdEeWljI6C4IDyxXO9zZinUOV1MXYMGA38
lCzvZweHJ6S8ppsTabvl/rtM4+/bFnNnF/0bRA6FkvOzR9tefX2ipuA74ISjJMKwMkk49pZyUS8D
ywfjKcqr5NfXe3IDCJWtBdzbmd0ejRRMfORSdt9UL3UHL4M9EG0qUzJWdAbXPaGkrvfDYEnG2DT9
/PNx1O5sKi+RvRMV1JGRyinRMrU1o8woC0I5hOT5aR8J58cweKGo7LaX4Aa5j9GlEk8tlVUSQOaE
0SoPRoFNrB63oiMpAu0aD12+1U44HJBm8vjATrS+eeOw0WTS9EY3JhK6YUvx/BjnohH7XlWi12JH
hrYoyseM3pNC/eYqlhmdnLHTWPLtd+V+xHoWgLwsz+UpjaIX3LTn/JsBMSKqa3TH/KwNfAUfFvUt
QFCbUzpWDYNkRyRfIl+wQ0wdtT1If7oluJ062/c3YcdrrFW0AL8pyusa86SjqjkojQ88DYud4Jmn
5sWxVF4I8//pUYJXFYznW8WiJt8gec/Whc7dJpsZRyCGdThwzoWeaTJm8ac29gF/UePMoodKIti8
HP5pC48PSkOXj6xMoEiD7ADEEuNxKUSlOVm4F38NWIp87sFfs7NYcv6TlAXvg54+RsGiYPZ3QuNY
feMK3+LkFOvRv8UR0HTQKtNg/jsY9PQYQ5qTqyx/OcJ1LGHhHNiziohC68OcEu2NQekxICEm8Go8
onUp6x+2+7WwY1zKu/j6KK/qyHjyBDDuYlo5PHMJUI5inWvdP0pP3RtGF5QqGX3VRac0kxzsVQFG
FgO+jQCZ4W0VcEh3Fm0EeNLwaaaOzH/8RtlSAy10G6JT6aVV96gV9u700nkL/9ZPJUNVEJaSOlpN
+wUebIschCmBGTUlnFWfrJg3p4K8QnXERoNKqezaQ3G920V0gTZr1GeEjsdnQ4oDSYPyD5kiq1ui
qXEkx/l9S8o+G2xpp0LHHlUks8w3Fy3ouLJYRGINZ5RPI9mqPG51pSRRNY1dfHOpcvbrQJSAcilj
3xbS28ccZRNup/yy9ecfWIB5yWY19pmlcxQVbDVs84OU9df4KldAhuDOmRM4SNbVPzWF6yzFyskt
V5KgfM9gyZI4PfQb8uwyDn7Bx9BCCOST2/K108EXn9SBYmqeUdYcFnEYtFQ3rh8sZ8FWBs79DrBo
Q45ahkgxYvAfTsjLW0WUazMuFv+IMdWE73zyw/8eA+HTDL3eIb8AVf8Gm7WuqUBdllY8gdI4xUv7
y6njXMgrfsNXaysR3Yk9t5i8kbXir+VPDaNy2OTfgOnApDhm9m2eUYwin6m3+RIg6mnlkqOIApC2
3H6+MJHtZqcG3bvg4aEw9VYT1dCTlHBaS75rvUdG6RbLlcCvgQnrZzxYQoBnm2/Y9tI0cOrzz4nN
PjzsUCxUk6RPt+dN/a2S+cxaU039V+SOe7VUBjuLbUDd+e1gmlNe/I8fevyLBepqFYZ/x/kVandY
yAsTKhE/bhb06emUJpFqq00acML34PQ16rhADnu4Hb/OLrXJi0LO43bfr4xmBHkkfNwLI6zCi3Kz
X70yoKJyybP77JNCV1NfjMk8t0tkxmbwOLjGH3y23KLQH8KCJXhmWNAoX4yJvih9uc9YcRBEK9Zw
zhGrJfXdByiBcJRItUDXuGVidXHkmXQcdkUmhoewV+633wx7MMFM0P++9c29KZBy4m4ksoFaQY3w
OErQKCCjD1eeaICLNEBHV994JdIH63xakd4TLLVOuHNOK2LgaqDDOjb9930FDi4LynF8k7rGEbYN
ISJhiEQBdG6/lUA8gkQBtCh737fU3xTzB+cS4O5Gr+48vEv1f+TmRVC5Tw3tZMbWAS+fgQyCrP//
4b8EAnXs60jaWl3iNmGpnHSexVmVvJH+r+Gz82gEsPUU9GnexTfWmH4Emu9sh7yyMeDB34HumdR4
hjyLQDUCjqG56ZDMVuL8LUiqe7pjMti6qfmexF73QxnzxpG6mzV44oE+nxm3EsWs0GQmPU3/mOtG
Iz3xQHFsIGw1LQaaK1yR8lFRgZxCZQiot7n9l5j+EIFKf3I7NpLQtb6x0cml0xkDYkBUZsji4sCr
PGg2Gbhzwk6MKyR/ghYEsJgntVFZRyrUCrzJ1sYGBwEwCAbF+X+hHafXaNVeHbuZpW75TUDwCV5o
bcbEujUbKMjRhHgRkZqMG4aU/pLA3G7yRkDWBj/lHSbCdrT5rczPA1Kmh/wWVqOnkezIUlshPnSy
CdkMGtUHsO9IVO78Ofx+Abl4ejWW8erw8JPKDI+gHg54PayQUWLa6qSu5KdJAsR4LqCuIeQB/p1G
DxJ4BISAGrZV0TG0wvaI5/RFQk3Tu4vuQYbqbByBe8mlgZVEkisHDgM0XBz+cI+uhpZmIUbR69GM
dwajtqembbaL+8q8AFe0H48NtDhA58/pvVna6+yeoXlMkcuEPGP6o7ITqFl+q++rZ0K26CEYiLF2
V+gtClKyhqpinPsMewMAKder67bHH1SeCN/2FAkIdhla+Zq0+Tfbmnv2nxZ3kwQRJ+HPI0n/os7g
9IXiHtVoK4GKEdQiUOOgvFxLxti9+ByFSl0bRMmzO4hxus+Uvi4vit6f7LZT8QGtGfgmCmH/AS35
ZzVjP2ALbEbZxrpOkSW08wzIM6Q+vnJbEIIxflzGQIa13HLMWRMSbK0J9hJ8cFVoqQYWCzPzIxgO
SPfNsjyZrdpdGmMoepFZTqIBafBBn5ocGKKW1IhJM1AtO+2ARxyypQjUasg0bVK6Pu2hz9Pp0L0m
yPZQuN01arcHAz8lSGwrYx7QH5ZPmXvD52GT6ILeRBPp5c1/W29bXwKVooQbF4Q2UQX5ZvEzptsD
7u4wlCWIMMI+bow9+iwBJqxmbfmqvho8czBFtRFd7bslc63r/UnkFCDpMZXHsfIRcIynKwYOLeEG
/3COpy71rJ69VZkumUrMo68TDssPqAY9UI9vSX5Uso1X/2mV2OSBhPUrzgBKotUgwcRfym6TApDJ
uCioBU3X8MSbS+QDVVtxP/TPev9YKCT4XWjQbJUS206Prrj/SzW99HYfUhgjnJZtztcpah+xJGRh
x13Ga7zEMHD2Atvh9d9Svgv2DurG5nOB+oC6oO4WDRmKCYCdQLxh65SvW+nrXa03D+hcas9Atico
bOAFcOzo3ScGGufnL4epJ1z0H3pVgfzklTu87vbRBS0yDuFTpRMSvxitDCtfTz2ZKgTKos8lBrS7
NBa9iWQg0thL4HVZCLj59EhoUbyCTtPV6KcuQ8wkQ9DUpDlcHFT64W34pfOXynw7DCpEEeMmxUy9
77m/tXWPPaguenyVwZY/pUYTJEA336DXedl5S5qSEK96Oo6gdLU+WMDZtyBGQ+qmh+WraMMC9oag
Vv/Hx+bwtmEei5dpDQ309+5JQ51z0gpvA+9wE3DXSiwzapd8NdsaB4D8xF43CdcIJvXFvGekudY/
sdOdIG6Q/hW6zEBKApylcII6hLPKqb/WuZx/oB5m7qkzyxLFaC9q+HCJ8crK/U5HnM9iQvwt9b1A
NSaZP2hiBLCw2IsK4b7CC+GV294IMjubciehP9PJV4bziWsyj+b6gLp27w8dqHVMcjOcHSz6nnww
ZxKkTWr6QMGC5EEXDPc4VYxsmFXEJVwvy5Jq3cpQLwtIIi5ZIhvfKVIsAmdbmetIC5mvO52V93D5
aAcmfw4GKMxA6nQnMfDEuN3LBwm24Oo74P+0mXAUDwZKSr6ecM39gsN02YA8GA8cNzLn0vqpDMi7
I4PJ/tHz+cvEO2bxYRt6+aB2kFL5Inb4SuVm4foa7fWfNEFieDe1wrDMR5gmP9sngkzLuVAU7RSy
KkMRN6KObG2uswkrZ0Q3/NOGPzzS38nhT5tWYfREhygDCm1Qe0OPW48tbpLGCpiX7qQoJEKin374
92nWlw15Fn4uMTk8ihNHuHJVMurl/21FxAMjRE7Oa3l2bcw9bd9a/Yd1frW3RYiOJZmygRj8wqoo
FYrQenK6DcBbcdhwvfxVbsNOr0EkzZZD5pKVDZsNKgDTLdiL/1rCsyBnMQogi81gEAkTje9PQP/v
60dNNGeUAB44WjjGbe8+q0dMf4ZeObFCmr4aOwJDEacjo7CVQ1k1sEJR9hG6mAsv9KOgu8w/LU9B
bW/t4gYShci4hLEt3XI+Ug4U8IL63rGluXxdh5BzCA4RfmtSG58JiDi4kGIe8z7SPb5WPOTj0AO4
hvR4RhXg7Sxup8N7nRB7FcsCu0b0x8+U1+7/c7bDGInFSw/BP/QpXvQ1KC7b75k/XnbAY/wdq54x
Zc3v9EwVEJvvTnPyjGzRJZBwVgU4anD20x4EQv9d/CVw90hhQiexD0D6vS/+f2PKtz8exaMwllEv
nBSEcg8o1UiRPSNOu5kb+jZrW9lYyxEAzjRaZc3JdWUEg3xc9sscvjJI8MxS3RzKLgmjpRorRU0l
1HIqPIQvK+J1B4d6QetnPCojo8701hHwV+76KKPmiGWEnAjjwAWNpSxyIVZzWN0kyOMm2hzDjw6h
FXh8Kjl0osXzuuXcuq0ybZU8QqNydoUsTbaDTMjVeZYaTwuk1706bBkoqGBOwv7U1tDAo5b6VlHJ
U9a0qNpbBuYIGGTro2vGjSrg4BKZ6fvOOhHAGkJ8z3sIjsGFEpmUGnjnB76wcG0/lH8xh1UiSMV+
MV3NjVoeNhn2rRIBG/oCG2jsIHeBpHjtH3RChVdS33459DVBHk6RoaeDh08w7U9vEtemj2No/ff+
Q9vvkuGjUg66by7Xphuk5Yv/pylicD2RunO0jq7PBxAcZN0VvI3Vg/lqt4DBiHVSgo1jDdHyHRAk
Ofv+0gRiBejqyPj4+LbtPSmw2iSKfh4/nNsaWqGey7k7i6pLSM4wG1h5VP+P8nGKwK2TkbEixMU2
p5fi++fVy1f7g6i8AyO+xpA6+zuyO/r48LQ7faA2lSpEN816EBmyQF1Eo/4x5TXyleOqhsjOQdSA
JVUihcWHH8Z0/QolASPcY5Mnyx5g8GC3rYSCnscbSjIFPvH56Hl7SMSUet4aJtABXoY3n22eJH7o
/ZSbz9DIFFl/h3wdOyc6ggv67gOqw38CEC3RqbGTTXHXJlHpvWX82mICu0DfjwHzblILmA715Vpb
3vKFx9cj1Z2gPTOyB2d9ljrpJ3st4jbUt4jP9rnG9UCrPzeV0fphmESIzsiBINFiUlBj40vMpoJg
n0tzItpGef3WRsZFwMbvXXEpl3zvVfOtOZl4U7Az3Ji6YgZ+syeyQ4S7N3FYCywm2xoiVe0JC4dR
IyLj99pgwhAq5Yo8vIVDhS0ZxgtuzPONUQzfXn/aMMPo9UJCMBMcur03hIL4AhXOCrTWOvOUdmQM
Lcq8IQXKmli7g8ahCpn8DQLrL0Jv3YSemq45+w47t/C9na8I2Dn5FXzKKvj3cLAcIua8AyTTbKbM
mnQaqF1TBmlt9ynvkc3Gg9qaw5LyE5jAWF5Yor03Xy2hbOoSF1mvlEHW4eCiWbu72m73ATErHzy3
doicUUA0toVVe5dws4DDnRZqmAi7unDW6x0LygJb2DlgxU9bX8CuO9APZjHEjnXlYWELWVzRHy6t
j8a8c5DAoEnoocW0qSlpnxCQq8m5ymxyVZ0QyI0sjzeH1OQpjBBm5Rxn/DJoJHUZgeezEUwdLUER
ZWy0rl7yIW+kNTaP0twtQYBeP5HznNlhGVHvuZ9JAr6e8WwxI3NhOP3CgqBRmQhstTAHdp7Ae3KH
e/NU11iXVuukmyq4SRYDuQ7lveQJ6CMPGdDi29j4L6uDdidOHIw46lmmqOdDEy0A6pP/Vlq7F2IW
gla6vW0EtsWWARaQObeCzd0OXh8yz8ebVOYoonVz3bxq6Dh1H7VaBIxYiYnelD3Rx1d+nsN6sHMQ
P/M5cQ92ZGmwYyn/WmhEcFCvHZql4EZwl2QuV0osQer4h9gzIlCRtGCCX9RTZmTkjaEP9PbKcuio
C0UBtcgWhb7Ck52e8KQPdd5UJHxkxmuhfc762E8JXKawAkBXV3lwhWk4nj9JwqAwMYSDOtypvFpR
jMZBMbNQP4x3/uz6N0pTB+a2FmKdFdWHNDKf1UXX0U9AxqnYmDPIDR6120zvs9D/c5wxtDtckiVY
YQe/eqNllap3jP5UVUie5T23O84bYtvHRtc+rS4mm76oASfMOW+Zq/bh5+0RbI3ql0Lm4qeAHxlS
GYZEOf6AGjSFkvyyLWh1udNyPBV+7Fpd55bXgIrdETGg6rDevV5w4HmytbPxOtnfGEbEj9X9lQrQ
F+t7/knzyy3aDJtH3x6I1xrIPwYMARSvlCcg9PtYUcPYT97t1fpS26a/x+a+ByuhOTLf6v4vB4OR
QO6kdL7RXo5AlUNfT6WO+xUmkb8VIvLBgPfilqXOATlFCcoRDnJIf8qBQJwH1u43ZlFX+mF5Diiu
7IZStp4fsZTJbCPVPVmzOjNxovs9iexsk4NV8DdUySlxxjat4ji2yJLVQ32j+lYuCSBBdec1Rhi+
bIaQKr7LjyEpcCwY5RCGHGI+w9GYoA2XCrPvo+Kj8vIyucg0J/Rt0V2kVvuDJNVkZTyVJpzCjzip
hkuGfp5pBqaX9t7ucCi+v2LNuZ9cQBYbpVHQDGikfiSdXTnyn40GLogSBTbjZVl4Xu4H65qKPHQ3
xCWFq6vSpaxc3imEb7oCkNdDbgaFJNG37EBzXpH/gt1s5rJwo9xpoCpO2dfvSUaqBE2QBN9arqvz
EI/plJc4Wa6JqijO3a/CzX0/mD8vbXylIw/kg5C27zqW0vHvNRl9LxljrFNK080KiEKnjnL1j2dE
IrVojl2AiAsU6opYMv9julPcK8wMAGK4rx1rU2Tzhcjymgg/dVXiVBzHCK+DhWbM1QE2iwR/y1e7
nPeJFVXfCDCQxmBVam93iHp1e5VWwT2lKnN4TP3bg+HfK/YEOqyhO8P1etn5H89julRh3mc9pKAD
CROKbtlDXiGLibAPutePSVGOR6nfXsA1f3sjk7x3oCcDS8KXUeUCWfrkVs++PJw5WjS2PkjmdSm9
CN1bwlLswYZQ0N1BcPKg4+5ucK4vqSkJOvcyJf/RMrazBwJyrga5rPu/vhxMXtt+MN2gaO4xyZa8
2Yj3J9Da6g/D/XdIix578N+NCpkTf5FOf9WlFAke/kJv5fXMhcWzKQ9WfVIVBbfussU1TrZBhm0K
SDlrWjkCFJt8TLB3v17XibktYm2pfXa00MGcErR0gPCaA6z2iNjnG5+AWlagT3tjRgMfq6bp9yOd
ev3iGxWGGIv0W2rCLNwLXTFJefKePx5281paYD5uVPWjRZIDKOOC+9dx32CmMQZKeqjSerZKoFnK
T8M7vJNi4SvvPaRGEUhmbhpxsJAFrK4K+ixukEhfrPiKrTjmY2euDVaxKUe1ZWcfCExlA5GbW/Xh
bTXLtt07dPliz8m+qpheAgqxVghwKMZ3WPWusvOva+YDmv20D71aeZI5SYOiA9VyrKT+ayBoVlF7
BP6HWQ549Mi1o8ZTf/9ZmBx9EwZNWCI/uVP+CokbiLgPN9uBXR++c+SdCZeG4ANyqWJpaq4nds4j
dwxANoS+AwS1+Hk2t/ERgdUwtGmrk2RWzdEePHPHqzV7QCA9YH4E1kl5PqF97hX4TmBUz7kCg/rq
rU8pp/+0HtF60yQ4lm00qly9gVWicCmHK/kHxptzVpsO0t5swbMApYKf0o+KqUmRcc7wV8LI6mvd
FeIwTYb6FHOjorelnKyhD1Z9ofH4TGL/lpo1A3OaWojrRZQQTwjcxmO5PDSaeXV0FozdwHpVpNk7
Tq2SpyVl7GfIFUrwgnC3kueULUEd3je/7LkGI38ECKdVgGWrOXqBhorf54cOIkATVkIIeGk4HEp8
AxPsOrbbMV1WnVsqdDWwueYC0FjNvkd6veWInr2KRaSS3bzcIx+FtJXhumqDuatvR5EUvywOtLnW
9k3PceXzcIEvXtwm/9wJBHWOVYBfwqt3ezMKftc62BO3coW4BoyABrDN2+EX6FYlgUfV/gZoMdWg
FTwk2Ftp5W/cOfWqnIsjUKvBlueVbv0D7lwxYXXCazJ85x9C7ybIi4A1atGUjiV6muexmAm6DYfV
wxMq2xaDbzZHhVLx74W6RD1kv+UBkkPUgAZnlvPH7vGUnxv0R+NTFLbzT4Jq/obewY0nYsN/r0r4
cHgYi1Y3h6Ya3OxYL5RV9gfZ/tEeWRtIb64+wWCLJrTIip2TP157sUd9VUlvrI9Ik1tj5dnekL7a
4vgwizmnRzpwyMvYeDOHA5uRK7MOqvApi1/hmTTll/W2Myr9Lt3nTAq7B1+T3KLhrgQKOCW5Eo7g
8bW75J/wa0ApCwZB+5Adyj1u0msBeoOl82gukBFQcBZzs4k1dFmSQwCJOpuZCpLu40IUEneMQ+v/
+mmtawbqJT7087QPfFfmv2Z/rX8Y4Ag6zcR1U14xQOXV0vNulGNWSYvQnerhNgsO2hwHB6ZQBYNH
j6vBUjMxMb159mmbBFWiCJv4MknCR3lm5LrM0QcyJVTQ7Y0eZTGGT6bJi+ZFcBx7QbopLEPW4Tzj
VCDyqKa508zbSYYXosAI1KzfrL7ouflvNdX6ckQISjZ8atozPvwzyyPzpkV5ZJKoyWEcthflGuNr
xZ3E9FRhUQGm4RsNFvdMMWHay3j0OC7TqQTeQammY9RcY0hPXQn57ujxccY8soz/vjanRkuxXd/L
YnWMTocgJQlX1Lj04btfeKfJzLawFr03gSLKo/3BnckXkRSfEUQmb7l72WXbA78mT4wADAv3TKIE
+sX7gRmmw4PnYGEz8ZRLrUDcmDM1y92ChSHm+P8nz5x6W9pCO9UmpwHRR5TDjFeQDO0fSaMtDqJR
8mB3LRxIdpnmNOG5/1kspum77S5Gga6bne5QM4OrUFD34pYEwAHBKvZuKo3nZ8s3Yi9aSsc5k9/O
DpTtfm5FtQFPGYqpuRGEpZ24mf9/PJPNIo/lbCD2HVkW4hoTW3JaWnjcoJklFaR3i5brbCNejibg
6L5mgp/Sy5pkAFtw1vPP81EwCeeQj+oQNe/NJbgzxcPK60IeB0sb0w/N+og/OTmHHJmFP+19V4p/
g529XjFGUyqaZHQvkE9joI7wy88fQMr0Hh5BwAWMrKLvbAdFIR8nRJ9tmRabGmjb8QoKKqm40W0b
Nrsc1DI2VQTOIBWLavKdmb/baUwL13qcbvq3vR6ShivQmc5dNl8qw5SpLGasF1vg4u7sxp+sfpT5
d8ifNyX18xLfy3qwmrhYUyyyJMDBHJIGWgs+3IZYs1te7OjqJMpoSLpzB3Y1K5iiB7FmGsTtHL/N
jun/Td4/oXbGk6m8/2llRXAfhIkcYpmDqS1mxXSAg2D6o58t5KjwqQoP9l6jv29393seGp8frwHh
VAmwAyUfVIsBaAG5VF4tobR8IO2vxeYeI3bRogbwW2nqgszGzBz5QclcHdFzwvTh8xGqCuEoI50u
wvzb0Z5+W4B/xH+jd79U7KKJml/CJPR/ikM4aSol2mbW7Sv1UcDCYzdCcnSy8aIyxcXWn+KK+0on
QGVMOD003ccezpzWKcsRWlqHu6pXrLDUD7yGUpzv9FHECQEW+Sc0XaIHMonbBvPH/Q0ZDAO42jUe
n3usNz+zoMp8B3wOlExp5WclxJ3r9BTgf8HY33UwJIA6Bz/QtJeIJ40FMVv/BpqvUuJZtLuqRLkk
wiB/6b2rdkNojRnecodyv67OosxJqVOTho7t8d0LPi2WyhX75FF/bVFy6/c5ba7DzuPTXcYa6yn6
PYeAOQjnXhu/T1cfuyUD9IEpD5guowk8IlYzxuYsERJqlbHDiCGEXbkLze7CgXAvGbJah3sF/PDI
leN73t3VA9qFQQkfk4NBihCBx5VJKFYDk9a1eq81RS9gWyynfxglWRw/3F3DziGIG4jcMDSpg1Mh
xxoptGK9y3mwh/cUS7XjfO1JsAZ8xgIgpVadLr39WEigRW2r/O/Roo9ZiQ+atAVHdcaP51bkD106
7xlsbwGTdLfsblOzJYKQ0s9mOesJbxHRGL6KFg0qHrNZzpReBmrh7loP3/wXnYfg8TLkiNVlDtse
3poOIlfTjL4oyj57G+kVQ5pfmGMnMkfbqiRNkA4pRISmoo/zl0/nOTYZQhI8jhIO6Wf01No4q82Q
I4gWV4Se5WA2yrMMlA+2HlfioLyitMXvIysYRK4w8UEboRslc4tfVp7pEMkkCgFssfdm+LyjqIdc
1/rEfQ9q4oi49HqGrYE8VJXVFWZeF9R1v+cE381nk/KQZOFmncSJJgWjOQt6mpUJhfKa0DqqtYNe
5IuHZq/Ohw7OXO3yXR8YKTnRz/zTVrw2jGtuPJGB96/G/j9uebjRxpbwE+FZsnG20vLIZIKQkh1B
bvhkzNClR8qlaMmADof/0xNCsElW1+em5KfEMBSltVNjYT0U3xtZf9kkjSG9s3NE2Skwhqda7GvY
8JP0vv+sdHXVQhh44DHQA/J/Qh3Me8aFIYpHX0eXVo05TQIDTqjOHlyBx/4GYpJAOpcR2V0JBiYe
7l3suniGkfn8WMNHbIPD8LZx3xNdmBT9HS9pqt4s1XwkMp4nTqCZa1hhDYvDaJsczn7yDR8sTxDh
2ifN145AW4Y50juYe8za9XZ3mJiEDPkhPdtRWkoQp5XaqX4c7kZo2pYZ54yFyaJEgccG1yqoEvQ5
prtbQMyq4AVlilrBpVgGgphscEmOWFprgkCRPuEpffR9OQ79VBkoK1SLDhHoIY7WlKKek80ArK2O
AiInYZyR+HzGkoO7bM53yOgXmQwaVoA3LsNCBlMGYBw38kGCF7h2DaWfkEdgSAPecMxRewUO0pBY
viWs2RoNZEMLbqv/qHhRp4ie6T7F77CZCKNf26/NNv/cBjkvzTbmzZGoPG966rzRLcDozKRDopJd
Cd0Qw1l1B+D7jvYjT+LQvBgKFkPf2AZfi25NKwO4VphTRDDV3KYPBWOQSNOasAhWRLFKknBHunIy
2i7WTVN677u5sgASlH2dw+/rAiXjbRBrRUWWsVP9+sMwwjtQVSBzungafMeSjlftP2PWSTnjK6ZN
39IucDU27RL6j/kDAmv1W2Q4chm0mWKPwddmheYIAxdUgNSEG2WTWo4Mn1neaekdeUO1qmwXQ0e4
ZSGRfLmMOi0Xj3zoUy9y9Un9II51WFhnDNbrk1TXh3PaV3jCMk97dyib6AGSzHI42E5pPtTDLmHp
V0reAbg9HCq8+q+2Eewn6eZ1dp+u53U8FVXRArv7jQRwiyTmTc6uYaLUtadWN4BB931rD6BWenrP
CPfIFxZv/sFHpeGZ9LUxC3n1KxJYRhPTy1VyxMwN09LJYlYJQz+XLHgb69Tlcp8sVI1tH8yZjVvY
x+Ig3amLUQV/T41ef0n956CRNhnqQg7fcawL2A9qChhFetaP81L//U8FfRmnQ/958y7WnDdQCUt6
47u8OEx5LavzIUufPn74orusMPGZOnW2YWTRlcoPjJ45I2hDpiiLQgCb6iY7y4URG90VzfBNBdzL
cAxeFS3lQglap5idBw+j5tyCfX2Swq3zS1d4QKBqZxyRCx8fsdSPMIUroXbPAhDlpuVJWILIS2/g
oIl/gHQ56f1eGF155Bh8lBBjimEqTjuOWfwj9yq+e0HkRLF/iz6gnGGkVGVQwz359+k8AbpLMm2B
XDd4dgEeRPEqe3A6RuseFO6KLE0BTnum91XrubxMrnoVdUvjK9IDTsNTxj8AoNtf/ey3jMeFjKN0
593FHPG7Y4qAkaae5KGthQLemX6tg0PZp2eNOX+IXIUfhCYY4igM7ASzQw5suiHXRCgglMlzR2mM
5eXaYuUglATt8Ha/X18iPVZEEinOXS1rJmHD5Iqa80Vn05E1NZk46Qw5ml6PDsH179f9/bdF0UTt
s3RLESp297QNmxhwCqWG4z2bKtLnv1erohbM9dDDLku6b+gt4zcKDg/sNiyUoDQPgvEp3xYRV01E
9AxxqGG63VCJzGh+VRGCnxqjmI2ljTHLEVDugQxTcs22EXh7BLk8YjZMbPocIrpIs0FIUNXW4UNo
oAXGX5BRm8Jq2738Pm7hazdfPVtc+3n5sjmTmJ17huj78b6PZjaOJmBS81InTe/AagKT8t3Ogpbv
6mI+8iYbKbzkSK7OvJ3TSSO7RsvOAEtwwaBd9ebugG+tkE8bBx7zy4DDbG+hMFIa8ObxxE5xQ9Xr
4orghKx2kiORj2yu95NfjFKfENxdJGOtfwoBtyORkztiZGTIr729fV7LZ6OEZG46Mz/JpOIerhsW
TJBtMvwlZ1thb7TsgBZ/QihLNxI1cwjxDLEpLazkcR1ccLyG/4oIXjsqu2EtjbOmFDqdMBkUbNgf
jgyFhh4WPw5dFzM2P7BGHtnn88aGefCe8F9BdTQ9Ob9OpkxNzuTSUdYvV41rYaaVtpssWaRFty6t
jFz3ibgeJ2KO6q28gKdCQXERi+1q2/0t6cB/+q3utttU9W5gs0gpU2VbviSw5InC7hCDX0f/tu3T
76ta5AhPeg8dOY1OFK25AFd0zKXaH9EPljEwjP7VsEd6WbFgXm996K4FtGuFX+ey9Mw6sszeMGLz
1lVj+TFfPIKShgRsrufRr6+ZPCLekNnb+5hV3wcGD7pZClXO2aYbOaWls3JbTupyFvtQMo1nsosm
lXfjDRIljodsYmmxhb/DgDqBNLzFhMq+ba8IrCYLehS1Yl41W0jQkVV6UXSNcnVFwU0k2z01YFyf
ksDT65vOzQRXrMGwpUgnvFnRcYGaunb2Qkb+a18pQAlZEHn9SpKXu1NK72TlN9hSJakzafy0Gb/x
Klq0zy2c6IQ/DawiORKsGgp4r05iVHMP0Y6Qr1Kc5aCaTF67J+UhAT1wPyACjg4c5Z1fJO73DTBf
T6VHTCJLmrepq8mYoRZrBeRoVMGa8MEcH8sv458JlOfrTNWSWfZl//ntBVarWTXyPxYreXaUlirN
KLLRaQ66Fg7+EMumOUOsHqujiFOWu7cJ5xz2dwih0l4QpIuLPAlQCHVZ6ZM7Wq8BcpFSsH0Bgq4k
QsAeTPpz4eLPQRu1nxc+NCJqO1psSiZDzwv7r9GhvDUkp4nLgfI5Ukvhf1bx7zZMG+3VOpFLvcj/
CCBHZVADNShiF6hY8SHc3yI52A1PL6BCqWCBLrIfjZze6WiQLxQQznH7hkwK4NnCTTvH1gkB/uf2
hXxWFc4Vhch+GOv99sgKSwKvjrb1mki7HQcZ4uAQsekaLkifrI5JXU2G2Bp8DPzfB93wmlzV6VFM
5srUd/ptF7CBR65bqjQVnfQfI+hpIF/ooyPw5uM9wZ0ZFICD1tMXBlm+mOKI1jP3wP7Svjr1FKBe
oCNkgbrA70Ll0ijSyYO6GxDxu1d/RcyUDUhkUBS8a1Zu9n7LP3Aju0UNh6LD/NAYpDZCeV/hKdSy
2GNHslM+DR3fDR7aa5C8kGGk+m9VdBRlyx+h9879Q7E0uzbH5w+q1WCEIpJXwtTpIDSwu2ITKRb0
MAH51rnr9P42vDCqpZwyIMajg0s4f6YUpyzn9eQKASWFXXizNvxjVdqnV1bQ5FXFzT3QAKDaAAG9
AviWROnN5mx/EXm0E95rdFDovLMjNUWVUXeIONVxeakCD3Q0ud/DhQpX0fwe2+kY1dhj2vtCix1a
yYcAwY2Fcn9+YYAZygvkyRTMYI2mXs8LbOU+o8K+pOE6DZvvQF8wJIxa/hk4TIhc87CPvP4DUEg7
uxnvvY6rrdOODToSrn65FR+/sldEsKtvIHOczxrOyt9jcjBvWhkG6QYyoDs5KMBlONRsuj98uuR/
rUhpyKOtp+rFaUP+YGDiotYueSdX1l3Y1DnNoWFDf3ZYiT+rHXNW3EsM/ZX13X7tSRF9ditf8KAK
rNsGALAY1tFU7BrYxYJxu+Mh3/ff/iJCS7vLwLYiQIz3thw/4HxB0uAFcGHDWbMGYWU2ATYvuyZ4
37AhmRBLtre5FVuJAVE8ukPYSrJXuNe7CxRk2wIq0fP5StZPBW/t9wGaQ0rjMZXPEhOiMFYA3otM
jPFNaNaAfitK7dZv7OTuc95ke+HsA7wCBZ2pKjLdsVoi4JFEMZc43pEFG/KhC/icmS1Ci/hfBxSa
zQhJTob7JSQm8H+4mAJxn0nXtgT8nuK/P+1P5zejCqlTDA5nb3spZ/G4ltg/o/EozOeHuziVgkQ6
zZIE4TSvOiQo29++2H9dD4S7gEUhyuoFVsw4aLMEGUm9RDg1dZD7awGotJny8kLNoVer8GXsnjiK
tRzW69yasRJ0wpXQMEGI+WNesUrI1fHm/tgYN8oBoeagNIXM/9H+hfgxvABTZO7YCiv15wSZI6Dy
0w0onvZD+W6q1e2VUvXpZqA/3DBm2SOYacGlhihTAwD9h5QdQW5o4RfcjIT7eWfJXACYvRHco6j1
khKsDgGPOgEyED+MMooHoRonm0kyuo5eIfWAwQMzzZwQT/1ByrX5Nxa7vetAFREPTnoU5KNhm1Af
+NuVQ1eeA4wC8H0iFTtPCUsFLjJRpbhpDttcyCx112bgK7OVAgJeGOXrKSFDrlwUlAvilPtCesp9
nLTlvecbr6Ag7G3urt7li9BdOrDuD5AAwb5W+tPLHAt6Fc41bah89x/QjAWqTmRJnj/ZiqU+K0RT
c4T6CxsbWdUNMi0vfRYwVxeIhZ5tnDCqUw01cGT2FMHMFgCkW57wpB/qhYLXON6hjx87bH423Tkq
nJHkbo5DyuLlzc9Qr3NdLHnElQFOm8PT4qrHEMALjYAiJd8bQcyQ61noKgjVGQWtX1Zpq/qP5TCw
BSA1jN59iNPXmZw+I4gSCz24sd0ldjThVlMR732vNK7tmXGvcN3U6977fwsCNVPQo3Ddiw/uhFxB
kE45t6ibBvC4YInyZu1gJ26CzLHyZu/8rEkS+mk9uHBtweazWLw6U4Tto8O73jOIS6rLBRpS6+5i
RLvMxt4ocFt9rdZ5VT9/Tk6fhkxzro6IzF33DyjS3K/vQE2pX4OTUAo4hzYM1GWqHl9iLF1wbk8A
s8jPus80/cADpuVt2OQcBq0UMqRsDD7KQ4tsfl1tu+gysfoR2EmStI2PeKfgCRfIik5fFjoObz76
AUH6irTZX+LrFJO+C2Dn40o2JLYvLbVM7745B7M128ceKlnVA6/tL2uKCcAYgKo8NNqsAibZn2ZG
L/U/fRdvhjvPXYEYbmCpkVe+EksXWZVD7Xadcx8f22PmaJOPWzYMUrWEAUFVznQqN7scRjSq43HE
JVKffplNbSnmDzWm1MyxddxddyFr4DYoDoE1qzF0Y46NOFkQjh24YGL1+S8B4PwC8QXyccVKRdlC
CAg7InML1WuwYZETID0jZunJXNIonSs2/DQT607cKOJUxXaAhdFO64ruXpURn4LowjJAp8tm3BRi
sTBCpAsjaGnyCl6KdMUeCH/0H5yrGzrlLkkd9VIxWrlMldXHjf3Anu394ooz1zPes9y1SHYhbxRU
2VYKOd6jStA584EEBdpSfi3R53D5p+AL1optX9wlqI47V5sZ9eRkeeQkZJDA+WFjauGotpUQsj0u
FuZ2jFj57+p/LM3o/0xeGeQnGgRCTwLU5UUwfOLlUi7cb0a7zr4BYEreGA7n51Lx+wn5Hm4cqABm
pMNxouIdbPomPOwHb5g/1Gs9FZHcvepfiBIHhzpeVtcv8REVTAaMOoeL+HPVPgoPircqypghGMqc
bnftKgYo4I2c8IxXWJ+RczmwTFwAbD2eLqxQzsiFX7AEPdhHZ2ccOtJjOrME6XfRHKMVZ/lGTuW3
DzQZpQdN1ZNV0Px+C92xWA1PHrGsest0ZGOWN0nvYSMP7I2eOnKazstIFavcdnlBD+oUdEsQeEyF
WSJYspSuOtOyEJBHUjPlSFiW9K+BqoZGy+WXR2hy74shEbzH4sQbbfw9TD5suPrGpEvI/8ieqUR9
chpC0+FOZWHYhCpDs7561tVT+NYgbfM25AwoK9fK33eYTaHD8uDhVSSaRyv8lsuFi3kQ7NWiNBEt
cUvvMPBaZSeSx449bhjPxheFZZhKhqGmwLZrcdugh2N2oOkOa1x9/hvpPFxQz/vmdhpweBzijHpn
OlZ+phDAZE5bXosG5uVhWQ0+GgEGrL5iumCioFbvTNOtWd7ZRKaQG4WVDs+XIVBaFI++xmGyLdm2
q89PvmExOkBSwFHmQmdvCPrqrLOHXJgiU9RA1Q7PINYMbSAl4+n988YQDaCKUfd5l4P1yaT9QiSo
XQoeGOsMN30+GDyIdgM3jcrBN+sdrvL6/X2cYs1LaxxthoRD5/6bS/cFqbtkjEiZsBCHdZkS5MdO
9Um9O8Im7nvZJUYTaUkd95wT2ujJMUlruQkvo3bqHPlIASpPhV0DVdsBVepX9XcFCaHUbR6md3TC
J/YLo8cKNqVO2LAvzdt5g25k2Af8ATGqX0XSie8tEJqRcJ5gyXeGk/1WZvtweLN6uJHx2+pFw/Nl
lSIJR4neVX0sful6ZcYEKy+3QZaZoTlsmrUAj9I0RuOnfrv51JYXtn/zDyR9f1V5nufbN40rROQ2
8dK6vWIn0qGkIOFySGW5Gq5W5sIkDy9KRNIV5gKcq/2aNq06+y4U6WwgOpINT9Px39so6hQEVVI4
Vthq63jRtNleLC9wwmSRShlRkpPZKTQ/pxCrMKVbo7cbQts8fMRDF7KAt83caD8XMG6Rj+GYpyAW
1VNuTOpB8+Qnp1tjaAqL6avLHOa0DFmfyvFYxkwrKDUtIeR8G6G+7GwLH6BIELC1R2vGKB8msW0e
WtyviupdCyBxeRMSNYu3rjLdzdVj4NpeqzIKvOAfT5WbgGjYi2QUMfn/SjskG3NluJ+6DTRXEVck
+/9AEMqKLViZBevGRkdy5bdJrhux8/b3FCaA4m7sXtf5feDybiYVH9OLcxuTEoIQHuZzxpgBeTVx
rLQgvJnJ3eMPjfaGN8yUqERH2GxLb5YkqcXGBGbgGaLL/WcT0fJxV5w3OIBFUXWPB2XBvUUKcjPG
2cRXk1nwfTTYha60iV+c0v/vd5WKKlFehC/dstDn5l8Q5HKp7dgciPnHw+jnCKiJ6Kxv99yGt78K
KISPw3N11X0F2goHBikPePP4NEht9VXUnJfweJUhvB9jdAuGd8j0e/EqgNDH1AIUnXAF+KCVOzVw
uwcpGJuHbx4e78MvA/kK0oL6ZgKU7ZdAia7nSt7svszxxHQxT/EIm2mFl0P8UTEwwFu4RYXtVTZ4
iDG8UV6p7n09h/TajPtjr6MyXY5i7BU2iMdO4+VZUUJm8n0XvP1X+mcwM2FH58M/EapLGyjAVvao
tugaV7PkvusaF3qlizcISpCkWET3GCRV9Bh2a0DeAnjlFo/oyX8nZ2uk8/x917LZ3b3CBIbLfLAX
KaYf5oYpUSpanAq6pun77eBMzFl8CaJdjm4UP0wuNgHgQO3+N30N4D5ymy2B9o9rCnMYqJeXmNLr
2M2mU3XJ5jgjM7PfVS8hpEomzBGnuTGzo7XoO9/VY82lFzuA23HL/eBZcvkeO3CPd2fh2hJ8Slls
hHceFGvRwoy+QeOoA3IaHys0MhZR4+4s3FQwhjWP/GLkrgPUqQqgG3Z9bJ5BgXEb9HpRVlfVB9Ef
mvo5ghxW7aGnoqpw9uSROQqPjKc9LYRIjDhpuacVxmk3no2Kn6yB4FUZt9wCLc7fdxjgEr9CYcuE
GHqtE5EZdkmIGf66cnYBLM/l+TXsqXCvgpA6lsDhxItgcPg5Ki15W29uS0Yg+NT5Lxl7dqd8J0+r
5heha5+Au/ChWrAZBYMbaKRQriu3/CrBaj6DsbUYR2qznqqqmIUojVAgSyuoCdkbOTugoWytkgZY
EQfRy1yD2KcxYABCjOrhhFB40hHq+tG1TatoTohcLK6nzCiM0yzzGgXPLpIyK19B/PMaUZIJ8ZeR
/6FZRX+W2ggbIX6omceR2MPmpNXRGmRYFiuI51D1hIRww6Rm7OMU6WJH1w5e8P/+TzIKQ6x2UiqW
H5YBUZCB9VyEpF5rWmvA2yzZObUs2YqUdnx8+cSSurLWzj8Uy7lf2uD8xL0MNJnBEERuTn2s9ScJ
HXEhVimMgS/U9ekPj7qaZALzT9S/TaVRXue8/v7+FzPo/cBBGu2i+d+rdqbPWVvNQ6kqVq/KIrPK
Del0qU5nP3Dj8pWoerbq2V/ypVS0JFA1kL4pMVPyuyCaxyx2gqBSxqNOZ9COcdKVgUBDnmvf0Zlp
dq1hitLJ+m59SgL8mNxRt5szwMm+6EoHc+sJbrKXG/BPW6oVJUeWczZkVOJ9UKdm8hxmoiaDbwpB
gutFC8yDsLunNFTqwg7Kot4U7HO5gvYGAHvFZIyf05ldn3PIT+zeIG03BywtCuSXrEYhkJ4RI0PQ
lFj0JGo4pLAtOgSzqbQuOB89qS6AGmKzdWnOOloOhIl3eWcanZATEwztWlLcgeOcRddRch68Vksg
s0S5w2HeK8fJjAAvfqvlOPTdo11pOcJFK5gSk+LfqVmvb6815Xhq8gReePLOX7rmwmwIixpoh2d8
b1eQk1vCqIGpkP+fAzA9qc5wFGeYGYZSk8oOiZMrKtyjaKQmOJB+D/0UThsTSzO1AujpXbzefmlM
u/wA53kuo4Gg+alttWqXYxLfQfAdaHh5N3vYxTzb+IE9VSBftrNVwikhuBrd16OwU1auKFz1SOWI
vSvKyiBVzbqKBoUr+pWuapVjH+21YygQfmGpIBjUxUxOtw/vENUOBXxvJnQ5wlSB+pChmO1vXVlB
2J3qQRLw+g8uZkQ7UryepS87vLzk3yIITUFWR2JhvOTOkXd8eDVYxUFAwtTGvg2aHyVNgKsLvQg0
CBHU0AkOLsJ9qG6KKl8T8Yw2svA6XfV7pInY3YUCKovlBM2cSIAMbTPtJJ7wTaxsinGu8hKrBS3e
pCVqs9DexzJwO6LTndPZ713iKL3m5trXvbJzABJJdP61dEM+It+3fhVsPOAI3aAifyRcieLwx9MJ
svLB3cjsY8JyJRBoD8kqEcLE2sI8jCQpHZMMgRnmDMaWMNsH9YWV7GTqBcDMFfP3i3Cl8bfSvoKs
wBuruQgLihRspxR6yUZvlEMSrjFdtjsUPAXE/+67TH6fgfvRggP/Dj3vWfOOs5raEnV1Doep962S
+Lmx7GceG8aigtHRL/BjVdV1IDweijE/9jmKVv2u0wWWyQnzBpeJBinvqyJeAMBAoXaDeqE/asV3
Iq3sCefYz4dzy91lGfjFNN6RYryEL8CBaoGRHCXx+dCMvfz9pnYnrkEWhCuLIePzT6+aqXxVCrfQ
q9pi4Ae9Im3fcg/n59kAUKRL/6l6vJXC6kjiDhG1V8Otyz9DFY4nZL+4bx96Fs54L4Aai25/50c5
+aomOdFbGbJwmcpF9z0iO2/3xDOXzJj1AXe41Tsf8MqPHroRrn+eX57Zx94bdEXVrCj7kwDzzlQX
3U1es7235F3Bl+IpH/ugXnGOiVK+5MLeRDnP0iOt6FcUXtpafmcAr3HcKI7ld1JgDSOPEP2ZgvsL
aopXrc/O00FTI3hQDDZDivr1tLP6ZjgQBw2t9dN8Vy9IxbBMO1jgly9iBD0VNIn8MG7BmOGNNwWN
4T74La9AXBKdfDjGZXBYM4CtzhdtaBdEHtIeEbaBRzFmNj53uRgpG/e5HOn/b5SzAGMTPRHUbpSv
n9+U8RlJxeuWehORBmCewxD27XxMVYI0WlvQ5NRSkZZrP0AMHr+jvpY5W8nYOomu1veos3MpjvLo
jONTVB3SRpsbYcqcBJ0ckNL5dY3807yvQMn90lwqvBNz7dGPM/CZzt7GxM+pVSjUo37hZmL4AL9g
d+7M7v4+hnnpbaVMj14h+gWNaREqWfnuQXQtUXrVYkBLvdsrPbxx44FDXgqtCiGNTOiaHjMAnz+u
HvryZ0+HDXkTvHXSQayJKmmhhXcQk3jTqpSp/fCPxvp7qMelvZgcnwN/jdSXRn/voODKcZSLILAm
CxDeFSFb0bs8MOpc2EoudT/WvGNUH7CQMB6LHejQQIIM/bhEkZUF5XtR7fJJyRqBISnZNlVjQW1R
8IXCHT/o6ylumXnXhzUetRgK3R1ZptXSuHCVnQ5FKN3GcyuXOf6bGScwjTkgR2V31mdU5+kw04pz
u3FpInck3MbysN28JawzXEiOvsdXznC5HjGf30tAJ8e7eGbeMoWZZSq1MDHu7zwIBSw5JDZJP+rJ
A6X3g9oHJ3QGj6KWmI/+sclG4G34O4/oG1lecv8Y1Ws/524F45OEVRwZl1V3sZ6JnxeX30njyfmL
Stbt0k8BepTk/mHIRmhnWYSDGbDQw9ouZ5Fcv+3hDTHcUN8PuiOitsDp5TN1xca3nq15PKNqXF6K
p2JSGNC9JHWdUxO4RQ81jYL8yIk+ea4suvWcAL/GBDiyV0VH68yZCDRzJ+tJm0rZXlWwm5G4xV6Q
trPr7rbsOXL28zEEnbVb8xE+cVWvgeVx919UlpviOV8wfdY57knNGPCfwRebMKsKDAkfWyxNhZdU
bkdRXSM45dLWUjL3U+tzYVAQyEXJEIvRS6U5kIKTl34LyZbZ4uFa6lm4HedEIvhxCBHMaAuQ6WVp
PVRVz8lA42G9D32XzSUWN47a52JUGgIa4uCAggroG9Xy7OoUbWeJ7d9iIkvPerX+h6D7A94nezS/
g0z93NzVahCebI+30A9IDiCzpRY0YK1m9SxDhcnnBY8mzZ3zX3sRcCkuIx8MEfKRXWBftN/v7yuR
+GD4DjxRll0rrFsasnqBhmAP0PLB3k0Iq3LnTcR4Us2tESlF/USm67XuIfst4LZYwO57KEVHH7xA
fbAhvmbuER6FlzrWo5XkZGugN7BousJkGteos4jsYlc4ETVYxqxPZCQcY8v4JnIPdfqFJm8990co
o7zqCSX3v0DNG5XZK0b8Vv6l25i4Z3rcbyZ7RK4JV+7uHYscc+TfnjR97dxwrOseBvt9B6AgNUS0
Lbhsl1X1RVKpCR2pPt0uMS9I9F3Qya4305DINYXfsAt/3Ncnw6uy+rS2G4O8L/ziZ00OJu3E4GGr
siyYWurWvoxnzdWXI9K+zd8afTBSOkry17gTGF5gifXRibr8oN+Da8xuDdoIwbB4rn7V+M6YQkhr
4Ex0Gt7XOYm58RbsM+q9YHVnlnDV2/3BR8JICq6NHOpZsLseBuP0PvSYtn6MtAXOUBL6IMOEadqi
wV8bv+Ib7EvbVCrjuKlHP9n/IvtwAnEHvvCNcFJvE8bulQEY2vrZSwRKQnBPs5SuNm/pBjyUyTrw
mBYTvK//9L6AV6eE/DtGqfq4ekefHbAx5DTd1uDzAAsCtNBz6oozx+cKYZeG0JBsnX9eowIFjhrE
zaHk7SYek/S98/yr/qZlAU52H7l7XAfalTgKx35xYILKAaZ63nz51ejcJfR9VDjJbq0H6ye8yWLA
MPVLjxRPkJjpfcT5a8ZLpvIclHtFZseUym3DQXnuFpr5kQsfxxMYsJTUaGJ49Wqi2XlEGxZ+giVu
P+RUxfRKZat6YzHHyzMnbCu42rDa2wckv3ShLYNlSN1nUsM8eOkQF/qPnuD5BPB7Zrdvrf2OkC03
pTvU8yni6mKKxH0OhyecYaJE3zTNQwwk4Y+MrSJdvvlbNmrt5giH7cSUglbCg4sRLvPxalXnGA4M
6c8LrML3HYHN2k69LNdKaaGdYI4+i1jtY0xkpDijMzaOkMCO1H0z6p2bcGcg7vJNBJaF9dzJSPqP
kNRwimPluspo7G08FJNBr7yWLqa6LZK3+ZU3TRf7ILGkv5ldeu/NEjwOOd5LVsm7q8JzFnPNS0l/
Lcf0gXJ3hbaNj0s6/3+drQ/axa+FFlZF8Aqfxg+kP4XZMgpjXff1YOh2kWGAfjrVRXRzRRdSgesu
w+mWmV2LBkr8abBulzQhM2P7HCM2LobD/c/Lq4cVUXebXu9CMCteAI4OxQggfXdZX4eyraBWLrO/
7eYN4oxu6/nrCnWSb6utcT4BWdIkrLEZsDRWiQ+IPiMNqdOWczJ1a11I87ZaxzLqqjYS8EQO2hfw
L60+6Qn8RIumUUpIPnjZAzHSLV3P39Kz/jg1bBkSWFCT5Rx1rg3YEmA22EBvdi7Qdq+d5s4AFt6L
Rg3gwURmOjVtG9P37tzCuZOJ+9ExVSylnbjETIc9PGjnJqTeBDMzqUYqLz+PV/Ov6U57TvhFyv4g
n9MwNF80D2JkAnAMjfHoyLBHifj15n06ckokdKltUqkz4wOoXlVfDGiDHzumnNX42nL5ADsx+DrC
b3ShPIGmiHN1R0NU/tyQPXglKJvIMZtHDGk5UTuFn9N8UFfL0CyYOREb0Nv+5xT215r5fwpbvZRW
b3t1rxMzJn0WVR9lpQ9dkd5ie2um7Jwim3r5eO7DnyJK/JDjx5bvqdJeIquXBxhy7GZ1CPC3Imcb
fkD6Q0s+hGadvOw7Hj0gnzBjCaK5GikquJs0ktW9ZCAr3m0wZZb6YCVsBbDrG01sll/j5ykCdLeU
Bcgu+0tBwZLXeYTZOtKfFJduOxHtgbmcZuY9du8LfnyUhJLwh2DFR3N3hXoFkgKhmJUQ/1RXtsKj
k7kazAV3Vk2QkBaw+nRYIgeXcVjePmfyUrpaLC8nZCIgXWYKKamQbwZ0G4idCp7x7ABGomn9f/Zi
p5DBKskxDni5aOkhfqpO39j9UH1ZoL3T2JjQUD6Z7Rd6qau8jFXYCotsO8wSJZysrAkm82Dqk0yc
K369esFLYYoNEn72BrZ+RSVWsJ+fHVsx1bBIKe0pRepMt76t1Fnyo0TQxh350gkYDQAy5dmjFcdc
KhP2/s38HqfCbc8vsxjg8St7/N13GOcXpzXkcVx8c9qq3U9uPZJh3N+AGnncUahC8nlXVtdTxAFx
mJyAlXFu62uH406HewEHCfWc/apOQ0LT0Nb8ZAxjnWqwBvX66Wb4aY26NJRpRciCIJjIZBJOOpX1
LYrVaachmCLJs3aPlYiz7gM+n9d0hjzpOYKGzqvRAnFJOJ+eZQ4xiOICxwIuyxHLCVtXBnQhk0fv
PX9TNYRyWqOv8or67CmZn+r5smdcaivKNdA7Wos1uJSziu5RlqZUWf9+/CY6OIq2B35YbBveGrSn
tQxIMoTmjAoLtLHn1GaxZsrflvHu1aUVGcbsCbTH4JLfcYeuLaLh7ldQznHpU8CqlEik6jp/FwSK
CYEQQOlciA23DhU8uluh8gIfEJcU/G9MCj3K4Cge98df1mu0EAXiLCb9fDZ8l6CmG3efWLzFkSCt
fGDn4CEaGG4oy8b8JPkineuSce1z9Bkmktr6xrYeaQOAALgleiTbE7foM1Uxw+s+Qz8Zdz8tlFJO
tL942V3sWWvBA0GybMifefRpvf/5GYt/BwV2nhJx/5iilQCBWkG4VVRKU1ScmHvarKKbypR4d1Yh
/+303wWVJ7k5sX3Qqw0DO5qMjVJC9698mxdfzYTcFzw65SnFXYCNBbDHFA5xRld0K5qxA6cgKJPM
f/kBc/lKgHglifRv6/kZ/llYHptZbJYLmBVjBQVrtyuzP1sx+WOhIXJlH6tiV307x/HV8zbp/DIZ
7JfNF/CXLuLTQlEHZn7wPAs12k7wyBRMofM6S0jRjd9gkJF5u8tTA9RsjZzAfHxZkbtUM1rhs0DE
6i/JfdY5ox52GonIy/QXCY2Z3K1fC/FIAM7rWpA4oyPbc547cU/Qf2tz4/oEeafoegU2FE+7qI3Y
fTBTXJ9vN43sLZdcUdNO1n35U1kAYvo3y001RMMnnIKmVDMJ3yD5KR3itpGkBn+X1k0VpYDf3gRj
EYLen6BNtVzfNEq+kg/v5AP8nNzKwUYuQAMhqEItbRR7XOR6pplAhk1scr3hnhGy2MscKwtrh4sz
ME5ROEHOdX5UiMAyTbrcvG4rTd/Ig22i5640Juh7yevNmu3NwZ89o9QrLN48xfF/Zh5NP+OewaoO
sky7l2FILhHD/6w9S/92LQjPRmAQkkJKYJu154P4L+bFLPDoZudglWzAgV6HYJw8rgHAZO+AVaHK
bqwvwYQk1HlrcmCNcUHYHnSOvpdE0ZpuOcA0eWEQcmfJX9k8j628lSq7ZJ+X8xZSQrFMltwyTPVU
sgaGl2AT6fAzd/rpBsBdDrhvFLWkOXMPlaZJVLp/uh7j+47nBOPp8VYdydKHnKNtohqEQ6qfgSbN
h6AjIjR5KkXPq4Ts2O4rGRio4HxKi3i4n3OEfoLWCHD6Z5luasG4Q0YiaRgNcdwTFChHmLp8QJYm
2Abbxw1k56UjxXfvBY0wzuAfGGJGDsW99juz8hGg7A710ZEH5zoknuc4QrbjAIUo3asJUlzm+Y9C
Ud+O0z7hIXNiTh0uPmxukFAX9gCFmbvobuGsqdocbB8WvBNP0JhX9kHJ+VwQGALSMhDIV6uAFWkq
c6S0xnh0xbIM4Ax1B9oYzzig4Z+irfOJtjcPXBPCb+kkzUBQoiRO35dgZwj8+vVWG1DX04Pjzyni
3aiHpCvBG/cTdmevaE6FZsxQ7gPyUDUCgwAowneOCXGajEKjtyKwgs/Xb3Dvb6UPF8HMyNpLT0tQ
mNINV0x7qmopCOC5wLP9pseKQnLjuXP/CGxWKISVarJgbb/VC9QwoOWtWSNFIDko8XODkyKITT3P
49L2pJEMUipbTPv3/O0iyPPi44k202UkT1//xtOMXQzQAZXYdJRekoC2Gli8e4jTiwwLs8pJ2WJh
95DpUm+OVp77cf4kxK7Oki4zmRBoSymPtK7C1n6TlmBQuij/pthlxM/4aHHhS6OgoFL1rd7qxJYE
IQG7F+flL+HFoyIT1y0RD079zCN5ZarML7kNDlyQUpAS/Ow7N/1RTlCQeL3U4h5fr499Jtux6KIA
AtX3YvtOZpbq06vL4dHzzIZ2/4TUoHDMLJK3g3HBktcSosl1ZHaVpq6fLIWrDGfy6wWXsaTZGLAF
Bhbn2FdLxY1jIt4rDF0/v0GngmrrxRg3XBNdpwjxOGU3LuE11MRqnsCTzpSSh4c84LY2QvUXdsI7
jwlBXyNwjr0YPtJ664HURvfOCm0z+D3uTb3x5yMg8AtHtvyWCIOQ6tChUqIMTpz2uaJjxmFe+e67
gcpyzZ00y7M4mIrJyPKU6vYqCtuk3oUR7ynAURVRlajooEHD2+Q+xn9jsZKFEVCslUue2mFUHvcM
mg18iqtW4BF6E1RfS2UqDxdpmCa976r8QHgxbBwUyh+ISY8VI/+bxUg6LH6EOL/eDHzTHswCU1Ua
NPwCcPkIKXvsMjclUXBsJmqqWcbgdotPnti7+qgCk0/LQ4MVBtalO5zFwUAMC5s5/zarPkqEhvSy
yWD5I6QcFnqqZTWhG7Hyh4triVJlIVBIG8j8TsaPNr0v1yk/R/gYSDdFd4Umecc/RM8LjCNlRuYj
0F70+YlzJ9SS2/AVy5ZAG+YLJZG1Efgk+Q4MzvPt6HZfJ5XVuanr1RMJ3001mJaEIdr7F7B54QSg
yy1DahMY6s3UcUrJZCHOWwRuRfWsY9/ExU6CG53YSrNi7mJZaKPTJf0TtXREwAr6/3QoECog2sSi
8N/Y688zz3qUA/WJVzPLExBGo+6+8tN7Ng0xbmgD/jpri/hwrmbMgxiFEKxx2YijWG79hYUaqnBR
zATTcICMIr7VwpCgokNIM3BDFxuo3ZnLUh4AM3MuT7MFrYmENRLMHAD+I8BetkURovczlw9OekAd
8K38GGDSoliHsAAIUmETmP+e4OYik+4LHYUTYs08qAxKDsr/a6pUPSJjMQearolQgfW/wnh8DCvT
NBAqrbfDDU0bI68cBnZsRHnAYtl5MItwJXL+5e1kaGS4nM/Qg4OwLChMvAZ2k1xazIIITIP/d/z3
iLgBzvyCr34x7bdJmk+5XjmDtdPWxIWmPIEu7uOm50QOL0q19g/qR6y7eL+G1txvrvWoYAVJrq5B
Po8V4RxFQE60Vh3pntewWMPrhphboaHMM9wEBFHRn/sAly9/NVQZs3mWB+X9AVI8PtDcSJV/aJq5
MQsqmlC5IR8OSKrdERptWre/ydfqA/bmP7tsMmTN+J5jiHq3ll5AijiPB7SlP3E3GAoX/Vzv2/o5
VCpSWH1ylIbxRUDTM2ufACe2yjtlHfYsRjkEAJvduZ+N0CcrHIvCy7YQdmc3umkY1lsao5KUsAVo
ZhHmDt+NiSQ06SdSwbDovcxO9dlcCTOLtpPOMdbxLPBicuf3qwY6garNMqzzj5GQy1zrnL2209mV
+o4vocLLUZyGH310XsH+CkepILSe8Ydf84Rqa/7Lo1zMhKW4SlQMceTXNUKtKMEGu7vNu4i7Irvg
76N8NNkP4BEX0gWrvRZ0dW5l81ekkpuVPfTFIdVG3gMaTXkJE+VOtCRA5TmRdj9Z6ak7gVLYFy7t
DeMrh0PkRF22EkGGJT1nH0OoYZI86c0/MbeyPpsIv3TXIKBLVTWb4WO8kJW81Lu0zhtfxBmt4YuO
Hs9Ym1v+CiDxRZZFdhPA/qxM5a9dlp6XEYBIbWr4FnmmGANZLeWql0xg8HBPS5lWKxU2nx7JW+pv
NtfRSmPlcq/ra1GARXA50/YkRIro+AazOCWqL6Qs7Umq9xgRowGMS52+HQrEChcpZhnHDrCUQuPX
NLNQK9qhA+WUFy3mMRzrfwW41P084mJdC1VKJ5lkUzETUVMxc2wJ8HmMlTzq8Re1qZpUoiRGA64w
39FprfNuCXIp9cD4ZIFHlsbHeo5kp+0d3z75V75Nk9ZMsSuEmYGZBUc00+otl0zz2czwfLMqUFH/
pRq3A39mx3+TQEMXYqwcWGutKJsn1rF6V0wWB3M9TTZ6bkzL3PqT7d6PSsywGnPD0qZOKL/WUIXy
HtW/d0kagnSoSY5nxtaKLh/r1S3b9pNdbfoC9KNhhwEP01n1HH9DR74Zn6FhNwiu5E5KED41+0QL
fAJNMkT559mKROWqL+FmYckOPcQxZPj6yZvG5s3GJdOJsxtfsqreBSmtTJfXLGN0qCL5UMPu7g20
OpsyWA9SptEkUYYsAMEwjPIr2Alv1DTlfnPG/It+4dY2EjBdqM3W8eRFZLI9nD0fm/r6rN0H6j5A
ksqo2eikLe9eKnpYHkl4DYl6h2+hp1gEXBQziROqRxvJZGIfb2UIr7akecy8tHKW3wXqIamDseii
MLqtMgENaqstnEvGXE4JZP5PTYBvfC+jAUFUZDlEvru7vUrwwTF0ndLFotFViX8/a0+tbAZYQy03
uQk7PNCvlexkTjcBh5XPs4Jlw3KRpUKFgWWFF93D2Gk7NSfL+0btydPBWcXeapzTH/7olJLmXZsD
M/+xjX10C7gabPVaXbmByt2h7qP2I2tOxpAOy5Gi1NDJ0c/6MwdiQbGRkeimY8mTJMuk0WTkqi0J
37xfvgDTF6TBj0Mdt1/HLy/s16FT6sREZ+ak85JSgYU8M46NwdD1M+QFTC0mpkB6RaHnyY2xNy3H
CF5XS/+dNXsPHcJ0NJRH2LCfIeSuL0h7xzk5rgFGu/k1uyqsOYbRHBLjqUYfgYy1+mm2npifIrHy
Cy0gKJI4AYCjmk02AzBGTX4e81lL2S/IMVidl2H+0GW5MgAGmu9goq41/94di/uJQ6OxC5Ip+8OG
uNzDj7WdhraUNOgJug3xC1lXOIaNz+fJtUA7xlHqP8521NbjXy21cLWaWrXvHBpbsIoETrZT9hJ+
ABFLUnzbHcosb/9WnKYKNEkNrVa0CJqN9p/AZFCKR3CpPbTdetgLc8wutJa0IFujd9DI36wGkC/C
avsG56hNXi2U6QgtKuGh+33OB8X363/LZBwWeuknEpuzBRsWmd4hV6uop5AlbMvR10f90JX9JBNP
6bQ+2YIo4c1GLSI/1iD/TuqD2fcf2JkzwQq2iPHxMcesWOKYA1NgHy8hvDlymzCryb9Oddnf/siB
XZxYKAqYiUID09pForaNzWP+JYtBWp9fCyIDrqJrqcPbJx4zflfHd5mNv9abVlBXMKHjPdbwQqJl
Joa3xNpDxDnQOYzOD4h4ua7b17z3XNPEf+9VLohX4LQ+dzSlzKjeSj73E4pEvNhs+3imkJC5TGPP
v24IFYTX69CsYAHeBTekBSN9KKffj7K5NBfp64yFubxIp62daSkvZywqefpzHHYmTBB/F+0Szasq
FD6IC7nnCJxY9c++UuRLT3dMRiHzUjuXg9tpyjree080cPfqv4/2A0BaBHkpcaJq1UYMVWdNxID/
auXMzifvqOAEKfx6qSsz5J7YTdd1ntOPcwZnXuHU+c1ovcuqubmKhg2gbLApjD4LA2RIW624piCt
7X4WCFmoZAjVquIxb7MPTyGmTjZUygaA6kySYKvp3zLAqeg2hpVBikcDd6zYVRIQBrFJzEONa3TW
1TxBKPrpSWH6Ic7lgm0+vcOYgcNiYrQKxdDq+rg8U+a8pESyhB1OOJGiUyJ16ksMnJSYspiDz2SG
CRiLRAor8oXo9TFRqXyYIv/9ginEeCoiXp50ZmMLACLupNuax52Fg+wBnev+3IXasbEhO2AwUebo
dl3Mhcsd4ELfhVkD9yiY8hOhsqmLPvsEnqB/q55JqLNnM5qjykaHW+fxAWVjl8qn1a12+rwtRkP6
5weFooEFMee6TopivuDNovC21K6MObZZPqA+d+fpe+yX85KHhqEZ2WJ6KuDBcSzTdwdyjWxWM0pq
POkCm1FOIItCZEp22VMAnd/6f12cYJdoqcA5OzOOtfK12A6hcsp3VDeurg+azdKmA3DekJQtysX7
n/NXw6wqchdM59D6L7v0EPMbazBs8YRPagkCkgPkaQEN4+WkUZ1uKwWUItOuL9UwsjVngnfVRySf
7h7K5hUUStI91L0l02LMtOtG8oz9hIb3U1faYHxxbOc1aumn7jWYs/NWU/AORE8w3POn4GFn14XM
scuhFYY62U+XEyt67lfO7vMXe07yUfWc6VhdXP72ODxDvqrbmxmTLAplIqjDtvA9npl1ShtrFquh
Vh6PCTWPsVHYwnjkG/Bwv7EHShPcjnw71Ys/Fx1wXhh+iw3uSJVgm+Xc/V62XDR5f0LAx6h507BR
EMzGIb9iejC9YjN32lAYGXEkitgh+bRG99mtuKLbxZknRGkf3d2YdkvKM7KsLVH9YoWZYq8FTQR3
sJRnKKpv0GEIY3nVUEvjIM7G9SNYGW91OFAyX6VO16NshDcPac0KhW5CI+TgBKaLSO/IqulbAGtV
POCTAiQ/3a88foz69il5BbIeeIqYfcI3FvRoXJB7yDI/uji/kjdkrip5wAgbSOGr3wnyHERnCvAQ
OhH/y5bF8zSVpcDWPf2Sy7BFSMAj/lCjuc7Wbv9cAXl8p3/TSgN4Bheimy10jAfex6DHpBTfAqJV
IS1vTLEHQSgCf61diDou8wYJepvw6DyMiZ+8UziMyoA2boJHiD84MjLJOOqHNMGKRVTdl0Cg9j44
HvwxAo3Rz7HTKN/Ya1L2dDnB16O0OLZPDeFgBzG3yeutnN0cyoTuR9AhFS0NNfADYhidxd75/3Lh
2Ylsos4Gdq5AtPTq05epnKk6IUxaTCMPgbPejSZhGOWGN0RNcz7veRKZK0JCPPbppdkW2r3Rzckx
VokvpQQMwEoTXWYFlKgc19zbPUBCu5ZxLhP78j70WZJR70hA1fzufeicL85YtHp0xB5kYW1tpca/
5kyYZh9HTsnJX/scshjKfkUAuByMimlsdSyRSj9bxtVy9Qs/cdN/F0Zlkj6+ETMtYt7s+wUC1ndH
cKYmHUpLx5ATIP2wd+VDVajdtXApOvCEstrLxVw4IE8Qz9ec1AyfTPrLSu2e4I+as1ZObzzYYq8/
AFnA79HV0LcCqD9gbGwZWgyAV9GqLaH3PylzAN/EB+gPOLozTHYCWYJrXSGIQ5Pd819qt4auLAHo
zb5PTrh2l4DM98ZE0eMUUdGMxtyLDOu5qBpIKL/UnPeY6tCuVYuGe5FpU/eRPiJcNUaP+BCEKAJd
M0ZxwN9/4Epuevwwp80Wdr3tNqhkVlTVLIzBZ8czW6+bb8/BBG3Y8UTzExnalTF9hND8UoWi3+pQ
yYrVi7LdULPW0Ifng7QeGCH8jE2SOL0kkaaDRgIjRY5wpvy1DW1nqY5G0YWqeyT5WBqFuG9zfwLo
ltk6pDp12Tk9R3JXWpb6VSNEsv3dgH8oQJlGPEljY0q2V3uELpeb9+cLWRPGo8WHr4SdVv995/0x
LF2HPYolNEXmhbeiETzpfV9mawQ6jj/u3p3FWGEaJZRUfedImTNAv5BN/g5hec2kobjsV0fjBH3m
gkGNM7uhbAmGwg1HLd6fFC5p+nhRYdNQlA2pOqeV43irmEj+7ptGNvcPQsvCvW3Vbp1MJX2jES1y
CUejJMJLFTpfGMnqHLGgdlAS2cLvP+MxXXAOLSJ5sOwWFwzPvDT9GOi98RS3lPVgq+b+3/D12vH3
BHquQWFCWwTmIBTW5dSGT6wW97L33JQoHtltjzu/R34+kAyfYErGRAIan1wRE9enQha2UEHdH6rN
suyX7xWo+IqTc9yAls79pSPgP6Poz32esg/lWw0UNiLfQo6yNCr6lhelfZ+BFGwqZ3de/TDg3MpH
fv0TnUep996W1cfSCNjwAz62+onJYMHIA4qConQILvHhzu18o43R7doxCw09OZ86uiOkchynmnd+
kKJX1m+t263FGaLAsVOopqwu/oWzYpHoQz8YBWtxx/mMV/1jENTnRiSHF/qiUdBUehj6Ip+UYoWb
+icPmxn6ntmK4Qr1vJ5D8aEpu2BsKRK+6pI+R1SFWEgFKYmCdI7hm6LpGbDck1s8uwbI+K2F3zrl
4yWsScxPdtPRROUcFf0FqDCotPfPpeY3qVwpyeihq7C/om7igkg4Ro4kqbqRQxwfJ9p+z7CdAg6b
kCJpxkzHpsTzRyEKdechZ3nj41NQeTcXzkq1QBJscbuLPYxdV7kioVg/GJMuX3PerJxgV7V90HEW
cEO220aeGOufkmqtbdprf0mgP1gJIWfjzsrEHqnISkEzzclrmQgkbGQgaaG4sjLFlJc9rKoxHli9
iZJ/6p01aaG48nFVRUj7DuiJu4l/CeiH0YORHcwcpHzFgIvq49laKb8F1NYEl1dLMBvoOL8JIXRY
Cf25lmKk0UlznsY9fYMAwJxOhGG3Hog1oXWQyZL2Fu4nwkUk4cx3vcd/hOFKD6L2CN7jx0ls1dwJ
Dk9njeLYut2ne89gVXcMwdFivai/hNWu/Cxe3mjX066OBq3+sNg/S1QsbrcepJdJDM1gLYZPG9aW
+icjdnWJtu6/mrReZOxNUOwwOUjN4FMK2L4fpnjnvQcyG5RnZABXp+6Jb5Xg+mb4AIi+ny9YstI5
iLNoPsptexu8ik6Jj5zgM6qMgLKTvULHqczFieYfpnwtmiVzuYQV8zb6vASX/VTtPU3UYCK6zeah
LCeF4xmrSgEHPWF01qWpmrnj+xCfQcKepogCI1a5P3gI9W/Q4ZB81NdrQAGR7F+/8yni3/ewjKmA
VDx1Z5vVtvgCRGlKw46UVQNXLS2a/I5jGeD0SEL9EtxaQCe5ehdF4oD4Wd054vnfY6WjxwPlsCIu
wZoU415/nlIoyrZ7gsTZ7YQbkoKZrA9D/c1OE6UJir+4wWGFAk6k9PohduKKOlKLjgsvnlfXDfAp
Duc7DwQ+Qq6h/9lxtMalOAMMIl01uD7LAWjY+IDT2/Hr3weZkUGZAjPwjM9oHuoWUMqUyKdeL8ZI
Ib7utHfQmsDVI6VJP+zSwD6KusfHI9JtyfjE6WASQlzxnF/ADuB0CqZoQjngou6LAGLQertSdZLE
9qT3hVqxeTtAcF5ofJUNLIFZvivZGzu0PMLa4kvFzWtmKc6MBIL4yd94oqtzWtpy1wG4+wLDe+TU
Ze026X5bluDaLC1YUhclquXhyKG6wrnqKlUILMYNANRd8aPiO+YB7Zh+nDVgmhWYgca2uNzquV7k
O2JcUyrwfoXf27hkCL3E2FKHSzgKAsMJu6T/+jyLjSAePCZrysDsRX9QJ68p7WZjMu07D2wYa/+J
xr+3hVpTs9GpQxmU90CatdbxuRSWM63nOqPdEi8auMSGM7PNryuI2R6QxdrYZdgP/+YZEkisuphe
kVJE93bL4/ghNNmZgFE3/SrxcCfDQe7xXxCPNY49rRUo7EL0lGzD5cRPyKTXz8K8ySewcRPRQ8TH
eeHuaqOO3ITZLAgOfepN7N6eH7k36STykltk6hQFs8CCLV27QAo9swzLeUi63ejc+tpB6kzu1kxx
TdvgnEYaD/6WXC3kMYEvTOoYAq8wEtA4rvwIX1Rk/nZTWfRM5MQMjgNA7FjRFvtzLOb0EY3zM8c0
Qgzeg6cQy73r0XWKvmS5HKuTxuCaTkr3bPAR6KltkyjRhjLJ35dPm/WlFAt8Jgb1W2BjrnqfQXnZ
JgLqZ7iS4LwRZE+dyYrFvR9qdjBQdc04U1ZFSiwENJkmFtNv2dm3eUGR5GS5TTO57TeZcxmawv49
V2VpTzYSfFyrT+qKVQJpZInMsrlp1FnHQ5yREWOA2tR/nWu1KCsZuU02BBhAunGxxuWxAgJMpzE8
fUsRUBibLqac2MCKNTmQJ4k+pa5PojNVmYS7kKa8wf5Q5jFCSGTqnVAKHe6+RD1CaF72tNGNdly8
lxbiOhbIisuLWUy1B9acu41XCl6cgMhtUjYx0JO/w1MORAMnICe4C79/uGBNpQavDsbLtpT1WXLn
WsjmGMfp+E+r+M19L2nlSkpELZQ4A9Yion9r7Oz2Iq9mG+Gt/aLud50Ta3l5ACLvlNbxWXSDPdML
HC3vrWaiOS6Xaxj+RhE/qDycsyQktiIT53umfurliPLygoVBhb2UexWaTuUkuNjtDxcZU87A8MRB
11VdcYM9/tGLc0AlUGwfjqnYj409UENcIH+dm7nRBxPcBMC1P0omPpZvHEEVZWTTsxcLfEnskBW6
Uk7tb5hJ/QpVd9BZzd7/FfaikTafexQh/3Ic4dakcTUdDMsdITyjXU64I8lNI2RrxyCAsLzx9mKX
+76ij5GC9V+Xbwm/exHPJkoegxLHUStqk5F/uYfq/1BrSo3D4zSwOgrjxy2wpbP1660FdJzrmIDT
LsrDp3Uj/S+OMI4dhTk/9cPXk1hVAEH8bfTpBPg/NqiSVwX/qtqVwU5y8HEUe9gkbwXk44/kMhdp
+ZILP3Jdq3wZgyzkYKArjjVniOP2d0Ipo9RCCZg+V6vTtif0fOQqv/fS4ntkvfqL9XkTB68AN0+2
P7oEY9WHqlI5YEUORX2RYQdSAdSqT+vr8OKYbaO5hXboICEcxYDAegwJEmsxqOTMMHEw4aYGLuDd
x2In6JxbTdkFim0IPcOtlvjBjjehqVoSJv0vj8+55Xy38Z4WnYjbD1DYle7BhXB2ITNRXXjdCCNq
+ui48ROXInFaayJEjsvbUSsClpUepiAUNM7NxRDWmVxkO9Ce0LsmBBFQXKwCrBwq0i4w3DucJAS/
81vHlAIoWC1FbQwsh5OruN8idOwGuTnIJnyWrwUCvoxJtsGV3/iFMpcXZ8xmaWri/2pbOfF3Io6a
O20JwEmxDLx5WwQfLCKXjHVtXF6kjOpdfkD7PF/8HOoJrGkZflp/iB1JQaPpHnUnz4Zb6CZgRl7n
/ubZJK+Kf3kfesvUFF1yER6R6QFMW5Hay0w6krX2Pg+l6G1rAvIvQaQoGZev/t1wtMtFXjANuMkc
otD0vTv5NsmSh1WlRGl+rBhVR9FCJ7YgL4DLTgEktjfds9zgSEzV/v6Qyx5WX9iv8MWxCqzzAbuL
+zb2FJlSpo9oV79t+5jh7ZwmdtMYd0nnlFw82OzQvypaoH/C17xQCUGl0XCKG1xvK4ZPv1Nbtw+k
Kg4NYyURnHLatdWOd5sqzpgjxzwr/fgQuzU0kvCCZU4h+hCkYqHGq09Mg5NEilQ8fD80Zpl+Cc9D
shivnd7M/0TrX0yIX50QdXozeIaTo4n9rcD6qe79UPx6+FGPxAI3RdFvHG8AP202xQorTHwkfFJi
rYfj4t1tOm2TA6u/JjqXY8HMp34dx6YaOAMoEZDY0bLLWPQ0iKYuGFgN6Ix4A94GmFc83NRxTWKg
b2frsiZlgCBc5RsO35RLzDVcCxmV0padGDlyV/yf5vFa9YV5adg2n/oVtmrWvOYU3FHBTPGr0UD4
gBP1sRytdu+HsMDiz7RKNoqo22zagEJvufTHpl07uNxKErOykh5R1uujV4tlkQ+xV++Qtjq9ld6g
/FQHNxf3c2l3Yo0A9skR9vNEcb/pjYsuU8j4ZmeDGsFYHXhUiui6W2AEKAogjkzdt7qTpqzkdKru
SxfGZH9EcJA7m9/oBNP81vAVvOhQSDq24acp2cIml9MoDqEaD2geUVO2WjRBNT35+EEiGv/XAZ/U
76GM+K27gxyqL6GXTih6ownyMF1EDIjDYsxRFnAmAhzyBeZUr81TrVOorfNbdDnz4M5IPWAx9PQQ
GtPp4o9ftnLxO0ozZ28FzScvi+obfLyy1lgKCnvJFUycq1R++wxb5j8neUzvq1w6VjLVOqwnrmVK
wyX2nwWC9QNYZonWCHX5UVIPpzSflqwGIbCR2ARQ9n8+104RfNAbKRnf/dK4yl1Tahs+W7Rt8j6U
zADRA14ZQvEyarJcWshgrDsKst2AsQQfqkcfAho3aIpd4kGRnAG2MW59qlNJCw2ri6fVQ/WIKeBU
Xyvvt3w7s+NiWrjDwx/LOK4dnwoqzjO7AjDlR3l71ftUCCMSfsmnunKLYZihp3JYMeiido0HZsC7
Oepf9ERuHy4Y+5yEtYRCM86ht2QsEsZdxc4zRhXoY0QKTErPJNTRANtm/mfUHp/hHO6zfvDj8hYk
U7uQicXZJuNiC8HwRWtf/rwglRGhTq7URp/f5mtIoQIm+oh4+RDESmcw7yE5S9Hskt25dxdZNEvj
kq/qJh6HrNknNzWR4jIKRXwKdWRyeLoZUlTq4K6ny0PlI/12TBCT9FymsdZi0rK3/bQQOv0NSLuA
foec05ZP7e+VU7CHLh0mKtEKHzE1bdYdXGo7gaqc9B3kKXMVukadQBDx9jpcNIi7fP69r+/wtf0p
325HsUEQYTow4Y4d79OGm6Prthwzve7xdJ6ibMhlval5OfSCAmTM/44oI2iGAohrY2B2ktW4z5yl
MEDphgFTRy3YWJ+M6i3PebQirvIuXjYYMWP9gILQRDmaxfmroJGYgGdk16p3UWL1Bw+NlZFMhGWK
MaydjebkPB4mGrZ1Jsd3Lwu1Cd+lmRSEHIR77SXHN2R4jkvAsY7oA86ICHWkOY47FTTHFb9+9RlA
pAUqQzIxb60/Wvf82XDevhMWCtiQmPlJjh4Qm+rhiiiiS1uDZ9SZijgt9UCVSL5c+MXgIHke7LvG
5CY0H6KedRCVw072ewNcQsrTVIbSKFw/qvFrU3u++BHdOhS6T7zpEBF+iXPE+X/X1q+OdoDfAXWj
pBajGIGHBQM6+iuK2CIwybXHAUeO37uHy56jm2C6mqIvgYIH8VHd7K61JNG42WOfWXbNbRLHC+U1
nYlGm9FWOM6tre5frE4AwIOuosAprlkU+X32in/1Fryr6G/Bfnj1iL6alkAu4RmoA2H/vUXbc3Au
CMSZaomEUQYrmOG0+Xd13fWgpdbyC5V1qTLjt0UNINjz8ne2bF4qLQfu8ws6DGMKECWi342aZ7BO
3i+OSZSe7BDxjAiEcqjEz6+LvozxkvW+oBMywqE5R2mhPqVwg64lU19ciSbb2x1cY8tknolwvRd5
DBrph4fgoKDs4LivBKKmRrX43HAsga3M1j2BJqXvENsPZIa5csqaCMGXK+6vAHH4E3NVWjG/fvbb
Y5/aYsE16giPm2aLOPqZ3Tn27ygZjgezVQc7rxwTkQjuY22To1dieYlJ2oCxo1rzRx7zMl7VPunR
YYfc/ggh5KEv/8YBeKjO7u0AtykOQJnAP1kleLhud+8sOlsybVzCyNoR+I1NJxHDeZaHt98O6vvv
fQGpvUuBVJdjvHXXDHTT4ziIOjlRfJA9GkOU7t/qpF5eh6+OPOePXiyoxDBA61rRPTXHG4qg/YzX
0L8L9AJ4160OMre7bAU9s0xEXKb63np6l2k0BCPWUhYla+CcsqvdZbx/IM1f5U4BupblU3mNmRzm
QC9Ht7GIVdcAVXPxwb5zkCI+XaqhoMqT3gUiE3CD1ZVoUIGT9ZZFs422bMrKofsNt9Kbqp+YuFWr
E7u4z4DafBzcaoB5eFKEoN/xfXRarDlBjDrx8NyrYMeu71RtsYk3G3/h0tKWzBISfh03YuPTy1FR
NOlVP/o/9xAszrCLVqB9E7uu0jrywXh1FL5c3qNI2pfBLuTBwYB8xa958vtfZOeAZgmhIw3gMS+F
P4zDw9eRLEmxK/ZQ5ibyfQ2+lP7+/eDFoesgKQi0mRIE/BFyc627aQnrLk8Ho/dQyVepbAUb2i1n
LA8zzdrW9XRozg59p4uu9Vn0Kq4gnQNLxWYXWu/eztK+4ap9rsLRxaLQca3Zw+TpUC72f9y6TCmz
zM/1eHOw69OO5P+BDoVft2MpH3Ps7mpTNmwOvzyhd7Hi5R8JjqTx+7FcBYhN6Nmwa0GjpM/L5Y3P
uDjZEGMTBqqATovEnlySf//KrBv1FEad1Cf7HF4KXpaD3XJ7aV2BhNnDah1ihcN35QGrf3dYm71s
fCfDDlbU5e+0kWcS9srxZpYF0hrm+chy2o0Fw/7YWhrCrdagS5SYVNDPzjBxe8aUCAxBy4kgvZsD
zgkokQVexmESi+XzUADflGDwoFy9mfd/Ls4UGKCig47wQHA5Um09YwNQ97eT8+bRV0bWQdKD+FX6
er4hI5s/Fhf6DqYPtDhVsrsFiKzOeLqA70iZXUptiZT6hunMVgG22SD+5WS0CcP+4hRFq8s757Jd
av20/z4Lor9ns4qYU6X12NH5p+llFUoAT0bbadKMKxeoMLgS77N7/vDKNFdGhhrGt0/abpmhxDCy
r7iuh9DZuR0Ml6A3kvvJJ5TPq8IpRV4nkaps0ZvvyMCxC3VDW0UnYPymhqpvUGBIu8noUTFW+Jfc
AU2KDunxkMwpt4tr1GMsTS8Bl2eqk3bfgp2b8IYhQ2FfZYv5AmYdvT4L1e2fjzXgYd+j/T3nNibm
6hVOWOerPErj4M6RKjMdaoLj3qjDQXB0ZqgLHS6nyj736x037bkIsF5w53y9cbOLpZgYQioPcuaG
pw0qLAHJc8wLsQxIUHumjUE4cK5TqXH01BUyrJWSjqkMxHCsBivtp6e3LTnsbNcEBiwTtmNE2vkA
jTPiF+X0+R7fNp15FYf88pV9stJBJ9nbFGf8p6A6Webt1mrbNHVEg9UweQtp8TUFCDBri6QdS65b
p+N1XbGg20lShV0hG1lmOX8a4IFRKfIid8fXd31tasuqnBGh8uUKhQfAn/vpnvRGERSJdpPk2VCI
Pl91bGvOH4sJrf93Wj80d0pn3CNKPg/NYHZ+CbY3eJRy4rFD+D9N9TIcqSXpz4P7g5s9HVllhbSC
mYe7bmcN6YADZWmJgWe/dBZjkF39WJ3mJOX133A3/Vgasi9ks5Om9R+AwO6x2eA4VYpSMcZHDg9n
5I6WYKgA1E19iW8lzVJ/n2gDVBjHje1b7aW8nFVMH7jO+IA6Jc7L70NwjLrSkythZEIzMacQlWkL
DtxmdznbHtWkwHXJrlJ79Urooupw0ocC5sT/r9MtmRWThY6Ni9ibSu0s+tlFYtma45Ar2FNrSsQ/
CfpVcWGNDA1aVEaaHODjCgCSz75p8/5DyxRXljhnTc88YcJ1VmGSmXgmNT1lf86/nAmLnhW70hmi
qoryPSebUxbDyR65zihhzh75bk2YpSm35Kxcspw64F3z1X67Cre7FEhA5200JKYSbpVhZTCENwGn
HU15Fg7ohobDGQQgBbMPpq1qmpUDJ/4aWEOAQYm5eKEeUWFfByABOw3HhCuKnuz/aIY43tluLnii
DQqtRlWdrvqmUJal874cc5vv03yVraDIJPuq+SAw8yyvTAZNlXedr9j9LaIgge7vQbBmX1knmE1D
25w2ZvvtTwZqUoH1hf6CEOH7q8LAWvPDfSY8THm2Vyn/EYDcRMwYjzsxFpuckoMA8VPveHDY4tyQ
dFLocYa1H9dUbgAfKB9Ho7hufSIO1dU7igxpgf3FQ61Vw3v9MnKuYU6ik1o/60mNbmtVlWs1ix2f
rHhWgO4aqfqg31L+Tn3aOKJmnRbM5QNmOFmQAXl11vGXueR1l/JJ4IQPfo4IaimzpPRvQZRZWYaX
QLNQyJFgkDU2bf4dlsGB7tRhjkVZdTF90JpDrm+IZ0/F46F/Vg0pTQ+n7tdfSFMYwsixtBLcAQ2R
HBRULghzN7sruP11KwGOiog3m2mKWJe1PGxt+5jjGP24tYiVTSMaPOik2681W3vkj9sfPpNyhB6d
xvDSXcb9PyhO/cFP9822dwQ/7TDQDltRz+WwoHVwgoboIlWCzIDCHATfCcAe45Ja+huD2aWwF2NC
VpQ+X5JKFwaWDwexaHIPfkKJsXYVXPCo+2f01Q+K78yzHjVO9vsC4HnnMQMYWQgRk+aa+d3X/T0r
SvQoq3xXh9WQa+BKfDpZomIasESX+sAU2W3+86ux8BerOC1lfESq6MExh0fwZokbfYOJEOZHjm6w
/rrpld4/xQWGOOA+xhx93BPz8fEFsmcyO9EHP6bt7p2r+fitefclUlSCfgY13ZITnfVGjEA//J8q
La7DREkAQgmul2v7WJrAQdyP8LT9Du3pIHBNMlj/GIGtHQ5KV2cQo5qC06K5NULUeRBM1V1gKY+X
mDcoZHwspDdBgR+W/HAPDvf1sVPyC/IhzB32WXBam21fnCR82u7dNccyGJSvC9OU9n80lcRH864w
IPLDqZrEQ8+JHj9NNnc/xijHmSn5P7AN1jQurMwkaIzREtvLlXVr6ZEYp62MUsc/w0Ou0xz5cqLd
4DswMAZxmUA9kZ5D32ygGcSeILibC5/M6Kzb4Y3opxpzaCCRmtAYjpZQVQozjk3jYuN6ZhBr0NgY
iM1m84H0beBBJG6fSYQCSkILJu4JNEGmidyjqY662u3DbHrCWBm2S0DPNZsfPltYOQByvtZ0roGJ
g+xGpTzoiaYUmOLojPXNgCVIHrtXvqPosFpO2IGl6IQvxRD2Ys0kIzbTCOYL7oU5moAHqwuAR5CB
KWQsoX/cZaTKbwRVB2PvMJT4bT7t/OcrIhCP59B0zM+Y8oZb55NTeCim8kxs826NBxtzmirLhtEM
KPE6HobmTIhDn73mJEA15fUnwj2h0rg0vPtMEnGvXsHhwIRs1EhCJ4/D0hleNr6nmhRrY036PGpq
dUZgKABZrR1+Gz+qdgiSA/vSle/Qmc3BgMF3mb2lJhywzq0q+t64CExOTjsKg1Fvn3XrDlIFwfrI
1bsNS+W22wgxobE5gUV2Em3VW2zqepsoxtZKW6/5cKSMIvh8C4hUO3eZUi0vL26a0DQxEXpsw1rP
3of/5W9Hy6HUX80l273za8/kg3l2V3WgXJ2RSUJpQio5/stVL85VYwxZduw7/bloqIIvu6OkSz+X
wetBP/sg4Prr5ojOyMJnmIm4pwtDNDWb57oMKW4jqylu+0NwpQzWtirk97zyXZIJWxwcET2tkMK5
jk4/mbt+cxxPgxF2i+E//DPO2+zGtemGhdgQdYV9y5IF6UtTjAp45bDM3vspAmP3VoOQn6iJn62Y
5UxPBCfFgQJpWXEw4XmXSCfhfGu6Ru/IMC9IszWnrWyinC40bWg+ng2wSCz2WUiKoKOHDW/IONSU
3ek6MftG39CML1EuAfDggTdTNSIUjUL0aYYsAS9zdY9ZJBxXpbgMDerQRDjyhUt3YosftIX7Tn2H
zCVlKTDS55PgtbgCjJCXboW+9kuk9fmRzeLjVsXJsK1YNzbDXY+FcILjHkG0LRMnFyVvaXkckJnP
XWdQo0BdlTBKfD9x/88ATMcdYgMORMfjS6OLfQHypSTFpsdwINSZerGwTXO7nlOAatdxWR0+uDlY
rfC+lgtYcWBnfTrkqAMB34YhbHHDuu0m6MpCwcM2VRbZaGfAwkyVTG65MYL27ruSIkkmvXMvfHhU
XzPw2CoAVpKgiEXMNyWEPeyfNZrK/rAUEDvc+eeZgsEGl4oGj/uc3k9aKZUM9OKY+N3C1PeO3j+S
3CCXALeNFs8cLqs3LAoTZFRORGwDIgZ8CODOEeuo6EXV5AeJ2jFaFQWQQQr5zCeAVSDeGsSmtEcn
bFbvEwi0Orh31IGPrPE+4nQ3/FidvpwblXPPrRvxbzVj3WTix8XXlQyBkaqXiBosn3kJ4OSS1lKH
3v6V1h2F1V7m6yoCLsQ1fIcI9ebPfwr5+ppI9jb5dU1+IXEpNTO5VKI+yZjm5ggaYhXuel0eRduY
gYaeti/HNtZJbA0UzxUu7daLOZyYrOL/8PG8knv4gSLrWMjmW8eJ0Hkza15tc4hdu0W7K/Oy1z+i
D0vUmwDa2D5NrSru2KvnxaTpaAFj0iwupAMmVcH98aqDWGWHu48Tp8K1wCr3167GDEcP3Ep64IFp
7EioSXdLhGDcLy2r2IV/0ffVUVSTbh4dSF+RNpgdwm9kE52/5SrQH8cf1Q0R8MN9/x4OBIR/nOTA
RQ2sdXghEnJrYK6Wy3x1KQXUhjRnHPnR01uFSTG0YUrjucP8rFQRK+ne842W+gqh+HBN3XJN3B6k
QkBa/2rYutigKek691a1Fl50KxgiS5SS+Au8r+t4vFEo+MVmDdRJIBicxeQ8nI1kuW7pbjZTpLtx
zVaMrAQyab5rnBIa397Ju5TvTZY2CRFzBwU9IH6OrT3bTprq+jtE25s5stpaijZgCtfAu5SNkD3f
M6Fl3va0NkzoXGB+QMzQjb/jp/OkjspnmKLXkCxeYElavS9wVyyWChwpNuofAAvq1yi7dSknHdpj
JC8VifyUh1UCL+YeKbk4/uMHDono0vjNELYg/otzMSGsGdpPj9KrifWNXJryniAMinhCTBSd+cuV
j1NO1W4twmckv225GJg9pYNuWCYMW/FaNC/huev1qYdt8YnUZJZwCyTf+de5rtTylYj9/IGeDYxK
iKGftioo5LSHCigxrZW4BkLAIFvOPuW7UXJdxhpPZ4Rkbnarqp5MiK/h3hw9snrcyF8AxRXu68xp
wgOE8B8Wc+zIJdWrM2bWGiMkL+W3E8yntL8VEHBvQw+VcWB+v7TU1QdRNtOGLsUl44CjSvtbeC9q
psiKckWM4hrPmFoubMfuX8etY7hOI4FOsDlr13g7uFpld1Xs3coLKILDOJKaTBFmRMPpm+8KbBkl
EhV0HcwIi3A0DgP84/4eO/RGP8GEhYoOwqD0PszBnRVDVYXafm/i2Bpl/QcEuRhlTUgyjWMCXeqh
qVLH8IRHs0dqk+/6fJ63RMe/tUn3joaePy7T1PG2uZoL8IeZjvkAG7rjsGKDxgjV5QylZLP0lW35
s/2luy8KdzCE/YI+Lq4uaFosdWxGCZ1Pxa4LNCS+CD0qRbstdWEtT0fGc+BepUOID1ypzd6Dv2bs
/Bbn2IM9joTiEMKTFQsuSKb9URDn2UnFaxHJZANnPyltg2KTD0YIWHRh01OOvC475oPrfuOdrBtM
OTnNG4VWblVfirMPhFZ++c72Ij+r3JvpEwSidnWo+ksSQUhLucFmhKb0t9LgOmBFBjHQwstMgWPT
yH3W/zzFk4cHfej4a3QynR+8DpdMLVr9g2xZIby0FoGxMd1onTGVAjUIlvFMhC1i5iC8rjTePcim
E7FN1RJrZoS+G6Ff+B55jXIXv/9c88GkEvChLJy0EntBFpgr59iWUAULKozpukmMRYZD1dtyl35H
DzE5TVL6tMDkLbY2nxyO5lg+Ie10NxH5DUqJOpb3vSqdD+ChWzdyZ4fbk766ErW6GjT3z6cEu+Ks
jyc7x3TEZ3eHcFi4GlXbH/wRPMOw9//OzKFnMBBlq2FqKFsqFgv0blPWJl6adEEP6uBpPJV8+kwj
74QN9OBz1WDnhUPHZSMfKtDbcujxvW0p8H97zdx9XcjqRbB/2E/HLgBkn+JyRkfBFZwPC2EyhLB6
PZ4L9SXCOGx7cGpnDYTjmUlUSEbzuNqiMjGIdBBioejcumKUM/sNY3tANpqZFoGWrTNqW8UGGwp6
Tghed02NwluwpfEM1GWFA6OZsz9KRjT0oxPfKoPOn7E2KmjhQ/3qCCy/CWvKdTcqGisg6sTiSOhi
zTVh8Fv18TgXyUTiA0TRsIJFWQ8ele9R5XAwcjVox9f8AdFmznx4EfkdFzDm50JH/OsHM9Cu6iia
P2SVDnSGLHnxQ9GTlRBzmc+9hwVJh1qNcSZmfFxAKfdWdPybljyIw3oxDdk6LShdSVqdErWHT0iJ
hCMtTIDxI+Z9wdshvyY7TcZmRMCfUEwIgnoDejyh9TKi5NX/ok+ZhS+fiM9wwa3zik9Ce7fDpXiW
lB84x8bfGYzYZ6gYYh4Bab8zlv6ZR5UYnEGf6rJ6tz5VBPppB66dZOKOb5Kgn7CxtlGb1u9IvpFq
Ic+5rQS5yMpk2M0FD3ENj3dduT6HQE6omR1AnLvtKI6zoOZ+6dZE3bh1qkm+R89DzJFnr3ZBsRYH
ERO73qYoC9+dAZcrKWKPCln3QKdes6N/qKbwPliaLIwxnDuCNYBo3IplwBoJKo2AF3ona40HnPqu
o7ILG6vkKwH065cpWLYBzthFecbFy4QwbL1UPftRg+7sRpZNZ9SVTcxlDB5kw3IZ8Vvn3ZaUOfJ2
BTOrP3/ldHWegRxLWnbpHg39JZl6NVGCpG3W5LUDyiAvRjxZg2FQi+hsnbu7jJT+Vb1XbDrPj6Gv
EgsaacUmTWK1v2kysTwviGfB9RV15gBopljvSZuZDd3DeBSAjWccXV2JvHaoi7ml9aBaEsbfxIoo
rX/K8gDWmm8jamSb4vTgDHyqQMRW1Y2uZzLuVqvjoPD0QDT9Cc4j+B98S7o/E4dXtfyd9j3c1puk
pFf5fej4GerymGTzNRymXf+DrdqcNUy2vEIUQDPoRjwwU7ApetA3g5XbbDPZvgFALRuMrWh7jhNz
x8amCuTjdeVM1ErHLTCeaqYalcR1thOByGBKw9YbIvKqRI4u8UA9otO6xWtyFfs5CtgYQYz3NiKI
SX8ooPN7XnWpwZ3d/puqpwBmJeWue4IzXhp8V+vrawiE7WpucSnyJzVKFut0BzZAuVH+sV7WZKvn
RypOx7Sc2onLw4T7kPtm6AprBwAnrcCCictz4xfQwksSfztKYiDEvCvHTp2crv2NWVKetcA/c5xo
7nz9pIlRQJz89w6WtTkGRsZzUGJ+2M/YGVHPIgvWc2au+msWepcxUia/dDySGMked4rR1KMLbf+o
sDOtsvbUn4LWEDsR1yqMs3ppArx3ptW6i3Htx0lhm1NJOrD0WZu6KjPH9DhZ5aoo/Rh1nN1RUDCK
I4IY/sddgUt5dBplTR/+C8Z6EJeKhGRSOUqo+l8eKWf+CPE95zNW2lSj1TrnuBRKAJsFYDgdAD+E
x9V+9XETP2mmDt7UftgEGW+psEJFWZyLHlNVhQYpUcuTJWvqTaW/FQzHJADEf27Cj0hSG6LurH4E
aUvrAsdfRs/wBhfedmGe2qw5Ekz+MWQG8EIT8J7ANdUmRabKdLcUqFvBY2wuzJ1jOVe4TLw716fS
IALUSseyAwRUXjLNm/ZX3dvfttDwNKPrb9f4hnMo0JpIb77pGmOxrPN5/kyJDa7BlPWCEIC2MDvv
zT+Ts+t/OPi1YKB4px5dFAsPZzYHfx+3PSCmnlnqp1bCECz16aBnfFG2uAxhing/THfbOKLNem7u
0lW6/4jiq4pFcq9FhBVNDhoYPMq+nMindMzAFf9kLyU6EvpbOJqe8AhWGwcZ77oBaJCJTqdqedhT
sG0d4jlc0wlBXWGHErV5zucmOfdImL+qKoSIELKC/JA1kHmBrtTXcUsoOR3ux6bGDW7zeGU+MzHv
3MmPKfEHRh58MJUxNJDZdzgmeWxHBKvYkHxGx4GTaVLYDBbNPa6TZggaL+gunxtT+D83eGNQ0D5d
LmRBPcQZddmCPVASjKgZpEQhqokDM3Z4C8mc1dz4bXp4aLF4z/26AM+8SrhjHPfo87ot5Tj5javY
INHI2Of1QYqvtoHg2crAgCiHFIvsqoACEGwJpYBJWpaCMclb4DkElzebDnrcv0qG0LzgfhsaolM9
6YXjhLE+7U5owbueHKaneqhze1zArUA5ia3OQZIS2sIvO3GRc0b/tFVJ6mFm97XTHDQqFvWtAl99
JRAnqwKeTVSzFlkZ7E14bV8KBODpdYz7QgXheXozZIR6FTNaOy9XFmLe1HkMurcVK5W1MfdGCcgu
Se5UeNtsfkeRf3le3p1AXoI03DW47abiZU1rHMxDL/BzKGSr0YRF0Pkwf5cT+dYAdfHwA++bKXRC
A6RlSP8vmoDJCDd09kLsElAvdrHAz3Vgo83qGt+Vg8ALrWvzkXAsjfnHZvxxtKjrqQ/AGvmxbanJ
6iQpJ0yX5CIavWeTt8riIpi+4wZxuUnTWpxI3pAF3cdsBzxuyIctnEsmE97GcJn2H7YuClR9B1BS
7yQ83t/rKDQj9oBRyNPLcvuB24vqcLzClHSZUnNaFemLSsK3x1HkHShf11f2OzWefoqcnkqGkrY1
LbwiPGlHfXaTIVW8/aa6Cg+8R2A/6qeDB1YlScF4HmPQA+cc1Pt3Luanq6buYoU07rBkRR6tLNv6
rsxX8jWYKfTbV6jnLPJ6nJiI52a7WMOa8pFm+mYkyjVq+/JQjZE/9702Rw2hMd61j7zbA1z8NPR2
vnGo2QelONHZESpW8Xdm7P1X5/xhErhwm03OlQladc5ZK/Dm+oeKI1ghwg0ixngjZzAvjVQjU/nL
fSyGAOFYErfl7CjXBhocCHHmE976SpK2WCB6Bt4KoMDRrW7WyKFRCHPzIRMeHoYquGQnEehYBUQU
W385qev7VTLPxwHiSU8gX1VO3jafwtX4ZD8KLjBJ3iMGtglyKeZSffNpQDtYc3G3Nrp46wRSGamL
ZqFA0CDv08v7BPNHxwVvIS+Eovq/A8nmlXs0dCXjJKX2qlQaVpf65VxxUfZjANpLjnhOn7cEH/2t
3ABFyTV+4peVsLNvQOuAldrAUlsvS7n+YIQjiZ5IPf7ALfTbQ7lK3H+KTBdEqaYJAuWw8L/sRn4m
5lQU7iAvg9WbrVipsLRqpCl3LIj4fgVm3Hii1B/it8BqC42A+LkyqSiA6JVT7m0/j3KiaYTkLIwo
qwLIq91XkjBezIpJ41GveTCLM9Fj/kdufsCABtIOWIHZE/3+4rfsX8EuVmHMuyiHO15VyQDfh17e
LLVZCbF1zHrBd5UwZbmSgakaQMXIoAs+1YXuSO/kN/H3s6EGwEufqxwXNVyWLLmiRfsZxD38pkXQ
hlhzpUY9nXbIb4DehR5bLwcM0bD+zNUMzt1HEhbl7XYfZr5KCvELZ4rYpTT5hBIUzP3aH+9cgi4t
9l9HV2ahsycetT9mT10brB/OMYTD66KL8Lou0Z12g+Icp35v+Acnk1ljFsRQfeypzryBhFQFATTz
34u9R5YEDpyCQLyqe0qrFWAAJyD4EMLgjNo7Q1doNkXqgQO4Uz4uIfp4yFA1wIOoggQC+JsyssUA
SobKhlz9DweYinADdDjaAjwSBvbVteKNhnoOmLxR18HETmdYVT8bSMrAzxs14/Gp7wDuAGzCZNTt
hJSU7HAdLB60eJYX3NFxFxpNPVFlL6SW/b7EA2V6eZnPWv5NhYqJ2Xs/gEHlW04AqLujoENeb9js
71Se73bt7PZ9JI9NsUcBi2so/KePa4DbEgomIP93L+vAw8Sa/6emw9dYFeHIunG4+KxxNrR0oDTo
Godr0va8K6s1coO0hVuoHCr7nIxsan1Ad8mrQ9rnVEi8vcoCPr1oHwAEMaNNqgEXShku06rxUFlB
CF4BjXTBu8nE+U4F9s1m+Ye/xNsZe592k1AZfSwHxgYIsD6W0YYvZK+1tXUf7D0HlQjANBJ/VKVl
Nw4Am4X/zlkBjVsiGZdOg0cE1QlwncYEAjj7np2puQdL+T/YCO9ebngifJ0rFMsD+cfVHJR1wCEK
/nBuAX7sKmMJ7F+A25Z73o1rMwz4kFgUpctKDvI9MOuw9OR7fZLE+LiVFcPWbtevDXaXe8ET7zcj
kq0sUf63uBtUfH61TRTE5j4J3Ij+IP4luebdkA3Iya+nNb5rDcz2OzMY6JO8x0zPw5yqHSBvFwny
cQmRATksqFgtOFDCg7hvsKmcukz/UrO7HYWEfWwf2pOB1WQ50lNQZGhNxxinYImuVgkScOYCnLp6
o90Xqtb+EwpzJI0qNL8M/tXx5WlE+7dlte6INktILyXC/2g6v2O4PjQWKDGYgXP5zDel0Ogj8Nww
SLHkt1qRoBvEeicc7cgJ+CMAqquBHpcpNJvlrJtxLK8rUqX+JEDYftg2SHaGC3EachCPiMzaNWha
9u40pvoXBAbdb/yFW/1tcJSaPlGJ+mh1suNM3FQaeCQG5UuavJRlTUFmxXsHD4oOWiFTxED34jxm
OfT9i52Ftl8zCurCq1I36MIZxuOkRQ8eTFnOW1SuvBc7BU2U851BR3NQegZOdcgPHWL/xZ6Jw4TT
AXqNRhHqykfAkfwCB57IL8gOXdISQsGm4yXOy/3arAQIr3UvDqs4HzxjrmJqv1QOg28s+og9mRxO
6k4aoKNVBu3kNTQU/hSxf3dTqVyXrdSHmXwnxpe3C6Q+j4YDx3rXJYk6mse+fdsgCJ8yjDov2ieX
7z6RS6GNwgHh5hxsNwA0vs5jPVURzbAx0EGpybvFeivD1dw0n8sWZXjZaprxTj894FDN3NWmGHwr
ISTvQh05Y31ov5hg9uvAeRiCyfLAa7Tw7C2MkbnnQzrXD64ODtWEmkgYB9NbqdzBpTF8m4mnLuQO
nkwM9f2IqAC9zzSwfUIBz1AmPjYXi5Dsyw1lyGF0/Egy7EQXdX0H9EsB9t/KiO/li4SLxlLHbkdC
0TP22Els/9CmEibSPMN8isBQxJ2LAV9nC8tHeMAaHi3AZLhDAPx8gT7laQmQIsLSdtSaxFOYm7Oa
TDFRRBlGC+9dZb+mECt4J+UN604ldyzdBq9g2nR7WFjOWnaUB49A5l6gKDBuWgEihgzaW3S+DRoc
DuV92KAFx5HAr9Tyl0igLZWRnR24qpR7HT1uAiAUJ6e0rp+ZRnew38yZTAYowo5tO/hh1ggLE7LY
tN4zy/9khPTssX0gjXg3P9lcZlj18b3weTl+6v3WKsevXFnK0b2NVSkZFt1DxeXAVmxAnCCmJ307
IbzzXJVXqIOgUuXdG9FBZcUhWbJWt03XkyPWQC/I98uq8hYAqKNRDhiQqt7yJXl4vT2xQ9jafQNI
lH+LI2ZLoGo8fgSKoE3xeFuKF1ucwOiAVxBWD79BsXOKmtz/Z/B75vomJFdaLZfXTllct0tRr+6M
REtTH8mPl5IiRY2Cu3pOh/tv/2FujKpd2DDI5Zz4plil0Vjc5eydOob8aaEl+FNQXIk+Dmj+kL3i
BZoebC0oF+VVRXraPwAgTgvdAWDcJV4OERMWORVTIoh7Zj/Ixs4BKFWDtK/iwwNyOOkqMCzTkLuK
zLy2H4n3D3zD5ZQy3b970uZbY6rm7l/EopCCHYFcJWaAKS+SfdeWHS1j861dEDZdiRw8wnuf8uNc
GfQZ3CyiQyZ3cIQuoEdrjVl0c4dHLQ4M8WZvJt8x/Az41mvtGpzt1DZFrT//U72D52SMyqsg8GFj
87jw+9bVN86gZi+6Gchp82RZ6HvQr4a2sA1mMaJ7PrI9qjrQbZfq+O+hr1i/59OFkVQQpq9JWCwz
MF2G09b8gHhkSjJD9291v0Km5D/Up6PxKoZRcf5W6Ca/MYRaquTXZoymxSiWuluwtMryDlVJKTrM
et8Mi1J5bkxC19gBWzU5ZKBtbcw5Esa4eZUCVrkxM5HO3dMCbMrAv56K549eQHR/sLeHd8GTdoWJ
+5N7oM8sC0mg8Z1zBq0tElByS7aUH0y/bHcAekqQ4VJNXGXsi8pY4IdWulCZv7x1ytAfJmCbSre/
X92MfxpBJGKjHT2DM72ysNAiMOFO55JAlTdyLOkfth4RfEtGHsOAvP7oZG5+NDGmH/ciBzKPJAZd
EjwNM29D4444dTUVpwS3dvGxnulOrmecSebvjiR0PgQQx62Ni3TyRtkjiOB3uoMiYhvi4UgyvCGo
SB0zNIPCg1Zh/OMNKs4t0SkDj128fqSjUZW4aN08avchxPaYJ5VkosLcoWoqW5H25iBjrgJpVJzW
6o2Qqecoxosx5wNCQcMq0AhXU/oCQfEKSSgOI1fpQBuTiHpi4WMqfXEkNh9Xb4O77TVf6kSXC13H
Ogp5dFcO++ug089VybRddo9tM5ASP44mbmNIz/Y8bffWt549S9mPMNcfBrMwpNX0sAzQ1/GG/ZlR
l+OIjjnTFHsT4yLOt9hvZEq0vmJuLpssXSOzaiG8lkgY7kWjztKyqoR+vMJ3LQ61sYiVyEgl/8UZ
4rCwsb7dlXISJr+6kLkBp3CbvcYq5VtwTMZ6Vjb8FGZ33V51aSZw2ZGdKPEXfiQwCyz4b2Ls/qgu
+lJm+hDMSZ+ZfyrC2OulsnbYLRK1cCXroiSF9QEsaqhlHe/9BvMb827QJ4GaWwxjDfr1oXQAB71w
abgGxS2KkamGqwHw2RXnk0AdXNhirnpp423OGLOzS8Frb8gG+kQrt3vy++vy940jA7rUQH+IfUkL
dTe72TYonAIgc1y2QYgVOPX8eWdgcn1r/FFai6voJfxIH2hNmvHF9qLq5cZ5gfLwfQvooUd+WKep
VOF4HALA6J3IUKQ9+VaCBojOVmGqszOQx75AvvM7iJ4bEZwcK6QwvuqtLzT0eKf5DwX+WgSe2PNC
C1SiRuyqqHqduLN66qeDeB9IebFXuDrzINAV4G5TKh/5dkFCa2ZhHym69SpTtlYHxMqAlbZ839rA
+h9UvvXF78xQ5l0cBxbhj0cCxiyL/hSQjL/5fvOLWtrhhq2doNVg2Hag6Z9Omhg1Jj4fyKuwd+l1
ialYvZ8D36tfhqs/H4xTDxmaEDtzpaViiJ5FIMor8nsn76ozkFOwTU13v33C3z8AANgOT4KY3btq
e2XOGJruuW7vGRnXeNbfrmZe4zI1kYKBu6L2ktXVPU7GzGF+vPDq6/SqAH1g3H9Q2loRBxFljDYt
48oHXiSTb1BChohs+xkd+MXNzc87KIQMJ26ZdDdLXyWNIaLgZ346Fe5JLQSv0eMAe0FNLR3EsdDy
U8mSm17AIlKFxebrUAO2G2WmaZaajpPq8Q7ETsWgSFO7rBa9MK5ZsXcgsU1mOEa5KyQXpSK82AIm
PIFYx0L4YALkzFRjnSVNNc3uV5c3K2R7r/qH7mZQzSpuOK8UvQDg2YQA273iFw0VTEjh24d34QIW
h2NAcRXwAgBWPOjJ3Hw4KpTvBzsriWOmfhKAjUrW16N/mvEyChqBrV5f3q2e9uUXey0560TvewrN
xoKFPSjBBClNJL9saGroE52ZhDYW/IIzXYYdI2/LZqjpv2JieQB5Wh6hbBtotrxQNt55v3rQVA3d
g+JLuFYULOXEW/SQqqQfEg+lZgzy3iwAraIwwUeofNAK67kKYuReuKTfrsC9Rfr8OYxFLom/khD9
ZvmdF8TWX46HETsZDF2MtYr4UXDYb4tK4RinvI9xQz65+ZQ3iCrkL3fYS6C31wUHQlAIthEk77Bf
XPhQt7fsWbTLTGr++s3zg6Mx7iQPnKsjgULjlWltbbJUQaL26JU1uT67YtFIO0IOPq1EgUESoaDy
KCndqFMvLHdPVObWgYV+Z8VqWgZuDQTLgm7LKVQgoslA6qYMzP6cEw1nQL+cjws51YWchEpmWBtY
d7oc7gknFD4va7kpkgdGv2HKpkff7PK6HwkBG4+S0WAbTTe+DLO6WjNDr0xoGI8PbskXWaeZKZ/E
/tCjG6MPUoGFOah0Cnvsx+d1Xd7bJNWNQKljpxZYpJDzzBXVGUJD+i6if5cSyolEuRIpdpO0jUNj
VgvcEO4JnlWjXd9Tsyw5nA1vSKPFDHtKGr811wLOO+YSWDWhNYvT1JHV/YLJH7oCvKN3FOYmjF+d
1WJBBqDyWRo0UchPWdBAN6ScgBXrLucNPmqo+PJVFQ/dp+jFQEz7kxhM9tZDY4TG/IY7qbnodeZG
gjjkcHRriAdp2XCRIESp/KqhK91zx+xsgYCPKtrdWsUc00aiwAfwwZW4X+YkH4JzneIm01fkQAe4
nEGa/jjRyOy/523sapMdkC32tAQviMaoayiRmq2FmOyH3wAdCHeOUFtJRF1AYlBNzvy60an9uMgC
uOJtX06TJ5SIsv4X2BcJzRidXLumy8zv57GhRpW5kKsywopIgNwJiVF1zc/QsizmTLBvanxlZaAK
h0MlkZ6sJcQvg64MPcBPzyC5Cidcp4xJZIA0NlFC468Viag68FRlTZGHFM0nch2PDQNfJR2tiDbi
g4rdBx9ZGKUUpUGKyZCgIb5Hx5sxBW/0HHyYvp8BoS8k7wRWhK7G7MrBOtZANaRT+GMVTmwF9IkR
naP6qWL95bzQmSAkhWg6q56Kq6nRWqc8R8Jue0KtUREZsXdU6xV0fCHcMgzSwm08033ewp0dM/yd
whEqVnqMd8noUix611t+oWickXEYE6kU+8SNveP/o+K2z2Uj5k8ck0OSmz3RIG6cJZ2b1iOXdHCe
FZhMtkO4czOaEIqtu6Xwg3oL5KbUqhia4yx/MwIuN2y53ui1QbtXRKlIJ7ZKUXlLIQCjsspiXfpt
KBFaL0YaN8rnM8xiRoPq5caH51BaS+sktnhCQnzEDys533DXnfHegkx31hodD/flIxoAShw6x3nS
IP8Af9wfuGhs4BGqhAFIZpHPWUEuh3cpQUFDdJu4B90/L456sLQv4MPfgy1S0R22H65jDRNfYjx0
pyztRXzo3fI4qtCxYFmGaJBv/Y54q9Dou0oHrSRN/dmQEKuyoTQZ0tBLzkGyHyBfx38SM9+t65oZ
Ax76ooFQ7eT+aotFgmCKdIkmP4Dah8TTlaZT4XxVSokSsx7Zh5gSCjhm+cmC2Way1LuZfuKTmG2q
KrZlv+AeUHBenx5P30QJwmzIaFGkyxl13dNtNblN2dSR5c7KsezGyMQDm2Peuj3hF9wzxyVDjrtq
BVm8c7TkIIlTh3ZvYexhtM1nr2vONjtvQNrqUVGG7wR9r3O3vcCiVC1MRdLv1v8EPGz3Nr0dx/DK
lIvf0yBVLACAWMnSSSMw7KPExIlI/vYjX4rvgoV82RZXuduTqpKGHrnQf5YHsJjoo0y6e3nRGrFo
ykD3Bodu/jTQHvROdoSlDadT1aBu5c7QmQduHeU3OLPmyTRCpdstLWxVODDpWpbIwOICckRwDP0G
fAPZBIO5DBs4TNsuTKxzpWDoEHXsF82mcYN18M9n/4KNkTKopyi9vOfHWCvbE1htDgYx1N6QL84o
oQXhHidYVrQW6uANE2EGI33iwNpIh/zr3YhJrPvl5pFBn+lQdlK/SRtNQSyP7d/cJ1SRjDzizSOE
UHC+CzVQvIAcrFSoZXVKq+wSPAK46TI8KKW6thk/3wD7/BvlYjMxvgXs7Oqrkh/Z8Yo4fao0PouR
obDUdhk9W/xzs8erd7exIkCAeYyqju4ZSmqI8ZhwWHX6oGDjeYqJANd9CtaQaQgsUHLVWMchwV+p
9cXDI88FatdKRek0kO94k5dJmYdyyzG19bRn09KNkMs9Y28UljNyC6gOaI+9uHnmJB8NblGr3Xv1
qdlZGjzHGy43zWovL6dWy4AJ7jNEvmomb68C6uuHLdo0Xd9/AUcpt5rlihcp8tuuhoXeWFGkWdYn
JKo3W2KXTs2R37LxvtXuIEdLUbhILNY8uy7lqy7HuoUdhNpXJ9iSjV1zmpF7PCxJoHDwmwk/borL
rVtx41lXwVv7FiaOArnaVc1QaWp7sj3NAizSIIgWoJNrrT5qMTOirTY+K4ZurXJuwB0lN+ksJRYm
cWc03QB38TqXfucsvKLn+0pCnz3LvLFDTJqr6XLoRjXGLGmB2zKUiE/6L/AKkFW2w20IOH/c3eEr
htl9e10CO9o37KQv+9JaZiElRVBRdMHJFEAg050sjwV+XMO1PDJzwZfWXeJJv3Y5Xcur5BrQUg1A
6riW2CbfyrOdfbotxghW1RLATZNsjXOxtvfnUufcC/BRh55CNp9N9ndpdT43B2o03fFTE+XUh25V
bs+1nbLddt+k2EExfb8paozuvYqteCMS+OpkhVfQmUshvKHQrijdhVLH6NmBGVpgiDi24BdLCoRA
Q7UcKA4XMK3auvkC655yvZ4pjUNNK6RhetH6MWokDa5xGlBT4Z6oIpVsfj67td+J9Qn3mXn2Tqx0
oHyGyINELy5Vlx7igmTqOJ2JC1hphnK72QHDFGKdgHdRIXogEZ278vkXrligQ63Bh4ZBLud7EoTz
EhUli2eKXcePYpfeI+51nwfZ4JZNEaDVJoH3ZXCnvbGt4wr8sOXRyiBVkKDkMykiYHjVJlNjKed9
AnR5Ww9X1lXORuT8+SmEPQ3Zkd9y69ekK177NnWduOxLAGdFCbm+c8qzUMArmyiaHdMqVn3kby8R
317DKbTM1LKoqYPUnVd8NQvhZvFYglLa67IRsxrw9V/Mzb2wNlgQQDV4EFvZ22B4fOYlcz8gr1q+
QcA69pGvzvMTTgt2TVLpdpH5nE5uFhjNpBcMDR+HliTNgNfgxpABb0JGo1RGB3SiR6QH2gOkcvaf
nJqLMHnwjf9ms53V7Z4FLS6BbXx7JPOgB9mj8vTwIPiIvNcMXb3op4+o4EW+OUZILNVjx0OVker1
VnDhvxytvZpLk0QGu4j8QHCfTr1YZNgBMOdtMYAxdFnjN8kZXxBp0HWu592wJqP89oo/tXxp61+L
bXs4FdcDBDvrj8d7+iZ0O+BK0O7PUjFr95BBdBGbZZ8oZhr66YhqJx9yc3HgGz5MW8GpJgd0Lv5s
OvqTGOjDXmA4gF8wznnhM0tA04eNulFvyhEJ4XjSWU0helU8ZvgjjdS7fulSREgyUAXsaidi7xaN
DldIFC6LbkIv4roaEFnvaA+vT02zL2Yb+I8MGOL7fn3hknAGmZNNojU/5p2g0LhDH+fIs2fyYgPm
FM8lfbjw/coZjGFCKEYQ/Yr2Vbab5Y1GoLydd0+yB/PqdKqunvU9ce4ojsecKQ3MkCaTaFyfTzwF
G+07uKIS5ipH6uQ9bpkhhfLo9XWK3v438LHTGZFYCwAMryP9TtFcgPDZ0OOJYuRV0YgDRF6J5SST
v/0S5B3uTRyD8sjDW8rOljitsMkv4ds2H+oRmI/HYvoAR8pnFigUytB4ArwggFFOXIbeGBbpLxF8
YlomP75Iu2fdzkvDIi8DtwjLpb9q+IERFSm9rVHOKgpwejpZAhIdLPOrXY4KkvblMd0Z94qjMtLE
vMwDTkbdkSao2epXgFgLx8eKbs/cgtEme/duQKPvJqFRZwgKHVPcdZHyHTdiUUo2hF0V/OdRYj75
/kPLtaVM0cM/NbVi4GQhBpU/Ta/mzPLEvjnxEJtaK56vC6zgE3m5JkfBqKwFfwTCvCFudd2rv+9a
4z/UIh9UjfbbhdvG+jyEkbMQSrfC56lcheoRvZsUUSD/mR/N65N+9GbltKR095uodUTQRYh8Ry9F
lWGnwkLiSFAvTjv9hgmAWkgtqI+7RwHGBFMGXgOLr9m0cZnjo95z9RTOfY/FFraZ6yxe8XT/irmI
KDB/3U1wRUqiOnSAkGjI3WuFgvxq8vnLjmR5KVm6wRGwUMW6SFG/eEb/ZyEnOX69Ye0AzB5GBEjB
A3FujlkKNd9JW5ygQVXXty+u0BT5gXtYrhVAMBSNOqqBqJ6weDS4dDC5M3xWepiSLqhhSIx61hTI
OxdlMDBWnJ0m2c2DslBkziyy59ELvJD+ZQ1OJGNVsewI50odJVJMqhhhjEFh0bnHxNQWydUfNFZu
lClFJgBeDV7uGWaIBmwOZTdsalXRMti7askLZLt/TSg74/C40IPihv3T0YG/AE3SzkTIxwO1pFEJ
Q2faQQ7aOqHSBx90bT5WVjn4lgqRu1aNEhgwlnrgYzR1cVoeAXtA70jCz5k05E884mLA2UnO6zyV
prpvG+JLFJSt2g22t+9pYrN5mcalObQ+Iwb9hx1cmz1mDm5MZ5/v9bPeke8DqerOTGLKZcfKkuWn
0TjR8zh673ORKjhIkY5KWxAoZaqZ+ICmUnqrtZIVzUKAoIKJ0CsvUBt5WRrXNvkEocQP2IqM7Zwc
myEe3UqDTG1kDfXlJhxvWb6EnLcfyUHNcr54EMLZIjGKLvOICCpavyN5gnYYx96Ebk0bmthV3fRe
ytLxGFy7+7hSkF/LNGlUsZ4+2MWslSBITi9SqA0cp/IbYYaDc1+PUdTLQMvhEGReNH9maBGm3SZv
c/yP+X3qfuObRkWx+G7TlWwWeJYYxpHG0fixODcm0FjeFwops6zVGnvoDpodEquRlPXxsWSyn+mQ
ujfZPon/RqHg0yS9C/BdIt4uRyZt5VlANypGn2zBIXx4kpTwFnsvN5si81bYzSH8YGy1xdaTJ5Oc
NvM8pa3R6xSYbNfD67BElpSSp6wgI1CtE6UQgMC+B0VP7GNnIz/76r1VeELkzBZDpjAd+zg+QAG4
UfMaec+wAGSFvjfNLOlMtyJUOJMTFiNykkinFMm5peXNiMhvdIr+XTSz3aEOBn8RUeM11TrMiByy
RD8YlZ7McRbQTaLy6fJuPEzci/SohefwJK5cF9j6FpbJWy2JyiIXz/0tDexV/QMre2mFxDBcwMXn
f100JHRKrfyNzhLc3s9Ul1ShlkDrizPF/NCJqZv/HlVoUpAd/E54HIfhxUA5Y9cRLRr4Aa+u/2yU
ADmybA/vLwfN5H5eAfU9J5iFcdTbW3icoGgESoAwe/YaabuZgeQ1qry5bhkoBuNLBsXQ8olY74V8
22S36cpCCMpf5wzqN/H1thnD5Gea7t48pDpCZSl/Cfg1bGp0glKIsDGqP4gXUCuUQb+arjtJXBH5
FTLca0x4QoQgFDR1CEAeYPMw8u3+lR+R+PfI3lSjnJrvqeJrUQ0lwYC8xsfo0oMm/11bshxyCJx0
lu3zUNtG7OvSnFtzLXJGRMrBTTmnB9FeuSEzq0EQC2kIGZQTkLCoS4vQp2Hx18dBbVsDO9JusEJ+
B3YkOEzcLFssytvTl64y9NI2wzqfGl9iN3MSpuAfvTte564yYL84Jji81TaY3cbXSSZOc/52U3+h
gceSLNH59VuF64NRJON1IPvdYMMaAnNcETVa9a+64C04e1Nl/X75W65M6aGkgmLC3YLx9AVHqFKi
0NDkFxoBItJKy8b/7Ge54+MDBnoSCTph22Voo+0shN9JaS2Ey2EXs/pphOfB2qEnSKJX8p7f0LQb
+QTKIkgU9dEzKr4qk/hu7P4bkOrVscDuEzpyaWHAe17g/xUNNBAgtEY92zTA2b9Ufr3+4Saleckq
ieCByJzy1TCflGKyyPXAtmi9zZEwxktmFXlu7nI/pwDUIU2rENiaM261pS/HQ+oONoSXOc+L+KLt
ubl8A6e9s5lskH8JnjI5HDgJpP2FrtuUFGWeJQ3bwZliX9S50WflUxzAmqi6Z3zSIQR/dbkJTMDq
qA5s7ke9mVL7WDtEkjoT4eXF6jEol1x2iKu7IBFFIaO4Ev+59p7/1NZqoT5M9mNW5MlHhDHzfvgW
p/wrpfTP8R2zzdcPgsgiL+MO2b4ZwhtM4x8SuFBfT48CA3K5lSIIj9Zib5ppkQekeU7VVjj6aldU
2ffgcjuj/cHjWKpXpYaLO8ijQlObuZCrUGIIG5X0FIT68HVKl7aoBbgxLlg2xvsKtIGfYITUpCbS
26AgE7zGonAkvhvMdyDm8AYZ4vp+aBqaPmQMBl3E6OqXuKeOiI8vtG3yL1pDD6yncfc6TRcZNXW1
Nf7XBpehUed+a/VVR9yOpFi2c8E+FfQRpGWk1w4UvSBQsw9p/9eL3JfnI8ICagGlG4y7AtQqi+zh
+RkuUV+SfZH4cnrIeHu+HxfM67D2HpCTbgS/dJUI7ZdY8unn/1QgBpinihxzbmKzVXvZX40C1GBa
XcObQVUvMbv+B4KviEUkqTzyMxJ9bc02tEJX6jmEInSLdgvKmX3vxdkFSJg9cUFo+oRWtm7RzKC0
ebw9qa/0hMjvE21tbDtAEM88XkJaqgQGxAljtPWHspo11zC+vV7zNhUQoCvaYpZIcWryRUgjAu8c
mU7qaY3rh9NA40l+Pz/o552PffTOLxfvO98LdhAklLp7rZaduV27vgIJv9S8OH6Pv064xptDBBFn
dh+eLU+9jM2HOp7i8Z6IOPzI7HYDFyekcawNrF5gGdoxvs2O6ST3xx/E37xzI03/knTLrAPlZt2l
bK2KWj1uUE6kffdbsktIgQoFipNIC2/RvW+kRiJONBqqsfJR0niXPNReIWa0PCpW+8kUa2SBRos+
83lafCMPpeua83cxltUGc+ElPWU+Jy5KMwW98L3O+ua2aiIvbN0CrsytQitYQfOwJGBXvp4rqK2q
J6S4z8QtqxotuJQMKruEPuX+zUc+AnZBVhIcKp5n+qr1baj4v6uLtpYSy4oohqABRa1mTdUohQ5e
MRXjFqKm7VhOfQWDJDDjX7Anexpm1s71ZprIF3RI/AezMMAKzIkhxbP7fBEO0voNUaCXk8y1NyEv
bBOs8qoSv6sRNCTJny65AEoWTyb+DvSveUcc1Bko877JCMvq2vIOSdEr+T4Wx0pYf9XqrmxShiu0
+3hi/FuUIG8dQ9bp21cr5fV+fRoRx4dctaT4hy7qpuvE4JIbE/kMBZ77OOsG3q0F/LU24G5EWC4q
x9kUMEf0fQc4GU3JWCGaSicglmH5g64Xx0CvbwfnUDynPug6KDsv1UJvqHqcy793HkaUPIjP7GZx
088pYJRXZyifi1LiQJ9tPOPStd/ziL7J4e4P+f9sRpDCuLJ/E6MTyIN8KKsKaw5SdWF7Zou2pbpP
9ZZM92LoHh5jjUcT5PQ5sWFwI9PF+7Lq7HU33cLBxHEtrMj+mwQ48ptCnQiKqvoa7Xm6QRKqCM/9
CtX67KfpIK3iBbVIQObGTW3uBWgEiznAJKi11wxLAof5+mrL1mtG6Fc52ksA6VigHfi0UTJIW8iT
i5R8usxmpq9zE+pSacKm0HaH3cNxEQXvc6h13bFAd+1uYfNkuQkuIejjJAqP+kQAiR0Xwde/9ByG
yj/UCw0GJOGyRv/JRh5G3Dp1GaYZq2d8MP3hK7m83UmQrXNttPXv2nT6HkSy8KktPNJxiWLd9Cf3
NAr0eHGLIgVXDkpgGljieFHneBPmYyHGLPgPqfD3PNTgbFv0cc/WcZG/sCcMsa6HYnu2cZZI73Ln
Kj1NkmaGv2bS9VryDeypp/1dv2Ddysh9HGvgucDDJ8/0qlV3WB/eKQtqehhQ5jcqPQZdBMUj/Tkt
56Yaq+b9laV5FPbJ3j8ZYQ8lEMd4PMQHYm+ikPhz94/HQtEzl7QS93n5nXF2J6LelrXyWwmyrX8f
sImbmrIAjmXmfw0WJL1UyESUUyLsug7uYcBZ0CEbSYKDszW3Reqz7FXYE39Cmhu2mb5SZcJZ3H7o
485lwHHw33KE5qMV/1NM2vnl2qQm1fchT3rjjcOPaktNC5a2S7YbTCTwYJHsQO4eyFuuJb1IMUWw
kkMhrGNH3mLNSeYLwbOnUJE01fim26G+ONGWApJ/SgECWbYZ6u/wy7FtW8aOLIcLZcEMDCGD5PiE
ixBIr868rNTWMlbvE2IR61nASrQKqC4BLZPNl5u0wuZ4iv57GOcrbm4iE0e3/weRG38cpUkQ4A0c
zE+95ayt45wzwxOx/eRdZErA3sszHrUJh7xBtx6YTvpPaW4sz2D+1K7ZtMXOE9ehRJg5cpw27ofv
7G6mrjyEOK7XBYo4rDXmAE/+7RM4hU2WqoaeDyjfMaoQ/vu7yZ6aUdjV5djAtZ2RG4niWLyfcG5U
ubT1+H+i1geBKrjFuKdXCL0TFy/xGFKMADjfCiCLmDVJFZtr0xLdwS3vxdRqtKgfTJF9lEG26+DW
82TrddB37ditTR+qU1rQ7xyO8pds9G+hsP6myTv7ociYwmXjbtr7CmjYxJHixRJMPEBUTly3a7Cx
YJVDcXSOiA3X5Espai8aa2tysh4XTdjENk2xluibzOQX60jUtAvpa1zjgpy7HGNxU9GBS172axxB
frMfHqSUnHzAl1wdAGlxzrHNGd1a6SovEdcpY2gnkQHmtFt9n8cpni4ycVmHDd+9V3LWPcbGSG+w
HJrndYynt0wHsH6PTtNXJRD10Aq8h+xwOqq0wb2OUcQVE6B7g0EdCx1fVjkli38UUAhM22ZOBhay
qJ11KYQF/Iqbzq81JQm77eiOJvN9CL9TmYa8zsNUz6asnnA3ynVj+BdPdiTWA4JZTiNjkiy0B0qs
0i5QEr542Igfg98QNAhyI1E9zM8XuRjriJ+2bYrnEEjn2GJdErI81QPJUL5zf1F1s64gJ2UuK3QK
13MPoWGqOL17qt9P1p1Ynt1W3Mf78tShmGgrAapUNEaLtHmtn/joNdKN4xyiSb1rgzn0/Ikn09JE
bnVxeXwnKjcpj1ivom6h84jr0VLQ427zNQDrl3elHEKHxWQw6VpS/GsPbO6GSMulS3QWUWhol+Q3
MlnpCh2a8I6idPmlzaJk55kU+w3F4t0vMyXX+5s28PQvwibWovQVXU4prkWLYBa0JAebqTKjVMsg
dupn8YBZrF7SsJh2by+2TfwhT1OB3q3jh+Gox9TKY2WysuUeoNVQMTj6O2uQm7M4/RJopVuv5uh0
65tRa1Zh4Fbnge3KpRneF7icGf/oYffuIPxUvtKR8FgV0eK18/PmR4Iq84Oe1KWSIS0NgNmmSu0O
S0uCD89HGdRPPddA7T+nQciHNIQrUfpJT/HIW+ADMpuOruscTdtHrOV6VzVmIhVdGNDKY5hcTUls
vsbvEvGUophTEpjre4gRnHJu/9Wb7zegDauECFaSgZTp12Ehh7leQqor2LbXeqPGozKOydiHJp6p
HqSSbcN/gG2E3wX6JIihd4OsHSOjA/FZ5EL/PmUseo8ew6m3b4H0HrQZ90SEOTsyOLIi5pwof3bB
y8Zzatv5wfNhOpenVebNjrGpTvIzM5DLrs5l+x84ONwFRSWqu7mJpHyXs5u9EX7poYaz5OOEhc8D
vuYewLqi/PdYk0Y0AmSlHzReS14LcyAA9J7HoR1r5rxhSSrFJyfJYk+3N+deYr2FiWFilO3BB0vQ
vv/ywt/4WO5dl0XUjA2r/8FWIUiVEb+v8WyY+d7w8DTnM4VlypmF25MlOdaFbsMSlgrs7PwX3q2G
Z3LuesCLM6bZh/rWwl8LI9NHVlJcDIU70p/LeU2HP3P8Eq7o8YdGEqNr2QnP+SO5qdJgZQHbUtW8
oCJacJ3479c6P/e229VCoScjNYYaXq5nAteELLEYE/SZRBw3znvSDJwK4Fe1C8c5YNabbtSU6fyn
X4gxTAjW4S7a4LLbYxhRxEiAGwIPz6M3lB1eHSc0zDsPuFOQMjXQi5PgnwbG4xTf0LuXmBQjKYPg
Luy0M2Fs5i2SfRN7vBMlzsag+fZTcOEe3lWPbwFyoRYKPVrQeKQYAwtkDsQ+ogxe8ZpimDyiosLo
oU4qhDJ+Qo6tP70RFreFr5e8W7wcQyeId1T5UCLC2mCZLxcFbZUFvYFHaAFaAVxvAyhNgDsnSS81
dakjs535IMUo8gWodbaC+UwGFWPTCjPiGHn4siRgaKIixwg8DTXwv+UdIt7SviZsgXZ4Pe6ESn/k
XrfjDvbRTgMm6QUFyXdNCEvhU2uKypjiwau0rjeMSFKcoHPd/G5wjePkXAbWH5Lso67d1qHNT7mG
uG8MDsnMnssH9Y8edlPIVSbk5Mth6rxpd936l8Aqpt9BaRJZJ/pijMRH3ADCU8tGXS8BDu9c7+ja
qTsUN4c7PnYRQb+msziUxEjn365KDYfrUCuqLYv4JJ+J01NLZYeqcyW89HYpy5wvZN8+UeUsjH3t
OffMbYpH6vj58nGheMgQFqeb2ybLNu6eFZgnog0sKxhExwf01UjHYF9X7p/QZjzqZeHUlze2G85M
pT0IpK1NMaMh08I0c6dZJaMf/AsC+5oWHTUDo4BNOKfzQU2E1rNftpSobH5GJihihjERCEMxFV38
f63h45NApi+JCMfe+Crs57OnqlKXlJW7iB6skn6u7muzO434nJSvoWDQgbK7mr8WdVXXHxcrnC3g
Ipxj4zLChpuO35W+RG8eqjPnD5Q/wudpvxJ+w/maiZ0d0lE9j7MLIhrUrH8pGNzTkHaoyUwYeU3k
+/g1CsTmtrSULq+hZdqdzlcIIoextjtYdJCkJ1p2A7YXSIWVYbywIX5/XUh6n9M6NV7D3W8+0ntG
XgYtD1sdC3m3bnLPL1yMojj0cspqVny9qHTaUOZudBvB4/KVE4Ufku80RAssY3I4Fk44zqb42GM3
p4S5MLy7CzVpGF54pY/pSyDMNFfz0Oty4aJGJprconESU+Rj+39z93rUqyk8GtqCis1FrxznNMXN
c9GMgK9XUP7a0/araBDKrbFBkLy2TgMs6wP5nxIkpXjf2aawHo0YZOA1fmCdK1hNJI2893CswITF
C05ALg0u8f156oJSHZH7Vw4mgx/b1O87aCd4gTm3lRR/BVD8Z9X3/KFFhqidjHMXIDXslg7LLQsX
5WjofpvPkMo1zMPR63AbXePw+76TspaDEDDaFwN9bF+56slFa0dknue5steZWCwAOGSDcWf4mE8N
dkwcRb62XOfPL8hDY6IVcni/4YZ6x10BWJIpq11gB1Xcsvyog0Qk9vBm2j9jvNl0UyTM8rEL9dMV
F/HeOeq2SVDg4+BLQ6GACqAjtOrESVJJ3RsrWv9QokswPb9LF1IvFlWUPQhQM92QXQ8gOQXad0b0
r2wBSsrBMhASLkdd/JTJe23/wquiKYmbxvnBxtEOV7xda3/k5sP9jOcZtU12ESyANd4j3D0fMrBR
bNaaGCNaKnphJVMl8NlnBpiBRmSk9ZkvhzV3pmbRN9RDzjjILzt9x3i0fhS8MirIXYKwcfllMKr4
ONlTGzI8h8vw9b3b9F8hB+NAVErlowIS+q5J4dW8dz0qykc0IYwg22/f379GT9oqVPLe6xeJ6zKA
YtK8oiX1m/OXgNYZqPgo7uQ+OlpyZf276qWZASBMg6tr/KaHTRUiGcGyz4hQRQstMwLng7EU6ikR
+NzdSEFfmSXSdkryUTPbex8Au7eZwbkyLBDXrcesl9+GCwVcQZgohlheFgnU0bXI9fhRnGN0OeLd
E7KIVsOJ6JSQxcAtYz8kb+vgrnRlrN4J2YyUPRY4uQi0YcpL9z1fX7rBeRziLcFdIZyqsF5VkhNb
EFgayat84khTsMZmrbKnwbIUzNN8pYgsdWIm/IycfpcpJAsaAfAls4WLpwuXVEDrZ2Ks2tqZPe+G
eTL+mTtDgvSh5uCBh0ijfNUrEoxREuEGn53+sIzf61ixyN7mkZWvE3g3B0tIo+9vtxwCv7se+W9F
2MtZ7TpkLXO9qHjdUc19pZnGBCDCj1zWFk2XkgJ91kY77AHu4crRvpLHhCfV9BLMxQEKiM/Bc4RZ
XPx04zTlnCX9HF1b8UMfxuhTnGJos1C5Y+DHFVrwD3mOKCgXUCHp4nMmmX8sYLaFLZZZbvEhX6Ix
6EBXCRTo90kMh0elN4H4PpC51r8VZ5MMMF84qANJnKhvPpPhe+XuQ6J77XBLJg2Etl4LiOLfh7Uk
hLVJHaAP0GTXQZbH5bRK5cT4tIqP6SZXb0xrTdZSzsAg1Oa+7dQPSTyYMO6Rrigi611+W9IJB6YX
yyLRWq3DMKqLMGwTQn6CLpjwujS774mEHtOkOLzjr8NgIEA/ScKOHccCmQNZrHsx/PolqDlY+WzC
G/pp03JERRKyWPI4OMX8jQ0YndFJCkN4WM1bSzltK68R5X5qK5f45y844+uXbAmtcAFVPINbIDdo
Gvspdl2XYSI2rxp/NJP5+oLKRPBwtNURIB6IBinC3MzD14nRhV9wMAdv5cIVqH4Z9dd0m5tFUos3
cb0uWgwxHlghZNyYO7JqlbK9BhgkG2eoXaiL6GznDGkG7M4nj+2LBSb/r5ZHE1c2LKknY3OOik+6
SzXoAdaXLKehHv8bYpyOMRs8h3gVyOoRJoy585ms1jAtlsGUy+aI3jyUWM8Gn/lhYEjbj8RLfCf9
AVtAjbETOveadNCASE8EfvP0TRXSNlTJOKM4Dr7CNuyc6N1YWDHTWPEjaHuBPK7Y/uV+dVUoX3O2
xsSjLSrWKsmd825nC2Fbe1P9TawIt8ezKWrLd23da9EzeZN93AF/pTGO3Dx91hgDDHlbmdXpVcKc
7wO+I9vBmerCcJRFrMmyXYwIb4AnwYdxmJD+Ai+IrtWLUHOinbfhT4Zqv7R90SKqAA3Wpasx2JBf
BqmHb26ZOdT2rhZ4tyz2BRWQaIqDtKL5mni/9FmknpVIFUpmi2d6dE6JquHnODN2AONDFdKZfT1Y
RbpguiOcd52IP5RYoU4OP4HQ26C3fjZz9MmTP4azoHr1J0ZB6b0z09tzTW5XWekMpM2xgqhM/Mhg
kuO9ph1xWAXxLa+iEvO+AC8I50z0MwP3q0rkBsPY6JgSjDpKLiERROZLJ9IxR7Rnv1TCWvapgVtw
K7Hltiy2aKYZXhy/PY1twkaRuNgznHQvhzo7dWXUfAvJ3Dq5g74g3DGNU9tad8I3MGUQ8ZtoQrEn
eUqX+S0eeyN3r0yxM74A61Mv9n7FHBaYTa4C3/EDCB2YSryAj4YGgNqH650Hly6wb0vm4gc0iki4
tM8C5Ow3aTPMbeeF44BJYn/FRWNJYk3OqndLjdOULU8M5CJUmeD+q/j0cBRe1Q2OktRMQe8MdR45
c9B05Zh5Jy6Ot5LXtibwGLiXWX5E/sfngCR/aI0OeTDgniG8Q69jQ8XMNkYpWsfyB6UnWSqpoNQ/
0LJr4A2zrUsToJ57RmihwgPn9uleBjBaoEy0P9Kyrv7K7BWP+FeBzbv78t7YMqQamoMSE20pgJbp
BvpIGSXL25n89mHE6+GqmZuRIiDwz3WZS0JeGzjRVqje6Dr2Y7DznLonVcGFaNCeEzRd++kq8cM9
PKecnR3eng2QmquhCuKgIgtON9W7co/mIu9cdYhCGIY/gGXeRHWC+4Lk8wtb8NiO85jgYmfUxW6A
Xo4lnjVBi090ecLk/ObIK9OHqig9uqPcWF7dVb5cLic9oUldYH4U4BIIc8m27Rtng4sPghCLw5Jv
U1OJue58qtIdIeY5NfZ0wUZ9NhVPqXdEUohAiEF2SknXeYa6hLE4tWy+1Zov9bYNtr1uJ/1pf3kV
ZB4eh1LYRhhoHNa/7WE5Dr2fXZTgXqOLkcRz8562J+kW880FB8gYrORVZguVZr19YFSoFZWBgLG3
TCIuhka8HuG+ZgsjrB6p7qgn8nCgQQ8acc5s+yq2JH5jovm4z2WqAdpWwjnH6XzWy0HfJXYJVHKi
LARlTSDgez9oJO+GwUmA6ajzjr2COiNdCPNnKo+K0K6KjHWQ51Nr1sffnVZ/b2K4VwAjjkJDXHQg
uLcZmajO6PzZBkkkUMA4tOSSPFKt7Ic+lkjYTAEpYBInZcIuBpYx2j+l//od8hQBHQD/vZ6BYfmK
m0tdLGzQBGz9GW01t3NgskoDlEzobhS8Bjcr67ffybQf2KxNZC2O9xjnOJIUKHG2qtOrUKJ+sGne
wbn2UipH/x4+B4xEbKv0V6rEhqZ2Cqc=
`protect end_protected

